* NGSPICE file created from Core.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

.subckt Core clock io_dbus_addr[0] io_dbus_addr[10] io_dbus_addr[11] io_dbus_addr[12]
+ io_dbus_addr[13] io_dbus_addr[14] io_dbus_addr[15] io_dbus_addr[16] io_dbus_addr[17]
+ io_dbus_addr[18] io_dbus_addr[19] io_dbus_addr[1] io_dbus_addr[20] io_dbus_addr[21]
+ io_dbus_addr[22] io_dbus_addr[23] io_dbus_addr[24] io_dbus_addr[25] io_dbus_addr[26]
+ io_dbus_addr[27] io_dbus_addr[28] io_dbus_addr[29] io_dbus_addr[2] io_dbus_addr[30]
+ io_dbus_addr[31] io_dbus_addr[3] io_dbus_addr[4] io_dbus_addr[5] io_dbus_addr[6]
+ io_dbus_addr[7] io_dbus_addr[8] io_dbus_addr[9] io_dbus_ld_type[0] io_dbus_ld_type[1]
+ io_dbus_ld_type[2] io_dbus_rd_en io_dbus_rdata[0] io_dbus_rdata[10] io_dbus_rdata[11]
+ io_dbus_rdata[12] io_dbus_rdata[13] io_dbus_rdata[14] io_dbus_rdata[15] io_dbus_rdata[16]
+ io_dbus_rdata[17] io_dbus_rdata[18] io_dbus_rdata[19] io_dbus_rdata[1] io_dbus_rdata[20]
+ io_dbus_rdata[21] io_dbus_rdata[22] io_dbus_rdata[23] io_dbus_rdata[24] io_dbus_rdata[25]
+ io_dbus_rdata[26] io_dbus_rdata[27] io_dbus_rdata[28] io_dbus_rdata[29] io_dbus_rdata[2]
+ io_dbus_rdata[30] io_dbus_rdata[31] io_dbus_rdata[3] io_dbus_rdata[4] io_dbus_rdata[5]
+ io_dbus_rdata[6] io_dbus_rdata[7] io_dbus_rdata[8] io_dbus_rdata[9] io_dbus_st_type[0]
+ io_dbus_st_type[1] io_dbus_valid io_dbus_wdata[0] io_dbus_wdata[10] io_dbus_wdata[11]
+ io_dbus_wdata[12] io_dbus_wdata[13] io_dbus_wdata[14] io_dbus_wdata[15] io_dbus_wdata[16]
+ io_dbus_wdata[17] io_dbus_wdata[18] io_dbus_wdata[19] io_dbus_wdata[1] io_dbus_wdata[20]
+ io_dbus_wdata[21] io_dbus_wdata[22] io_dbus_wdata[23] io_dbus_wdata[24] io_dbus_wdata[25]
+ io_dbus_wdata[26] io_dbus_wdata[27] io_dbus_wdata[28] io_dbus_wdata[29] io_dbus_wdata[2]
+ io_dbus_wdata[30] io_dbus_wdata[31] io_dbus_wdata[3] io_dbus_wdata[4] io_dbus_wdata[5]
+ io_dbus_wdata[6] io_dbus_wdata[7] io_dbus_wdata[8] io_dbus_wdata[9] io_dbus_wr_en
+ io_ibus_addr[0] io_ibus_addr[10] io_ibus_addr[11] io_ibus_addr[12] io_ibus_addr[13]
+ io_ibus_addr[14] io_ibus_addr[15] io_ibus_addr[16] io_ibus_addr[17] io_ibus_addr[18]
+ io_ibus_addr[19] io_ibus_addr[1] io_ibus_addr[20] io_ibus_addr[21] io_ibus_addr[22]
+ io_ibus_addr[23] io_ibus_addr[24] io_ibus_addr[25] io_ibus_addr[26] io_ibus_addr[27]
+ io_ibus_addr[28] io_ibus_addr[29] io_ibus_addr[2] io_ibus_addr[30] io_ibus_addr[31]
+ io_ibus_addr[3] io_ibus_addr[4] io_ibus_addr[5] io_ibus_addr[6] io_ibus_addr[7]
+ io_ibus_addr[8] io_ibus_addr[9] io_ibus_inst[0] io_ibus_inst[10] io_ibus_inst[11]
+ io_ibus_inst[12] io_ibus_inst[13] io_ibus_inst[14] io_ibus_inst[15] io_ibus_inst[16]
+ io_ibus_inst[17] io_ibus_inst[18] io_ibus_inst[19] io_ibus_inst[1] io_ibus_inst[20]
+ io_ibus_inst[21] io_ibus_inst[22] io_ibus_inst[23] io_ibus_inst[24] io_ibus_inst[25]
+ io_ibus_inst[26] io_ibus_inst[27] io_ibus_inst[28] io_ibus_inst[29] io_ibus_inst[2]
+ io_ibus_inst[30] io_ibus_inst[31] io_ibus_inst[3] io_ibus_inst[4] io_ibus_inst[5]
+ io_ibus_inst[6] io_ibus_inst[7] io_ibus_inst[8] io_ibus_inst[9] io_ibus_valid io_irq_motor_irq
+ io_irq_spi_irq io_irq_uart_irq reset vccd1 vssd1
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09671_ _09688_/A vssd1 vssd1 vccd1 vccd1 _09727_/A sky130_fd_sc_hd__buf_2
XANTENNA__18828__D _18828_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18869_ _19293_/CLK _18869_/D vssd1 vssd1 vccd1 vccd1 _18869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14210__S _14218_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09287__A1 _12935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16137__S _16145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10974__A _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14446__A _14650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15976__S _15984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09995__C1 _09602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16493__C1 _12749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09938_ _10283_/A _09937_/X _09696_/A vssd1 vssd1 vccd1 vccd1 _09938_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09869_ _10176_/A _09863_/Y _09868_/Y _09936_/A vssd1 vssd1 vccd1 vccd1 _09869_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11601__D_N _11534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _12097_/A _11855_/X _11899_/X vssd1 vssd1 vccd1 vccd1 _17690_/A sky130_fd_sc_hd__o21ai_2
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14120__S _14120_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12645__A_N _12651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _12880_/A vssd1 vssd1 vccd1 vccd1 _12880_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10868__B _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11831_ _16268_/A vssd1 vssd1 vccd1 vccd1 _16213_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12806__C1 _12805_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14550_ _14550_/A vssd1 vssd1 vccd1 vccd1 _18852_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11381__A2_N _11380_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11762_/A _17429_/A vssd1 vssd1 vccd1 vccd1 _11763_/B sky130_fd_sc_hd__nor2_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _16925_/C _12775_/X _12777_/X _19702_/Q _13500_/X vssd1 vssd1 vccd1 vccd1
+ _13501_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11180__S1 _11179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10713_ _09707_/A _10706_/X _10708_/Y _10712_/Y _09739_/A vssd1 vssd1 vccd1 vccd1
+ _10713_/X sky130_fd_sc_hd__o311a_1
XFILLER_42_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14481_ _18414_/A vssd1 vssd1 vccd1 vccd1 _14481_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11693_ _17379_/B _11693_/B _11693_/C _11693_/D vssd1 vssd1 vccd1 vccd1 _11693_/X
+ sky130_fd_sc_hd__or4_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _16219_/A _16219_/C _16219_/B vssd1 vssd1 vccd1 vccd1 _16220_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13432_ _13432_/A _13432_/B vssd1 vssd1 vccd1 vccd1 _15276_/A sky130_fd_sc_hd__and2_4
X_10644_ _11386_/S vssd1 vssd1 vccd1 vccd1 _10644_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__15771__A1 _15770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15886__S _15890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _16151_/A vssd1 vssd1 vccd1 vccd1 _19490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10575_ _10571_/A _10572_/X _10574_/X _10307_/A vssd1 vssd1 vccd1 vccd1 _10575_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13363_ _13363_/A _13363_/B _13397_/C vssd1 vssd1 vccd1 vccd1 _13363_/X sky130_fd_sc_hd__or3_1
XANTENNA__10596__B1 _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15102_ _15102_/A vssd1 vssd1 vccd1 vccd1 _19083_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_23_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12314_ _12314_/A vssd1 vssd1 vccd1 vccd1 _12314_/X sky130_fd_sc_hd__clkbuf_4
X_16082_ _13178_/X _19460_/Q _16084_/S vssd1 vssd1 vccd1 vccd1 _16083_/A sky130_fd_sc_hd__mux2_1
X_13294_ _13454_/A vssd1 vssd1 vccd1 vccd1 _13358_/S sky130_fd_sc_hd__buf_2
XANTENNA__13534__A0 _19923_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15033_ _19053_/Q _14433_/X _15033_/S vssd1 vssd1 vccd1 vccd1 _15034_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19910_ _19919_/CLK _19910_/D vssd1 vssd1 vccd1 vccd1 _19910_/Q sky130_fd_sc_hd__dfxtp_4
X_12245_ _17199_/A _12267_/C vssd1 vssd1 vccd1 vccd1 _12245_/X sky130_fd_sc_hd__or2_1
XFILLER_123_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10443__S0 _10390_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19841_ _19876_/CLK _19841_/D vssd1 vssd1 vccd1 vccd1 _19841_/Q sky130_fd_sc_hd__dfxtp_1
X_12176_ _11818_/X _12088_/B _12175_/A vssd1 vssd1 vccd1 vccd1 _12176_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11127_ _11127_/A _11127_/B vssd1 vssd1 vccd1 vccd1 _11127_/X sky130_fd_sc_hd__or2_1
X_19772_ _19817_/CLK _19772_/D vssd1 vssd1 vccd1 vccd1 _19772_/Q sky130_fd_sc_hd__dfxtp_1
X_16984_ _19753_/Q _19752_/Q _19751_/Q _16984_/D vssd1 vssd1 vccd1 vccd1 _16994_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18225__A0 _19968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18723_ _19314_/CLK _18723_/D vssd1 vssd1 vccd1 vccd1 _18723_/Q sky130_fd_sc_hd__dfxtp_1
X_11058_ _18966_/Q vssd1 vssd1 vccd1 vccd1 _11059_/A sky130_fd_sc_hd__buf_2
X_15935_ _15935_/A vssd1 vssd1 vccd1 vccd1 _19394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10009_ _10910_/A vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18654_ _19503_/CLK _18654_/D vssd1 vssd1 vccd1 vccd1 _18654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15866_ _13178_/X _19364_/Q _15868_/S vssd1 vssd1 vccd1 vccd1 _15867_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14817_ _18961_/Q _14462_/X _14819_/S vssd1 vssd1 vccd1 vccd1 _14818_/A sky130_fd_sc_hd__mux2_1
X_17605_ _17688_/A _17602_/X _17694_/A vssd1 vssd1 vccd1 vccd1 _17921_/A sky130_fd_sc_hd__o21ai_2
X_18585_ _19560_/CLK _18585_/D vssd1 vssd1 vccd1 vccd1 _18585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15797_ _15796_/X _19347_/Q _15801_/S vssd1 vssd1 vccd1 vccd1 _15798_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17536_ _17958_/A vssd1 vssd1 vccd1 vccd1 _17725_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14748_ _18926_/Q _14468_/X _14750_/S vssd1 vssd1 vccd1 vccd1 _14749_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16465__B _16465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__S1 _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17467_ _17467_/A vssd1 vssd1 vccd1 vccd1 _17601_/S sky130_fd_sc_hd__buf_2
X_14679_ _18299_/A _14917_/B _18295_/A _14844_/D vssd1 vssd1 vccd1 vccd1 _16134_/B
+ sky130_fd_sc_hd__or4_4
XANTENNA__10794__A _10794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19206_ _19302_/CLK _19206_/D vssd1 vssd1 vccd1 vccd1 _19206_/Q sky130_fd_sc_hd__dfxtp_1
X_16418_ _13376_/X _19566_/Q _16426_/S vssd1 vssd1 vccd1 vccd1 _16419_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17398_ _17507_/S vssd1 vssd1 vccd1 vccd1 _17504_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19137_ _19395_/CLK _19137_/D vssd1 vssd1 vccd1 vccd1 _19137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16349_ _16353_/B _16348_/Y _16303_/X vssd1 vssd1 vccd1 vccd1 _16349_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19068_ _19290_/CLK _19068_/D vssd1 vssd1 vccd1 vccd1 _19068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18019_ _18019_/A vssd1 vssd1 vccd1 vccd1 _18019_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10733__S _10735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16475__C1 _12908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16420__S _16426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10034__A _10040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18216__A0 _19964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09723_ _09723_/A vssd1 vssd1 vccd1 vccd1 _09724_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10969__A _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12500__A1 _10137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09654_ _09723_/A vssd1 vssd1 vccd1 vccd1 _09787_/S sky130_fd_sc_hd__buf_2
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ _11491_/A vssd1 vssd1 vccd1 vccd1 _10623_/A sky130_fd_sc_hd__buf_2
XFILLER_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12264__A0 _12260_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11162__S1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16806__D _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12395__S _12395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14176__A _14222_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15753__A1 _19908_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10360_ _19913_/Q vssd1 vssd1 vccd1 vccd1 _10360_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10291_ _10312_/A vssd1 vssd1 vccd1 vccd1 _10291_/X sky130_fd_sc_hd__buf_2
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12030_ _12116_/A _12024_/Y _12029_/X _11977_/X vssd1 vssd1 vccd1 vccd1 _12030_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10425__S0 _10367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18207__A0 _19960_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13981_ _18626_/Q _13710_/X _13983_/S vssd1 vssd1 vccd1 vccd1 _13982_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10879__A _11319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15720_ _15719_/X _19333_/Q _15720_/S vssd1 vssd1 vccd1 vccd1 _15721_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09452__B _18343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12932_ _12932_/A vssd1 vssd1 vccd1 vccd1 _18437_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17430__A1 _12553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15651_ _14663_/X _19317_/Q _15655_/S vssd1 vssd1 vccd1 vccd1 _15652_/A sky130_fd_sc_hd__mux2_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _13343_/A vssd1 vssd1 vccd1 vccd1 _12863_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14602_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ input62/X vssd1 vssd1 vccd1 vccd1 _18370_/Y sky130_fd_sc_hd__inv_2
X_11814_ _11763_/B _11766_/B _11763_/A vssd1 vssd1 vccd1 vccd1 _11815_/B sky130_fd_sc_hd__o21bai_4
X_15582_ _15582_/A vssd1 vssd1 vccd1 vccd1 _19286_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _18198_/A vssd1 vssd1 vccd1 vccd1 _18413_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17321_ _19882_/Q _12880_/A _12883_/X _11665_/B _17355_/A vssd1 vssd1 vccd1 vccd1
+ _19882_/D sky130_fd_sc_hd__o221a_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _13793_/X _18845_/Q _14535_/S vssd1 vssd1 vccd1 vccd1 _14534_/A sky130_fd_sc_hd__mux2_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11745_ _12116_/A vssd1 vssd1 vccd1 vccd1 _11745_/X sky130_fd_sc_hd__buf_2
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17152_/Y _19851_/Q _17258_/S vssd1 vssd1 vccd1 vccd1 _17253_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14464_ _14464_/A vssd1 vssd1 vccd1 vccd1 _18823_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15744__A1 _18451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11676_ _11678_/A _12606_/A _11648_/A _11638_/A _12602_/A vssd1 vssd1 vccd1 vccd1
+ _11676_/X sky130_fd_sc_hd__a2111o_1
XFILLER_168_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _16203_/A vssd1 vssd1 vccd1 vccd1 _19514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13415_ _19948_/Q vssd1 vssd1 vccd1 vccd1 _16332_/A sky130_fd_sc_hd__clkbuf_2
X_10627_ _11438_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _10627_/X sky130_fd_sc_hd__or2_1
X_17183_ _17242_/B vssd1 vssd1 vccd1 vccd1 _17195_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_167_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10119__A _10909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14395_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14395_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16134_ _16134_/A _16134_/B vssd1 vssd1 vccd1 vccd1 _16191_/A sky130_fd_sc_hd__nor2_8
XFILLER_127_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13346_ _19757_/Q _12892_/X _13345_/X _12896_/X vssd1 vssd1 vccd1 vccd1 _13346_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10558_ _10569_/A _10558_/B vssd1 vssd1 vccd1 vccd1 _10558_/X sky130_fd_sc_hd__or2_1
XFILLER_128_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16065_ _13009_/X _19452_/Q _16073_/S vssd1 vssd1 vccd1 vccd1 _16066_/A sky130_fd_sc_hd__mux2_1
X_13277_ _15244_/A vssd1 vssd1 vccd1 vccd1 _13277_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10489_ _18652_/Q _19243_/Q _19405_/Q _18620_/Q _10439_/S _10397_/X vssd1 vssd1 vccd1
+ vccd1 _10490_/B sky130_fd_sc_hd__mux4_1
XFILLER_108_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15016_ _19045_/Q _14408_/X _15022_/S vssd1 vssd1 vccd1 vccd1 _15017_/A sky130_fd_sc_hd__mux2_1
X_12228_ _12228_/A _12257_/A vssd1 vssd1 vccd1 vccd1 _12232_/A sky130_fd_sc_hd__xor2_4
XFILLER_69_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19824_ _19859_/CLK _19824_/D vssd1 vssd1 vccd1 vccd1 _19824_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12159_ _12026_/X _12154_/X _12155_/X _12158_/Y vssd1 vssd1 vccd1 vccd1 _12160_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_150_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09643__A _10968_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19755_ _19756_/CLK _19755_/D vssd1 vssd1 vccd1 vccd1 _19755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14483__A1 _18324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16967_ _19748_/Q _19747_/Q _16967_/C vssd1 vssd1 vccd1 vccd1 _16970_/B sky130_fd_sc_hd__and3_1
XFILLER_84_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11384__S _11384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10719__S1 _10754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__A1 _11170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18706_ _19553_/CLK _18706_/D vssd1 vssd1 vccd1 vccd1 _18706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15918_ _15918_/A _15918_/B vssd1 vssd1 vccd1 vccd1 _15975_/A sky130_fd_sc_hd__nor2_4
X_19686_ _19720_/CLK _19686_/D vssd1 vssd1 vccd1 vccd1 _19686_/Q sky130_fd_sc_hd__dfxtp_1
X_16898_ _16898_/A vssd1 vssd1 vccd1 vccd1 _16919_/A sky130_fd_sc_hd__clkbuf_2
X_15849_ _13009_/X _19356_/Q _15857_/S vssd1 vssd1 vccd1 vccd1 _15850_/A sky130_fd_sc_hd__mux2_1
X_18637_ _19484_/CLK _18637_/D vssd1 vssd1 vccd1 vccd1 _18637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09370_ _20013_/Q vssd1 vssd1 vccd1 vccd1 _12688_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12246__B1 _11890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18568_ _19449_/CLK _18568_/D vssd1 vssd1 vccd1 vccd1 _18568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13612__B _18297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17519_ _17549_/A _17549_/B vssd1 vssd1 vccd1 vccd1 _17798_/A sky130_fd_sc_hd__or2_1
X_18499_ _19482_/CLK _18499_/D vssd1 vssd1 vccd1 vccd1 _18499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11413__A _11562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12549__B2 _12548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12943__S _17808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16415__S _16415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09818__A _09899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16999__B1 _16860_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09706_ _09706_/A vssd1 vssd1 vccd1 vccd1 _09707_/A sky130_fd_sc_hd__buf_4
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09637_ _10264_/A vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13803__A _14628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09568_ _09761_/S vssd1 vssd1 vccd1 vccd1 _09568_/X sky130_fd_sc_hd__buf_2
XFILLER_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09499_ _11481_/S vssd1 vssd1 vccd1 vccd1 _10824_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11530_ _11603_/A _11530_/B _11530_/C vssd1 vssd1 vccd1 vccd1 _11604_/A sky130_fd_sc_hd__nor3_1
XFILLER_169_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15726__A1 _15724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__S0 _10893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11461_ _19513_/Q _18925_/Q _18962_/Q _18536_/Q _10649_/X _10754_/A vssd1 vssd1 vccd1
+ vccd1 _11461_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14634__A _14634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18125__C1 _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13200_ _19784_/Q vssd1 vssd1 vccd1 vccd1 _17070_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10412_ _09750_/A _10401_/X _10410_/X _09757_/A _10411_/Y vssd1 vssd1 vccd1 vccd1
+ _12656_/B sky130_fd_sc_hd__o32a_4
XFILLER_109_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17479__A1 _17866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14180_ _14180_/A vssd1 vssd1 vccd1 vccd1 _18710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10646__S0 _10644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11392_ _11395_/A _11389_/X _11391_/X vssd1 vssd1 vccd1 vccd1 _11392_/Y sky130_fd_sc_hd__o21ai_1
X_13131_ _13115_/A _13132_/C _19932_/Q vssd1 vssd1 vccd1 vccd1 _13133_/A sky130_fd_sc_hd__a21oi_1
X_10343_ _18591_/Q _18852_/Q _18751_/Q _19086_/Q _10390_/S _10333_/A vssd1 vssd1 vccd1
+ vccd1 _10343_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10274_ _18592_/Q _18853_/Q _18752_/Q _19087_/Q _09924_/S _09929_/A vssd1 vssd1 vccd1
+ vccd1 _10274_/X sky130_fd_sc_hd__mux4_1
XANTENNA_input55_A io_ibus_inst[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ _19928_/Q vssd1 vssd1 vccd1 vccd1 _16219_/A sky130_fd_sc_hd__buf_2
XFILLER_152_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12013_ _16226_/A _12011_/X _12012_/Y _11668_/X vssd1 vssd1 vccd1 vccd1 _12013_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_78_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17870_ _17705_/X _17862_/Y _17868_/Y _17869_/X vssd1 vssd1 vccd1 vccd1 _17870_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16060__S _16060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09463__A _12933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16821_ _17073_/A vssd1 vssd1 vccd1 vccd1 _16845_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_181_clock clkbuf_opt_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19768_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16752_ _19688_/Q _16755_/C _16723_/X vssd1 vssd1 vccd1 vccd1 _16752_/Y sky130_fd_sc_hd__a21oi_1
X_19540_ _19540_/CLK _19540_/D vssd1 vssd1 vccd1 vccd1 _19540_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_171_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13964_ _18618_/Q _13676_/X _13972_/S vssd1 vssd1 vccd1 vccd1 _13965_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15703_ _15811_/A _18444_/Q vssd1 vssd1 vccd1 vccd1 _15703_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11374__S1 _09957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ _19348_/Q _12864_/X _12756_/A _19538_/Q _12914_/X vssd1 vssd1 vccd1 vccd1
+ _12915_/X sky130_fd_sc_hd__a221o_1
XFILLER_47_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19471_ _19565_/CLK _19471_/D vssd1 vssd1 vccd1 vccd1 _19471_/Q sky130_fd_sc_hd__dfxtp_1
X_16683_ _16783_/A vssd1 vssd1 vccd1 vccd1 _16731_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13895_ _13895_/A vssd1 vssd1 vccd1 vccd1 _18587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15404__S _15406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15634_ _15634_/A vssd1 vssd1 vccd1 vccd1 _19309_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13713__A _15276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18422_ _18340_/A _18413_/X _18414_/X _18421_/Y vssd1 vssd1 vccd1 vccd1 _18423_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12846_ _12995_/A vssd1 vssd1 vccd1 vccd1 _12846_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11126__S1 _11065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _18353_/A vssd1 vssd1 vccd1 vccd1 _20021_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15565_ _15565_/A vssd1 vssd1 vccd1 vccd1 _19278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _13342_/A vssd1 vssd1 vccd1 vccd1 _12777_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17304_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17313_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _13767_/X _18837_/Q _14524_/S vssd1 vssd1 vccd1 vccd1 _14517_/A sky130_fd_sc_hd__mux2_1
X_18284_ _19994_/Q _12825_/X _18283_/X _17243_/X vssd1 vssd1 vccd1 vccd1 _19994_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ _12604_/A _17391_/A _12604_/B vssd1 vssd1 vccd1 vccd1 _11733_/B sky130_fd_sc_hd__or3_1
X_15496_ _19248_/Q _15270_/X _15500_/S vssd1 vssd1 vccd1 vccd1 _15497_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13859__S _13867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17235_ _15822_/X _17229_/X _17234_/X _17232_/X vssd1 vssd1 vccd1 vccd1 _19844_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14447_ _18818_/Q _14446_/X _14450_/S vssd1 vssd1 vccd1 vccd1 _14448_/A sky130_fd_sc_hd__mux2_1
X_11659_ _17394_/A _12664_/A vssd1 vssd1 vccd1 vccd1 _17391_/B sky130_fd_sc_hd__nand2_4
XFILLER_174_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18116__C1 _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17166_ _17166_/A vssd1 vssd1 vccd1 vccd1 _17166_/Y sky130_fd_sc_hd__inv_2
X_14378_ _14378_/A vssd1 vssd1 vccd1 vccd1 _18796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16117_ _13433_/X _19476_/Q _16117_/S vssd1 vssd1 vccd1 vccd1 _16118_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13329_ input10/X _13303_/X _13306_/X vssd1 vssd1 vccd1 vccd1 _13329_/X sky130_fd_sc_hd__a21o_1
X_17097_ _17122_/A _17097_/B _17097_/C vssd1 vssd1 vccd1 vccd1 _19794_/D sky130_fd_sc_hd__nor3_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_134_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19391_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_170_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16048_ _13453_/X _19445_/Q _16056_/S vssd1 vssd1 vccd1 vccd1 _16049_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15375__A _15443_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19807_ _19859_/CLK _19807_/D vssd1 vssd1 vccd1 vccd1 _19807_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_149_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19804_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10190__A1 _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17999_ _17725_/A _18000_/B _17998_/Y _17722_/A vssd1 vssd1 vccd1 vccd1 _18002_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12511__B _19605_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12467__A0 _12463_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19738_ _19852_/CLK _19738_/D vssd1 vssd1 vccd1 vccd1 _19738_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10312__A _10312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_145_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11365__S1 _10691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12524__A2_N _12667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19669_ _19671_/CLK _19669_/D vssd1 vssd1 vccd1 vccd1 _19669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09422_ _17815_/A vssd1 vssd1 vccd1 vccd1 _11625_/B sky130_fd_sc_hd__buf_2
XFILLER_25_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09353_ _19882_/Q _09345_/X _11877_/A _09352_/X vssd1 vssd1 vccd1 vccd1 _09354_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_52_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17158__B1 _17123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09284_ _19997_/Q vssd1 vssd1 vccd1 vccd1 _18293_/A sky130_fd_sc_hd__clkinv_4
XFILLER_138_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17749__B _17749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16145__S _16145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10628__S0 _10678_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__A _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15984__S _15984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12942__A1 _11135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10800__S0 _10073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10961_ _09611_/A _10951_/X _10960_/X _09619_/A _19900_/Q vssd1 vssd1 vccd1 vccd1
+ _10961_/X sky130_fd_sc_hd__a32o_4
XFILLER_141_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ _12700_/A _12700_/B vssd1 vssd1 vccd1 vccd1 _17247_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13680_ _15251_/A vssd1 vssd1 vccd1 vccd1 _14628_/A sky130_fd_sc_hd__buf_2
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10892_ _11002_/A vssd1 vssd1 vccd1 vccd1 _11114_/S sky130_fd_sc_hd__buf_4
XFILLER_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12631_ _12637_/A _12631_/B vssd1 vssd1 vccd1 vccd1 _12631_/Y sky130_fd_sc_hd__nor2_4
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15350_ _19183_/Q _15267_/X _15356_/S vssd1 vssd1 vccd1 vccd1 _15351_/A sky130_fd_sc_hd__mux2_1
X_12562_ _12559_/Y _12561_/X _12562_/S vssd1 vssd1 vccd1 vccd1 _12562_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ _14301_/A vssd1 vssd1 vccd1 vccd1 _18763_/D sky130_fd_sc_hd__clkbuf_1
X_11513_ _11506_/Y _11508_/Y _11510_/Y _11512_/Y _10063_/A vssd1 vssd1 vccd1 vccd1
+ _11513_/X sky130_fd_sc_hd__o221a_1
X_15281_ _19155_/Q _15279_/X hold9/X vssd1 vssd1 vccd1 vccd1 _15282_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12493_ _19843_/Q _12491_/B _12492_/Y vssd1 vssd1 vccd1 vccd1 _12494_/B sky130_fd_sc_hd__o21a_1
X_17020_ _19763_/Q vssd1 vssd1 vccd1 vccd1 _17027_/C sky130_fd_sc_hd__clkbuf_1
X_14232_ _14232_/A vssd1 vssd1 vccd1 vccd1 _18733_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10619__S0 _10617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11444_ _10632_/A _11441_/X _11443_/X _09577_/A vssd1 vssd1 vccd1 vccd1 _11444_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_51_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19503_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11736__A2 _12631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14163_ _13764_/X _18703_/Q _14163_/S vssd1 vssd1 vccd1 vccd1 _14164_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10095__S1 _10691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11375_ _11371_/X _11373_/X _11374_/X _10732_/A _09964_/X vssd1 vssd1 vccd1 vccd1
+ _11375_/X sky130_fd_sc_hd__o221a_1
XANTENNA__18270__S _18273_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11292__S0 _10977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13114_ _13115_/A _13132_/C vssd1 vssd1 vccd1 vccd1 _13114_/X sky130_fd_sc_hd__or2_1
X_10326_ _10534_/A vssd1 vssd1 vccd1 vccd1 _10326_/X sky130_fd_sc_hd__buf_2
XFILLER_124_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18971_ _19727_/CLK _18971_/D vssd1 vssd1 vccd1 vccd1 _18971_/Q sky130_fd_sc_hd__dfxtp_1
X_14094_ _18674_/Q _13643_/X _14098_/S vssd1 vssd1 vccd1 vccd1 _14095_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output161_A _12519_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_66_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19574_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _19740_/Q _12912_/X _13044_/X _12917_/X vssd1 vssd1 vccd1 vccd1 _13045_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _17760_/X _17762_/X _17922_/S vssd1 vssd1 vccd1 vccd1 _17922_/X sky130_fd_sc_hd__mux2_1
X_10257_ _18656_/Q _19247_/Q _19409_/Q _18624_/Q _09904_/S _10151_/A vssd1 vssd1 vccd1
+ vccd1 _10257_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10188_ _10188_/A _10188_/B vssd1 vssd1 vccd1 vccd1 _10188_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17853_ _17853_/A _17853_/B vssd1 vssd1 vccd1 vccd1 _17853_/X sky130_fd_sc_hd__or2_1
XFILLER_79_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17903__A_N _17899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16804_ _19991_/Q _19990_/Q _19989_/Q vssd1 vssd1 vccd1 vccd1 _16807_/B sky130_fd_sc_hd__nand3b_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14996_ _19036_/Q _14379_/X _15000_/S vssd1 vssd1 vccd1 vccd1 _14997_/A sky130_fd_sc_hd__mux2_1
X_17784_ _17729_/A _17783_/X _17719_/X vssd1 vssd1 vccd1 vccd1 _18050_/B sky130_fd_sc_hd__o21ba_1
X_19523_ _19542_/CLK _19523_/D vssd1 vssd1 vccd1 vccd1 _19523_/Q sky130_fd_sc_hd__dfxtp_2
X_16735_ _16898_/A vssd1 vssd1 vccd1 vccd1 _16773_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13947_ _13947_/A vssd1 vssd1 vccd1 vccd1 _18610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19454_ _19666_/CLK _19454_/D vssd1 vssd1 vccd1 vccd1 _19454_/Q sky130_fd_sc_hd__dfxtp_1
X_16666_ _19663_/Q _16663_/B _16665_/Y vssd1 vssd1 vccd1 vccd1 _19663_/D sky130_fd_sc_hd__o21a_1
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13878_ _13780_/X _18580_/Q _13878_/S vssd1 vssd1 vccd1 vccd1 _13879_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15617_ _15617_/A vssd1 vssd1 vccd1 vccd1 _19301_/D sky130_fd_sc_hd__clkbuf_1
X_18405_ _18409_/A _18405_/B vssd1 vssd1 vccd1 vccd1 _20038_/D sky130_fd_sc_hd__nor2_1
XFILLER_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12829_ _12856_/A vssd1 vssd1 vccd1 vccd1 _12829_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19385_ _19481_/CLK _19385_/D vssd1 vssd1 vccd1 vccd1 _19385_/Q sky130_fd_sc_hd__dfxtp_1
X_16597_ _19639_/Q _19638_/Q _16597_/C vssd1 vssd1 vccd1 vccd1 _16600_/B sky130_fd_sc_hd__and3_1
XFILLER_43_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15548_ _19271_/Q _15241_/X _15550_/S vssd1 vssd1 vccd1 vccd1 _15549_/A sky130_fd_sc_hd__mux2_1
X_18336_ _18336_/A _18349_/B vssd1 vssd1 vccd1 vccd1 _18336_/X sky130_fd_sc_hd__or2_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12621__B1 _12395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18267_ _18267_/A vssd1 vssd1 vccd1 vccd1 _19987_/D sky130_fd_sc_hd__clkbuf_1
X_15479_ _15479_/A vssd1 vssd1 vccd1 vccd1 _19240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19986_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13177__A1 _13060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17218_ _19839_/Q _17226_/B vssd1 vssd1 vccd1 vccd1 _17218_/X sky130_fd_sc_hd__or2_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18198_ _18198_/A _18198_/B vssd1 vssd1 vccd1 vccd1 _18255_/A sky130_fd_sc_hd__nor2_4
XANTENNA__11188__B1 _09752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12924__A1 _18461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_71_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17149_ _17149_/A _17346_/B _17149_/C vssd1 vssd1 vccd1 vccd1 _17229_/A sky130_fd_sc_hd__or3_2
XANTENNA__10086__S1 _10691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10307__A _10307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09971_ _18789_/Q _19060_/Q _19284_/Q _19028_/Q _10735_/S _09970_/X vssd1 vssd1 vccd1
+ vccd1 _09971_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10163__A1 _09569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13101__B2 _19519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10977__A _10977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13353__A _13353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _16808_/D _12820_/B vssd1 vssd1 vccd1 vccd1 _11952_/C sky130_fd_sc_hd__nor2_2
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14883__S _14889_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09336_ _16808_/A _16808_/B vssd1 vssd1 vccd1 vccd1 _09336_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12612__A0 _19988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _17325_/A _11684_/A _09265_/X _09266_/X vssd1 vssd1 vccd1 vccd1 _11622_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11601__A _11601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09198_ _20034_/Q vssd1 vssd1 vccd1 vccd1 _09272_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12915__B2 _19538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17854__A1 _17976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ _11582_/A vssd1 vssd1 vccd1 vccd1 _11160_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10111_ _10910_/A vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__buf_2
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11091_ _11091_/A vssd1 vssd1 vccd1 vccd1 _11170_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14123__S _14131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12432__A _12432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10042_ _18789_/Q _19060_/Q _19284_/Q _19028_/Q _10700_/S _11496_/A vssd1 vssd1 vccd1
+ vccd1 _10042_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14850_ _14580_/X _18971_/Q _14856_/S vssd1 vssd1 vccd1 vccd1 _14851_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13801_ _13799_/X _18554_/Q _13813_/S vssd1 vssd1 vccd1 vccd1 _13802_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09741__A _09741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11990__B _17772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A io_dbus_rdata[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14781_ _14781_/A vssd1 vssd1 vccd1 vccd1 _18944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11993_ _19965_/Q _11355_/A _12077_/S vssd1 vssd1 vccd1 vccd1 _17457_/A sky130_fd_sc_hd__mux2_2
XANTENNA__09847__B2 _19918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17909__A2 _17971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ _19614_/Q _19613_/Q _19612_/Q _16520_/D vssd1 vssd1 vccd1 vccd1 _16529_/D
+ sky130_fd_sc_hd__and4_1
X_13732_ _18535_/Q _13731_/X _13736_/S vssd1 vssd1 vccd1 vccd1 _13733_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10944_ _19105_/Q _18871_/Q _19553_/Q _19201_/Q _11305_/S _10943_/X vssd1 vssd1 vccd1
+ vccd1 _10944_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16451_ _18365_/A vssd1 vssd1 vccd1 vccd1 _18412_/A sky130_fd_sc_hd__clkbuf_4
X_13663_ _15238_/A vssd1 vssd1 vccd1 vccd1 _14615_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14793__S _14797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10875_ _10875_/A vssd1 vssd1 vccd1 vccd1 _10875_/X sky130_fd_sc_hd__buf_2
XFILLER_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15402_ _14615_/X _19206_/Q _15406_/S vssd1 vssd1 vccd1 vccd1 _15403_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ _19288_/CLK _19170_/D vssd1 vssd1 vccd1 vccd1 _19170_/Q sky130_fd_sc_hd__dfxtp_1
X_12614_ _18118_/B _12614_/B vssd1 vssd1 vccd1 vccd1 _12615_/B sky130_fd_sc_hd__or2_1
X_16382_ _13089_/X _19550_/Q _16382_/S vssd1 vssd1 vccd1 vccd1 _16383_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13594_ _13594_/A vssd1 vssd1 vccd1 vccd1 _18504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18121_ _18121_/A _18121_/B vssd1 vssd1 vccd1 vccd1 _18121_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15333_ _15333_/A vssd1 vssd1 vccd1 vccd1 _19175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12545_ _19845_/Q _17234_/A _12545_/C vssd1 vssd1 vccd1 vccd1 _12564_/B sky130_fd_sc_hd__and3_1
XANTENNA__10826__S _10826_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18052_ _19917_/Q _18051_/X _18085_/S vssd1 vssd1 vccd1 vccd1 _18053_/A sky130_fd_sc_hd__mux2_1
X_15264_ hold10/A vssd1 vssd1 vccd1 vccd1 _15277_/S sky130_fd_sc_hd__buf_2
X_12476_ _12473_/X _12665_/B _12474_/X _12475_/X vssd1 vssd1 vccd1 vccd1 _18068_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_17003_ _19758_/Q _17005_/C _17003_/C vssd1 vssd1 vccd1 vccd1 _17004_/C sky130_fd_sc_hd__and3_1
XANTENNA__11709__A2 _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ _14215_/A vssd1 vssd1 vccd1 vccd1 _18726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11427_ _11438_/A _11427_/B vssd1 vssd1 vccd1 vccd1 _11427_/X sky130_fd_sc_hd__or2_1
X_15195_ _19129_/Q vssd1 vssd1 vccd1 vccd1 _15196_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_153_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output86_A _12414_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ _18698_/Q _13743_/X _14146_/S vssd1 vssd1 vccd1 vccd1 _14147_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11358_ _11578_/B _11579_/A _11579_/B vssd1 vssd1 vccd1 vccd1 _11575_/C sky130_fd_sc_hd__nand3_1
XANTENNA__11657__S _11657_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15129__S _15131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ _09820_/A _10299_/X _10304_/X _10308_/X _09588_/A vssd1 vssd1 vccd1 vccd1
+ _10309_/X sky130_fd_sc_hd__a221o_1
X_18954_ _19504_/CLK _18954_/D vssd1 vssd1 vccd1 vccd1 _18954_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14033__S _14035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14077_ _14133_/A vssd1 vssd1 vccd1 vccd1 _14146_/S sky130_fd_sc_hd__buf_6
X_11289_ _10920_/A _11279_/Y _11284_/X _11288_/Y _09735_/A vssd1 vssd1 vccd1 vccd1
+ _11289_/X sky130_fd_sc_hd__o311a_2
XFILLER_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13028_ _19707_/Q _12989_/X _12990_/X _19675_/Q _13027_/X vssd1 vssd1 vccd1 vccd1
+ _13028_/X sky130_fd_sc_hd__a221o_1
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17905_ _17705_/X _17894_/X _17904_/X _17869_/X vssd1 vssd1 vccd1 vccd1 _17905_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18885_ _19314_/CLK _18885_/D vssd1 vssd1 vccd1 vccd1 _18885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13872__S _13878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17836_ _17836_/A vssd1 vssd1 vccd1 vccd1 _17836_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17767_ _17627_/X _17836_/A _17632_/X vssd1 vssd1 vccd1 vccd1 _17767_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA_clkbuf_leaf_18_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ _19029_/Q _14459_/X _14983_/S vssd1 vssd1 vccd1 vccd1 _14980_/A sky130_fd_sc_hd__mux2_1
X_19506_ _19508_/CLK _19506_/D vssd1 vssd1 vccd1 vccd1 _19506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16718_ _16728_/A _16718_/B _16718_/C vssd1 vssd1 vccd1 vccd1 _19677_/D sky130_fd_sc_hd__nor3_1
XFILLER_63_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17698_ _17702_/A _17702_/B vssd1 vssd1 vccd1 vccd1 _17698_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19437_ _19502_/CLK _19437_/D vssd1 vssd1 vccd1 vccd1 _19437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11405__B _12649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16649_ _16674_/A _16653_/C vssd1 vssd1 vccd1 vccd1 _16649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19368_ _19464_/CLK _19368_/D vssd1 vssd1 vccd1 vccd1 _19368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18319_ _18319_/A _18333_/B vssd1 vssd1 vccd1 vccd1 _18319_/X sky130_fd_sc_hd__or2_1
XFILLER_31_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12070__A1 _20028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16336__A1 _19538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19299_ _19299_/CLK _19299_/D vssd1 vssd1 vccd1 vccd1 _19299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10059__S1 _10037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11256__S0 _11003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10037__A _10037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09826__A _09826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11008__S0 _10893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09954_ _09954_/A vssd1 vssd1 vccd1 vccd1 _09955_/A sky130_fd_sc_hd__buf_2
X_09885_ _19509_/Q _18921_/Q _18958_/Q _18532_/Q _10175_/S _09858_/X vssd1 vssd1 vccd1
+ vccd1 _09885_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14878__S _14878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15563__A _15574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13389__A1 _15782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10660_ _11448_/A _10660_/B vssd1 vssd1 vccd1 vccd1 _10660_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09319_ _20045_/Q _09449_/B vssd1 vssd1 vccd1 vccd1 _09319_/X sky130_fd_sc_hd__or2_1
XFILLER_51_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12061__A1 _19524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ _18810_/Q _19145_/Q _10591_/S vssd1 vssd1 vccd1 vccd1 _10592_/B sky130_fd_sc_hd__mux2_1
XFILLER_139_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14118__S _14120_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10072__B1 _10606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12330_ _12330_/A _12330_/B vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__nor2_2
XFILLER_31_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13957__S _13961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11247__S0 _11057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ _19595_/Q vssd1 vssd1 vccd1 vccd1 _12263_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14000_ _16371_/A _14000_/B vssd1 vssd1 vccd1 vccd1 _15301_/A sky130_fd_sc_hd__nand2_4
XFILLER_141_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13561__A1 _13546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ _11221_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _11212_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11021__C1 _09975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09736__A _09736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12192_ _12188_/X _12651_/A _12191_/Y vssd1 vssd1 vccd1 vccd1 _12272_/D sky130_fd_sc_hd__a21o_1
XFILLER_122_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11143_ _10899_/A _11142_/X _10980_/X vssd1 vssd1 vccd1 vccd1 _11143_/Y sky130_fd_sc_hd__o21ai_1
Xoutput75 _12148_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[13] sky130_fd_sc_hd__buf_2
Xoutput86 _12414_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[23] sky130_fd_sc_hd__buf_2
Xoutput97 _11864_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[4] sky130_fd_sc_hd__buf_2
X_15951_ _19402_/Q _15244_/X _15951_/S vssd1 vssd1 vccd1 vccd1 _15952_/A sky130_fd_sc_hd__mux2_1
X_11074_ _19489_/Q _18901_/Q _18938_/Q _18512_/Q _11237_/S _10083_/A vssd1 vssd1 vccd1
+ vccd1 _11075_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11324__B1 _09341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14902_ _14902_/A vssd1 vssd1 vccd1 vccd1 _14911_/S sky130_fd_sc_hd__clkbuf_4
X_10025_ _11032_/A vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__clkbuf_2
X_15882_ _13293_/X _19371_/Q _15890_/S vssd1 vssd1 vccd1 vccd1 _15883_/A sky130_fd_sc_hd__mux2_1
X_18670_ _19487_/CLK _18670_/D vssd1 vssd1 vccd1 vccd1 _18670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16263__A0 _19525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17621_ _17560_/X _17595_/X _17598_/X _17620_/X vssd1 vssd1 vccd1 vccd1 _17621_/X
+ sky130_fd_sc_hd__o211a_1
X_14833_ _18313_/A _16811_/A _14831_/X _14832_/Y vssd1 vssd1 vccd1 vccd1 _18403_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output124_A _12661_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14089__A _14146_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14764_ _18937_/Q _14385_/X _14764_/S vssd1 vssd1 vccd1 vccd1 _14765_/A sky130_fd_sc_hd__mux2_1
X_17552_ _17524_/X _17530_/Y _17551_/X vssd1 vssd1 vccd1 vccd1 _17552_/X sky130_fd_sc_hd__a21o_1
X_11976_ _12027_/C _11976_/B _12029_/C _11976_/D vssd1 vssd1 vccd1 vccd1 _11976_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13715_ _18531_/Q _13714_/X _13715_/S vssd1 vssd1 vccd1 vccd1 _13716_/A sky130_fd_sc_hd__mux2_1
X_16503_ _19667_/Q _19669_/Q _19668_/Q _16673_/A vssd1 vssd1 vccd1 vccd1 _16684_/A
+ sky130_fd_sc_hd__and4_1
X_17483_ _17477_/X _17481_/X _17674_/S vssd1 vssd1 vccd1 vccd1 _17483_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10927_ _10051_/A _10926_/X _10056_/A vssd1 vssd1 vccd1 vccd1 _10927_/Y sky130_fd_sc_hd__o21ai_1
X_14695_ _14695_/A vssd1 vssd1 vccd1 vccd1 _18901_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19222_ _19286_/CLK _19222_/D vssd1 vssd1 vccd1 vccd1 _19222_/Q sky130_fd_sc_hd__dfxtp_1
X_16434_ _16434_/A vssd1 vssd1 vccd1 vccd1 _19573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13646_ _15225_/A vssd1 vssd1 vccd1 vccd1 _14602_/A sky130_fd_sc_hd__clkbuf_2
X_10858_ _11383_/A _10858_/B vssd1 vssd1 vccd1 vccd1 _10858_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19153_ _19906_/CLK _19153_/D vssd1 vssd1 vccd1 vccd1 _19153_/Q sky130_fd_sc_hd__dfxtp_1
X_16365_ _19544_/Q _16364_/X _16365_/S vssd1 vssd1 vccd1 vccd1 _16366_/A sky130_fd_sc_hd__mux2_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _13577_/A vssd1 vssd1 vccd1 vccd1 _13577_/X sky130_fd_sc_hd__clkbuf_4
X_10789_ _18645_/Q _19236_/Q _19398_/Q _18613_/Q _10751_/S _10112_/A vssd1 vssd1 vccd1
+ vccd1 _10790_/B sky130_fd_sc_hd__mux4_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11241__A _11250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15316_ _15316_/A vssd1 vssd1 vccd1 vccd1 _19167_/D sky130_fd_sc_hd__clkbuf_1
X_18104_ _17705_/X _17667_/B _18103_/Y vssd1 vssd1 vccd1 vccd1 _18104_/Y sky130_fd_sc_hd__o21ai_1
X_12528_ _19985_/Q _11537_/A _12528_/S vssd1 vssd1 vccd1 vccd1 _12529_/A sky130_fd_sc_hd__mux2_4
X_19084_ _19308_/CLK _19084_/D vssd1 vssd1 vccd1 vccd1 _19084_/Q sky130_fd_sc_hd__dfxtp_1
X_16296_ _12772_/B _16295_/Y _16318_/S vssd1 vssd1 vccd1 vccd1 _16296_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13867__S _13867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15247_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15247_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18035_ _17607_/X _18032_/Y _18034_/X _17543_/X vssd1 vssd1 vccd1 vccd1 _18035_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13001__A0 _09341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ _12459_/A vssd1 vssd1 vccd1 vccd1 _12482_/A sky130_fd_sc_hd__inv_2
XFILLER_173_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11158__A3 _11156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09646__A _10849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15178_ _15178_/A vssd1 vssd1 vccd1 vccd1 _19120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15829__A0 _19921_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14129_ _18690_/Q _13710_/X _14131_/S vssd1 vssd1 vccd1 vccd1 _14130_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19986_ _19986_/CLK _19986_/D vssd1 vssd1 vccd1 vccd1 _19986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18937_ _19487_/CLK _18937_/D vssd1 vssd1 vccd1 vccd1 _18937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14698__S _14702_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09670_ _10176_/A vssd1 vssd1 vccd1 vccd1 _09688_/A sky130_fd_sc_hd__buf_2
X_18868_ _18973_/CLK _18868_/D vssd1 vssd1 vccd1 vccd1 _18868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17819_ _17917_/A vssd1 vssd1 vccd1 vccd1 _18000_/A sky130_fd_sc_hd__buf_2
XFILLER_94_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18799_ _19486_/CLK _18799_/D vssd1 vssd1 vccd1 vccd1 _18799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09287__A2 _18293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16926__B _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12291__A1 _19532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16418__S _16426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_clock clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_15_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__11477__S0 _09967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17506__A0 _12529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09937_ _19508_/Q _18920_/Q _18957_/Q _18531_/Q _10173_/S _10271_/A vssd1 vssd1 vccd1
+ vccd1 _09937_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13806__A _14631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ _09868_/A _09868_/B vssd1 vssd1 vccd1 vccd1 _09868_/Y sky130_fd_sc_hd__nand2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _19480_/Q _19318_/Q _18727_/Q _18497_/Q _09726_/S _09730_/X vssd1 vssd1 vccd1
+ vccd1 _09800_/B sky130_fd_sc_hd__mux4_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_193_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11830_ _12420_/A vssd1 vssd1 vccd1 vccd1 _16268_/A sky130_fd_sc_hd__buf_2
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11762_/A _17429_/A vssd1 vssd1 vccd1 vccd1 _11763_/A sky130_fd_sc_hd__and2_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14637__A _14637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11760__S _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _19638_/Q _12839_/X _13499_/X vssd1 vssd1 vccd1 vccd1 _13500_/X sky130_fd_sc_hd__o21a_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _11448_/A _10709_/X _10711_/X vssd1 vssd1 vccd1 vccd1 _10712_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14831_/A vssd1 vssd1 vccd1 vccd1 _18414_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11704_/B _17395_/B _11692_/C vssd1 vssd1 vccd1 vccd1 _11693_/D sky130_fd_sc_hd__or3_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13431_ _13428_/Y _13429_/X _13430_/X _13554_/S _13351_/A vssd1 vssd1 vccd1 vccd1
+ _13432_/B sky130_fd_sc_hd__a221o_1
X_10643_ _10648_/A vssd1 vssd1 vccd1 vccd1 _10764_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11061__A _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16150_ _19490_/Q _14596_/A _16156_/S vssd1 vssd1 vccd1 vccd1 _16151_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ _19945_/Q _13362_/B vssd1 vssd1 vccd1 vccd1 _13397_/C sky130_fd_sc_hd__and2_1
X_10574_ _10574_/A _10574_/B vssd1 vssd1 vccd1 vccd1 _10574_/X sky130_fd_sc_hd__or2_1
XFILLER_167_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10596__A1 _11464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ _14631_/X _19083_/Q _15105_/S vssd1 vssd1 vccd1 vccd1 _15102_/A sky130_fd_sc_hd__mux2_1
X_12313_ _19533_/Q _12206_/X _12262_/X _12312_/X _12212_/X vssd1 vssd1 vccd1 vccd1
+ _12313_/X sky130_fd_sc_hd__o221a_1
XFILLER_166_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16081_ _16081_/A vssd1 vssd1 vccd1 vccd1 _19459_/D sky130_fd_sc_hd__clkbuf_1
X_13293_ _15247_/A vssd1 vssd1 vccd1 vccd1 _13293_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14372__A _14453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15032_ _15032_/A vssd1 vssd1 vccd1 vccd1 _19052_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13534__A1 _13533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12244_ _19833_/Q vssd1 vssd1 vccd1 vccd1 _17199_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19840_ _19876_/CLK _19840_/D vssd1 vssd1 vccd1 vccd1 _19840_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10443__S1 _10333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ _12175_/A vssd1 vssd1 vccd1 vccd1 _12175_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_123_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11000__S _11000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ _19488_/Q _18900_/Q _18937_/Q _18511_/Q _11004_/S _11065_/X vssd1 vssd1 vccd1
+ vccd1 _11127_/B sky130_fd_sc_hd__mux4_1
XFILLER_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19771_ _19817_/CLK _19771_/D vssd1 vssd1 vccd1 vccd1 _19771_/Q sky130_fd_sc_hd__dfxtp_1
X_16983_ _16993_/A _16983_/B _16983_/C vssd1 vssd1 vccd1 vccd1 _19752_/D sky130_fd_sc_hd__nor3_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16299__A _16299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18722_ _19476_/CLK _18722_/D vssd1 vssd1 vccd1 vccd1 _18722_/Q sky130_fd_sc_hd__dfxtp_1
X_11057_ _18672_/Q _19167_/Q _11057_/S vssd1 vssd1 vccd1 vccd1 _11057_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14311__S _14319_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15934_ _19394_/Q _15219_/X _15940_/S vssd1 vssd1 vccd1 vccd1 _15935_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12620__A _12620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16236__A0 _19520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10008_ _11225_/A vssd1 vssd1 vccd1 vccd1 _10910_/A sky130_fd_sc_hd__buf_2
X_18653_ _19406_/CLK _18653_/D vssd1 vssd1 vccd1 vccd1 _18653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15865_ _15865_/A vssd1 vssd1 vccd1 vccd1 _19363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11236__A _11236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15931__A _15988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17604_ _17662_/A _17604_/B vssd1 vssd1 vccd1 vccd1 _17694_/A sky130_fd_sc_hd__nand2_1
X_14816_ _14816_/A vssd1 vssd1 vccd1 vccd1 _18960_/D sky130_fd_sc_hd__clkbuf_1
X_18584_ _19559_/CLK _18584_/D vssd1 vssd1 vccd1 vccd1 _18584_/Q sky130_fd_sc_hd__dfxtp_1
X_15796_ _19916_/Q _12127_/A _15795_/Y vssd1 vssd1 vccd1 vccd1 _15796_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10808__C1 _09602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17535_ _17813_/A vssd1 vssd1 vccd1 vccd1 _17958_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14747_ _14747_/A vssd1 vssd1 vccd1 vccd1 _18925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11959_ _16226_/A _11957_/Y _11958_/X _11668_/X vssd1 vssd1 vccd1 vccd1 _11959_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18019__A _18019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14678_ _15589_/B vssd1 vssd1 vccd1 vccd1 _15445_/B sky130_fd_sc_hd__buf_4
X_17466_ _17463_/X _17465_/X _17573_/S vssd1 vssd1 vccd1 vccd1 _17466_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19205_ _19557_/CLK _19205_/D vssd1 vssd1 vccd1 vccd1 _19205_/Q sky130_fd_sc_hd__dfxtp_1
X_16417_ _16428_/A vssd1 vssd1 vccd1 vccd1 _16426_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13629_ _15212_/A vssd1 vssd1 vccd1 vccd1 _14589_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14981__S _14983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17858__A _18127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17397_ _17397_/A _17397_/B _17324_/X _17396_/X vssd1 vssd1 vccd1 vccd1 _17507_/S
+ sky130_fd_sc_hd__or4bb_4
XFILLER_121_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19136_ _19394_/CLK _19136_/D vssd1 vssd1 vccd1 vccd1 _19136_/Q sky130_fd_sc_hd__dfxtp_1
X_16348_ _16347_/A _16347_/C _16347_/B vssd1 vssd1 vccd1 vccd1 _16348_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10131__S0 _11449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__B1 _13591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19067_ _19389_/CLK _19067_/D vssd1 vssd1 vccd1 vccd1 _19067_/Q sky130_fd_sc_hd__dfxtp_1
X_16279_ _16213_/X _16278_/Y _15745_/Y vssd1 vssd1 vccd1 vccd1 _16279_/X sky130_fd_sc_hd__a21o_1
XFILLER_133_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18018_ _19914_/Q _17758_/X _18017_/X vssd1 vssd1 vccd1 vccd1 _19914_/D sky130_fd_sc_hd__o21a_1
XFILLER_172_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09824__S0 _10245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19969_ _19971_/CLK _19969_/D vssd1 vssd1 vccd1 vccd1 _19969_/Q sky130_fd_sc_hd__dfxtp_1
X_09722_ _09722_/A _09722_/B vssd1 vssd1 vccd1 vccd1 _09722_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16227__A0 _15688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09653_ _09653_/A vssd1 vssd1 vccd1 vccd1 _09723_/A sky130_fd_sc_hd__buf_2
XFILLER_27_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09584_ _11012_/A vssd1 vssd1 vccd1 vccd1 _11491_/A sky130_fd_sc_hd__buf_2
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17768__A _17772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16672__A _16672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10290_ _10466_/S vssd1 vssd1 vccd1 vccd1 _10465_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10425__S1 _10291_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14131__S _14131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13980_ _13980_/A vssd1 vssd1 vccd1 vccd1 _18625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10189__S0 _09881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12931_ _18437_/Q _12928_/X _17808_/S vssd1 vssd1 vccd1 vccd1 _12932_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09452__C _17339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16847__A _17073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13970__S _13972_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11056__A _11114_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _15650_/A vssd1 vssd1 vccd1 vccd1 _19316_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _13205_/A vssd1 vssd1 vccd1 vccd1 _13343_/A sky130_fd_sc_hd__buf_2
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14601_ _14601_/A vssd1 vssd1 vccd1 vccd1 _18871_/D sky130_fd_sc_hd__clkbuf_1
X_11813_ _11813_/A _11813_/B vssd1 vssd1 vccd1 vccd1 _11815_/A sky130_fd_sc_hd__nor2_2
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _19286_/Q _15289_/X _15583_/S vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__mux2_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12255__A1 _11562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16058__S _16060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12793_ _14479_/C vssd1 vssd1 vccd1 vccd1 _18198_/A sky130_fd_sc_hd__buf_2
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14532_/A vssd1 vssd1 vccd1 vccd1 _18844_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17376_/A vssd1 vssd1 vccd1 vccd1 _17355_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11744_ _11867_/A vssd1 vssd1 vccd1 vccd1 _12116_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15897__S _15901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14463_ _18823_/Q _14462_/X _14466_/S vssd1 vssd1 vccd1 vccd1 _14464_/A sky130_fd_sc_hd__mux2_1
X_17251_ _17251_/A vssd1 vssd1 vccd1 vccd1 _19850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18273__S _18273_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11675_ _11675_/A vssd1 vssd1 vccd1 vccd1 _12602_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ _13414_/A vssd1 vssd1 vccd1 vccd1 _18491_/D sky130_fd_sc_hd__clkbuf_1
X_16202_ _19514_/Q _14672_/A _16204_/S vssd1 vssd1 vccd1 vccd1 _16203_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10626_ _19370_/Q _18984_/Q _19434_/Q _18553_/Q _10625_/X _10604_/A vssd1 vssd1 vccd1
+ vccd1 _10627_/B sky130_fd_sc_hd__mux4_1
XFILLER_139_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17182_ _17197_/A vssd1 vssd1 vccd1 vccd1 _17182_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14394_ _14394_/A vssd1 vssd1 vccd1 vccd1 _18801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16133_ _16133_/A vssd1 vssd1 vccd1 vccd1 _19483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15198__A _18293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13345_ _19343_/Q _13154_/A _12704_/X _19533_/Q _13344_/X vssd1 vssd1 vccd1 vccd1
+ _13345_/X sky130_fd_sc_hd__a221o_1
X_10557_ _19113_/Q _18879_/Q _19561_/Q _19209_/Q _10560_/S _10461_/A vssd1 vssd1 vccd1
+ vccd1 _10558_/B sky130_fd_sc_hd__mux4_1
XFILLER_128_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14306__S _14308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16064_ _16132_/S vssd1 vssd1 vccd1 vccd1 _16073_/S sky130_fd_sc_hd__buf_2
XFILLER_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ _13276_/A _13276_/B vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__and2_4
X_10488_ _10548_/A _10487_/X _09695_/A vssd1 vssd1 vccd1 vccd1 _10488_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15015_ _15015_/A vssd1 vssd1 vccd1 vccd1 _19044_/D sky130_fd_sc_hd__clkbuf_1
X_12227_ _19973_/Q _10555_/A _12303_/S vssd1 vssd1 vccd1 vccd1 _12257_/A sky130_fd_sc_hd__mux2_4
XFILLER_64_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18302__A _18302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16457__B1 _16455_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19823_ _19859_/CLK _19823_/D vssd1 vssd1 vccd1 vccd1 _19823_/Q sky130_fd_sc_hd__dfxtp_1
X_12158_ _12855_/A _12156_/Y _12217_/C _11920_/X vssd1 vssd1 vccd1 vccd1 _12158_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11109_ _19102_/Q _18868_/Q _19550_/Q _19198_/Q _11000_/S _11065_/X vssd1 vssd1 vccd1
+ vccd1 _11110_/B sky130_fd_sc_hd__mux4_1
X_19754_ _19756_/CLK _19754_/D vssd1 vssd1 vccd1 vccd1 _19754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16966_ _16993_/A _16966_/B _16975_/D vssd1 vssd1 vccd1 vccd1 _19747_/D sky130_fd_sc_hd__nor3_1
X_12089_ _12366_/A _12084_/Y _12088_/X _11871_/X vssd1 vssd1 vccd1 vccd1 _12089_/X
+ sky130_fd_sc_hd__a211o_1
X_18705_ _19552_/CLK _18705_/D vssd1 vssd1 vccd1 vccd1 _18705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15917_ _15917_/A vssd1 vssd1 vccd1 vccd1 _19387_/D sky130_fd_sc_hd__clkbuf_1
X_19685_ _19720_/CLK _19685_/D vssd1 vssd1 vccd1 vccd1 _19685_/Q sky130_fd_sc_hd__dfxtp_1
X_16897_ _16897_/A _16897_/B _16906_/D vssd1 vssd1 vccd1 vccd1 _19730_/D sky130_fd_sc_hd__nor3_1
XFILLER_65_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18636_ _19485_/CLK _18636_/D vssd1 vssd1 vccd1 vccd1 _18636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15848_ _15916_/S vssd1 vssd1 vccd1 vccd1 _15857_/S sky130_fd_sc_hd__buf_2
XFILLER_92_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18567_ _19511_/CLK _18567_/D vssd1 vssd1 vccd1 vccd1 _18567_/Q sky130_fd_sc_hd__dfxtp_1
X_15779_ _15808_/A vssd1 vssd1 vccd1 vccd1 _15801_/S sky130_fd_sc_hd__buf_2
XANTENNA__17709__B1 _18019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17518_ _17721_/B _17542_/D vssd1 vssd1 vccd1 vccd1 _17549_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18498_ _19481_/CLK _18498_/D vssd1 vssd1 vccd1 vccd1 _18498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10352__S0 _10325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11413__B _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17449_ _17446_/X _17448_/X _17500_/S vssd1 vssd1 vccd1 vccd1 _17449_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15600__S _15600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18134__A0 _16219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19119_ _19570_/CLK _19119_/D vssd1 vssd1 vccd1 vccd1 _19119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_141_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14216__S _14218_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12525__A _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16431__S _16437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09834__A _10509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15047__S _15055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ _10043_/A vssd1 vssd1 vccd1 vccd1 _09706_/A sky130_fd_sc_hd__buf_2
XFILLER_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09636_ _10403_/A vssd1 vssd1 vccd1 vccd1 _10264_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_66_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09567_ _09567_/A vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14187__A _14209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11445__C1 _09603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _10872_/S vssd1 vssd1 vccd1 vccd1 _11481_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_168_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10343__S0 _10390_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10799__A1 _10775_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10894__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ _11460_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _11460_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10411_ _19912_/Q vssd1 vssd1 vccd1 vccd1 _10411_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11963__A2_N _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__S1 _10645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ _10652_/A _11390_/X _10655_/A vssd1 vssd1 vccd1 vccd1 _11391_/X sky130_fd_sc_hd__o21a_1
XFILLER_137_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16687__B1 _16667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13130_ _13130_/A vssd1 vssd1 vccd1 vccd1 _18475_/D sky130_fd_sc_hd__clkbuf_1
X_10342_ _10494_/S vssd1 vssd1 vccd1 vccd1 _10390_/S sky130_fd_sc_hd__buf_4
XFILLER_109_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13061_ _19927_/Q _19928_/Q vssd1 vssd1 vccd1 vccd1 _13094_/C sky130_fd_sc_hd__and2_1
X_10273_ _18784_/Q _19055_/Q _19279_/Q _19023_/Q _09926_/S _09858_/A vssd1 vssd1 vccd1
+ vccd1 _10273_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14650__A _14650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13370__C1 _13369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ _17176_/A _12034_/C vssd1 vssd1 vccd1 vccd1 _12012_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input48_A io_ibus_inst[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16820_ _16820_/A vssd1 vssd1 vccd1 vccd1 _17073_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16751_ _19687_/Q _16748_/C _16750_/Y vssd1 vssd1 vccd1 vccd1 _19687_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13963_ _13985_/A vssd1 vssd1 vccd1 vccd1 _13972_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_111_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12476__B2 _12475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16577__A _18281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18268__S _18268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15702_ _15702_/A vssd1 vssd1 vccd1 vccd1 _15811_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19470_ _19470_/CLK _19470_/D vssd1 vssd1 vccd1 vccd1 _19470_/Q sky130_fd_sc_hd__dfxtp_1
X_12914_ _12914_/A _12914_/B vssd1 vssd1 vccd1 vccd1 _12914_/X sky130_fd_sc_hd__and2_1
X_13894_ _13803_/X _18587_/Q _13900_/S vssd1 vssd1 vccd1 vccd1 _13895_/A sky130_fd_sc_hd__mux2_1
X_16682_ _16728_/A _16682_/B _16682_/C vssd1 vssd1 vccd1 vccd1 _19668_/D sky130_fd_sc_hd__nor3_1
XFILLER_47_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18421_ input53/X vssd1 vssd1 vccd1 vccd1 _18421_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15633_ _14637_/X _19309_/Q _15633_/S vssd1 vssd1 vccd1 vccd1 _15634_/A sky130_fd_sc_hd__mux2_1
X_12845_ _19861_/Q _12842_/X _12696_/A _19828_/Q _12844_/X vssd1 vssd1 vccd1 vccd1
+ _12845_/X sky130_fd_sc_hd__a221o_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11514__A _19923_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11436__C1 _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18352_ _18352_/A _18352_/B vssd1 vssd1 vccd1 vccd1 _18353_/A sky130_fd_sc_hd__or2_1
XANTENNA__12779__A2 _13527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _19278_/Q _15263_/X _15572_/S vssd1 vssd1 vccd1 vccd1 _15565_/A sky130_fd_sc_hd__mux2_1
X_12776_ _12776_/A vssd1 vssd1 vccd1 vccd1 _13342_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17303_/A vssd1 vssd1 vccd1 vccd1 _19874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11727_ _17378_/A _17325_/B _09265_/X vssd1 vssd1 vccd1 vccd1 _12604_/B sky130_fd_sc_hd__a21oi_1
X_14515_ _14572_/S vssd1 vssd1 vccd1 vccd1 _14524_/S sky130_fd_sc_hd__buf_2
X_15495_ _15495_/A vssd1 vssd1 vccd1 vccd1 _19247_/D sky130_fd_sc_hd__clkbuf_1
X_18283_ _18283_/A _18311_/B vssd1 vssd1 vccd1 vccd1 _18283_/X sky130_fd_sc_hd__or2_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14825__A _14831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15420__S _15428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17234_ _17234_/A _17240_/B vssd1 vssd1 vccd1 vccd1 _17234_/X sky130_fd_sc_hd__or2_1
XANTENNA__17201__A _18289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14446_ _14650_/A vssd1 vssd1 vccd1 vccd1 _14446_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11658_ _11658_/A vssd1 vssd1 vccd1 vccd1 _18930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18116__B1 _18115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10609_ _10609_/A vssd1 vssd1 vccd1 vccd1 _10609_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17165_ _15688_/X _17153_/X _17164_/X _17142_/X vssd1 vssd1 vccd1 vccd1 _19822_/D
+ sky130_fd_sc_hd__o211a_1
X_14377_ _18796_/Q _14376_/X _14386_/S vssd1 vssd1 vccd1 vccd1 _14378_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11589_ _11570_/Y _11572_/X _11576_/Y _11588_/X vssd1 vssd1 vccd1 vccd1 _11589_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_10_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16116_ _16116_/A vssd1 vssd1 vccd1 vccd1 _19475_/D sky130_fd_sc_hd__clkbuf_1
X_13328_ _13326_/X _13327_/X _13554_/S vssd1 vssd1 vccd1 vccd1 _13328_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17875__C1 _11657_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17096_ _17095_/A _17095_/C _19794_/Q vssd1 vssd1 vccd1 vccd1 _17097_/C sky130_fd_sc_hd__a21oi_1
XFILLER_142_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16047_ _16047_/A vssd1 vssd1 vccd1 vccd1 _16056_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_143_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13259_ _15241_/A vssd1 vssd1 vccd1 vccd1 _13259_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19806_ _20044_/CLK _19806_/D vssd1 vssd1 vccd1 vccd1 _19806_/Q sky130_fd_sc_hd__dfxtp_1
X_17998_ _17998_/A _17998_/B vssd1 vssd1 vccd1 vccd1 _17998_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19737_ _19737_/CLK _19737_/D vssd1 vssd1 vccd1 vccd1 _19737_/Q sky130_fd_sc_hd__dfxtp_4
X_16949_ _16957_/B _16946_/B _16860_/X vssd1 vssd1 vccd1 vccd1 _16949_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16487__A _16487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09332__B2 _09339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19668_ _19671_/CLK _19668_/D vssd1 vssd1 vccd1 vccd1 _19668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10573__S0 _11428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09421_ _17914_/A vssd1 vssd1 vccd1 vccd1 _17815_/A sky130_fd_sc_hd__clkbuf_2
X_18619_ _19049_/CLK _18619_/D vssd1 vssd1 vccd1 vccd1 _18619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19599_ _19601_/CLK _19599_/D vssd1 vssd1 vccd1 vccd1 _19599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09352_ _19894_/Q _09350_/A _19893_/Q vssd1 vssd1 vccd1 vccd1 _09352_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17158__A1 _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09283_ _20037_/Q vssd1 vssd1 vccd1 vccd1 _12935_/A sky130_fd_sc_hd__buf_4
XANTENNA__16426__S _16426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10628__S1 _09813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13785__S _13797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16161__S _16167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11902__B1 _12137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10800__S1 _10609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15505__S _15511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10960_ _09473_/A _10953_/X _10955_/X _10959_/X _09601_/A vssd1 vssd1 vccd1 vccd1
+ _10960_/X sky130_fd_sc_hd__a311o_2
XFILLER_55_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10564__S0 _11428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09619_ _09619_/A vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__buf_2
X_10891_ _18965_/Q vssd1 vssd1 vccd1 vccd1 _11002_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12630_ _12639_/A vssd1 vssd1 vccd1 vccd1 _12637_/A sky130_fd_sc_hd__buf_8
XFILLER_169_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12561_ _12561_/A _12581_/C vssd1 vssd1 vccd1 vccd1 _12561_/X sky130_fd_sc_hd__xor2_1
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11512_ _10039_/A _11511_/X _10655_/A vssd1 vssd1 vccd1 vccd1 _11512_/Y sky130_fd_sc_hd__o21ai_1
X_14300_ _18763_/Q _13608_/X _14308_/S vssd1 vssd1 vccd1 vccd1 _14301_/A sky130_fd_sc_hd__mux2_1
X_15280_ hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__buf_4
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12492_ _12492_/A _12545_/C vssd1 vssd1 vccd1 vccd1 _12492_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14231_ _13758_/X _18733_/Q _14235_/S vssd1 vssd1 vccd1 vccd1 _14232_/A sky130_fd_sc_hd__mux2_1
X_11443_ _11443_/A _11443_/B vssd1 vssd1 vccd1 vccd1 _11443_/X sky130_fd_sc_hd__or2_1
XANTENNA__10619__S1 _10682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14162_ _14162_/A vssd1 vssd1 vccd1 vccd1 _18702_/D sky130_fd_sc_hd__clkbuf_1
X_11374_ _19111_/Q _18877_/Q _19559_/Q _19207_/Q _11429_/S _09957_/X vssd1 vssd1 vccd1
+ vccd1 _11374_/X sky130_fd_sc_hd__mux4_2
XANTENNA__11292__S1 _10006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17321__B2 _11665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ _19931_/Q vssd1 vssd1 vccd1 vccd1 _13115_/A sky130_fd_sc_hd__clkbuf_2
X_10325_ _10337_/A vssd1 vssd1 vccd1 vccd1 _10325_/X sky130_fd_sc_hd__clkbuf_4
X_18970_ _19727_/CLK _18970_/D vssd1 vssd1 vccd1 vccd1 _18970_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16071__S _16073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14093_ _14093_/A vssd1 vssd1 vccd1 vccd1 _18673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _19852_/Q _12842_/X _12863_/X _19819_/Q _13043_/X vssd1 vssd1 vccd1 vccd1
+ _13044_/X sky130_fd_sc_hd__a221o_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17921_ _17921_/A vssd1 vssd1 vccd1 vccd1 _17921_/Y sky130_fd_sc_hd__clkinv_2
X_10256_ _10256_/A _10256_/B vssd1 vssd1 vccd1 vccd1 _10256_/X sky130_fd_sc_hd__or2_1
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output154_A _12348_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17852_ _17865_/S _17851_/X _17723_/X vssd1 vssd1 vccd1 vccd1 _17852_/Y sky130_fd_sc_hd__o21ai_1
X_10187_ _18658_/Q _19249_/Q _19411_/Q _18626_/Q _09723_/A _09868_/A vssd1 vssd1 vccd1
+ vccd1 _10188_/B sky130_fd_sc_hd__mux4_1
XFILLER_120_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10413__A _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16803_ _19706_/Q vssd1 vssd1 vccd1 vccd1 _16812_/A sky130_fd_sc_hd__inv_2
XFILLER_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17783_ _17845_/A _17782_/Y _17694_/X vssd1 vssd1 vccd1 vccd1 _17783_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14995_ _14995_/A vssd1 vssd1 vccd1 vccd1 _19035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15415__S _15417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19522_ _19837_/CLK _19522_/D vssd1 vssd1 vccd1 vccd1 _19522_/Q sky130_fd_sc_hd__dfxtp_2
X_16734_ _16737_/B _16737_/C _16733_/Y vssd1 vssd1 vccd1 vccd1 _19682_/D sky130_fd_sc_hd__o21a_1
X_13946_ _18610_/Q _13643_/X _13950_/S vssd1 vssd1 vccd1 vccd1 _13947_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19453_ _19726_/CLK _19453_/D vssd1 vssd1 vccd1 vccd1 _19453_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10559__S _10559_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16665_ _16674_/A _16670_/C vssd1 vssd1 vccd1 vccd1 _16665_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13877_ _13877_/A vssd1 vssd1 vccd1 vccd1 _18579_/D sky130_fd_sc_hd__clkbuf_1
X_18404_ _18404_/A vssd1 vssd1 vccd1 vccd1 _18409_/A sky130_fd_sc_hd__clkbuf_2
X_15616_ _14612_/X _19301_/Q _15622_/S vssd1 vssd1 vccd1 vccd1 _15617_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19384_ _19480_/CLK _19384_/D vssd1 vssd1 vccd1 vccd1 _19384_/Q sky130_fd_sc_hd__dfxtp_1
X_12828_ _16635_/A vssd1 vssd1 vccd1 vccd1 _16528_/A sky130_fd_sc_hd__clkbuf_4
X_16596_ _16783_/A vssd1 vssd1 vccd1 vccd1 _16631_/A sky130_fd_sc_hd__buf_2
XFILLER_90_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18335_ _18335_/A vssd1 vssd1 vccd1 vccd1 _18349_/B sky130_fd_sc_hd__clkbuf_1
X_15547_ _15547_/A vssd1 vssd1 vccd1 vccd1 _19270_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12621__A1 _12620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12759_ _13245_/A vssd1 vssd1 vccd1 vccd1 _12759_/X sky130_fd_sc_hd__buf_2
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18266_ _19987_/Q _19608_/Q _18268_/S vssd1 vssd1 vccd1 vccd1 _18267_/A sky130_fd_sc_hd__mux2_1
X_15478_ _19240_/Q _15244_/X _15478_/S vssd1 vssd1 vccd1 vccd1 _15479_/A sky130_fd_sc_hd__mux2_1
X_17217_ _17217_/A vssd1 vssd1 vccd1 vccd1 _17217_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14429_ _14429_/A vssd1 vssd1 vccd1 vccd1 _18812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18197_ _18197_/A vssd1 vssd1 vccd1 vccd1 _19956_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12075__A _19968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11188__A1 _09745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11188__B2 _11187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17148_ _17230_/A vssd1 vssd1 vccd1 vccd1 _17164_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15386__A _15443_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09970_ _09985_/A vssd1 vssd1 vccd1 vccd1 _09970_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17079_ _17079_/A _19788_/Q _17079_/C vssd1 vssd1 vccd1 vccd1 _17081_/B sky130_fd_sc_hd__and3_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11350__A1_N _11135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17106__A _17122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13634__A _14592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10320__C1 _09605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12860__A1 _16528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09404_ _19886_/Q _09404_/B vssd1 vssd1 vccd1 vccd1 _12820_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09335_ _20019_/Q vssd1 vssd1 vccd1 vccd1 _16808_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12612__A1 _12593_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09559__A _10296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _09426_/A _09266_/B vssd1 vssd1 vccd1 vccd1 _09266_/X sky130_fd_sc_hd__or2_2
XFILLER_138_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_180_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19620_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15995__S _16001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09197_ _20027_/Q _20026_/Q _20025_/Q vssd1 vssd1 vccd1 vccd1 _09275_/D sky130_fd_sc_hd__or3_2
XFILLER_147_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13809__A _14634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10110_ _10110_/A vssd1 vssd1 vccd1 vccd1 _10110_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11090_ _18576_/Q _18837_/Q _18736_/Q _19071_/Q _11147_/A _10007_/A vssd1 vssd1 vccd1
+ vccd1 _11090_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10041_ _10041_/A vssd1 vssd1 vccd1 vccd1 _11496_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13800_ _13832_/A vssd1 vssd1 vccd1 vccd1 _13813_/S sky130_fd_sc_hd__buf_2
XFILLER_63_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14780_ _18944_/Q _14408_/X _14786_/S vssd1 vssd1 vccd1 vccd1 _14781_/A sky130_fd_sc_hd__mux2_1
X_11992_ _17820_/A _11992_/B vssd1 vssd1 vccd1 vccd1 _11995_/A sky130_fd_sc_hd__xnor2_1
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13731_ _14666_/A vssd1 vssd1 vccd1 vccd1 _13731_/X sky130_fd_sc_hd__clkbuf_2
X_10943_ _11260_/A vssd1 vssd1 vccd1 vccd1 _10943_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_17_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_133_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19488_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16450_ _16678_/A vssd1 vssd1 vccd1 vccd1 _18365_/A sky130_fd_sc_hd__buf_4
X_13662_ _13662_/A vssd1 vssd1 vccd1 vccd1 _18518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10874_ _19106_/Q _18872_/Q _19554_/Q _19202_/Q _09983_/A _10084_/A vssd1 vssd1 vccd1
+ vccd1 _10874_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15401_ _15401_/A vssd1 vssd1 vccd1 vccd1 _19205_/D sky130_fd_sc_hd__clkbuf_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12613_ _18118_/B _12614_/B vssd1 vssd1 vccd1 vccd1 _18121_/A sky130_fd_sc_hd__nand2_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _13592_/Y _18504_/Q _13598_/S vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__mux2_1
X_16381_ _16381_/A vssd1 vssd1 vccd1 vccd1 _19549_/D sky130_fd_sc_hd__clkbuf_1
X_18120_ _18121_/A _17607_/X _17543_/X _18119_/X vssd1 vssd1 vccd1 vccd1 _18120_/X
+ sky130_fd_sc_hd__a211o_1
X_15332_ _19175_/Q _15241_/X _15334_/S vssd1 vssd1 vccd1 vccd1 _15333_/A sky130_fd_sc_hd__mux2_1
X_12544_ _17234_/A _12545_/C _19845_/Q vssd1 vssd1 vccd1 vccd1 _12544_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_148_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19671_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18051_ _17624_/X _18049_/X _18050_/X _18007_/A _12436_/Y vssd1 vssd1 vccd1 vccd1
+ _18051_/X sky130_fd_sc_hd__a32o_1
X_15263_ _15263_/A vssd1 vssd1 vccd1 vccd1 _15263_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12475_ _12475_/A _12475_/B vssd1 vssd1 vccd1 vccd1 _12475_/X sky130_fd_sc_hd__or2_2
XFILLER_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ _17005_/C _17003_/C _19758_/Q vssd1 vssd1 vccd1 vccd1 _17004_/B sky130_fd_sc_hd__a21oi_1
X_11426_ _19127_/Q _18893_/Q _19575_/Q _19223_/Q _10690_/X _11371_/A vssd1 vssd1 vccd1
+ vccd1 _11427_/B sky130_fd_sc_hd__mux4_1
X_14214_ _13838_/X _18726_/Q _14218_/S vssd1 vssd1 vccd1 vccd1 _14215_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15194_ _15194_/A vssd1 vssd1 vccd1 vccd1 _19128_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_188_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ _14145_/A vssd1 vssd1 vccd1 vccd1 _18697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13719__A _13719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ _11580_/A _11580_/B _11580_/C vssd1 vssd1 vccd1 vccd1 _11579_/B sky130_fd_sc_hd__a21o_1
XFILLER_125_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10308_ _10378_/A _10306_/X _10307_/X vssd1 vssd1 vccd1 vccd1 _10308_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output79_A _12260_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18953_ _19504_/CLK _18953_/D vssd1 vssd1 vccd1 vccd1 _18953_/Q sky130_fd_sc_hd__dfxtp_1
X_14076_ _15301_/A _16809_/C vssd1 vssd1 vccd1 vccd1 _14133_/A sky130_fd_sc_hd__nor2_4
X_11288_ _10986_/A _11285_/X _11287_/X vssd1 vssd1 vccd1 vccd1 _11288_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11017__S1 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13438__B _19950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13027_ _19611_/Q _12911_/X _13026_/X vssd1 vssd1 vccd1 vccd1 _13027_/X sky130_fd_sc_hd__o21a_1
X_17904_ _17995_/A _17904_/B _17904_/C _17904_/D vssd1 vssd1 vccd1 vccd1 _17904_/X
+ sky130_fd_sc_hd__or4_1
X_10239_ _10240_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _10241_/A sky130_fd_sc_hd__and2_1
X_18884_ _19311_/CLK _18884_/D vssd1 vssd1 vccd1 vccd1 _18884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17835_ _17971_/A _17828_/X _17834_/X _17796_/X vssd1 vssd1 vccd1 vccd1 _17835_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13454__A _13454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17766_ _17922_/S _17592_/X _17694_/X vssd1 vssd1 vccd1 vccd1 _17836_/A sky130_fd_sc_hd__o21ai_2
X_14978_ _14978_/A vssd1 vssd1 vccd1 vccd1 _19028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19505_ _19566_/CLK _19505_/D vssd1 vssd1 vccd1 vccd1 _19505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16717_ _19677_/Q _16717_/B _16717_/C vssd1 vssd1 vccd1 vccd1 _16718_/C sky130_fd_sc_hd__and3_1
XANTENNA__13173__B _13173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13929_ _13985_/A vssd1 vssd1 vccd1 vccd1 _13998_/S sky130_fd_sc_hd__buf_6
XFILLER_34_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17697_ _17785_/A vssd1 vssd1 vccd1 vccd1 _17697_/X sky130_fd_sc_hd__buf_2
XFILLER_35_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19436_ _19561_/CLK _19436_/D vssd1 vssd1 vccd1 vccd1 _19436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16648_ _16648_/A vssd1 vssd1 vccd1 vccd1 _16653_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19367_ _19557_/CLK _19367_/D vssd1 vssd1 vccd1 vccd1 _19367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16579_ _19633_/Q _16582_/C _16578_/Y vssd1 vssd1 vccd1 vccd1 _19633_/D sky130_fd_sc_hd__o21a_1
XFILLER_148_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18318_ _20006_/Q _18310_/X _18316_/X _18317_/X vssd1 vssd1 vccd1 vccd1 _20006_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19298_ _19552_/CLK _19298_/D vssd1 vssd1 vccd1 vccd1 _19298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11421__B _12661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18249_ _19979_/Q _19600_/Q _18253_/S vssd1 vssd1 vccd1 vccd1 _18250_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11256__S1 _11059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13629__A _15212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09953_ _10082_/A vssd1 vssd1 vccd1 vccd1 _09954_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11008__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09884_ _09884_/A vssd1 vssd1 vccd1 vccd1 _10233_/A sky130_fd_sc_hd__clkbuf_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10767__S0 _10644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_11_0_clock clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__09842__A _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10988__A _10988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15055__S _15055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19504_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14894__S _14900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19287_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09318_ _20044_/Q _20043_/Q _20042_/Q _20041_/Q vssd1 vssd1 vccd1 vccd1 _09449_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__11612__A _18138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ _10590_/A vssd1 vssd1 vccd1 vccd1 _10590_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10072__A1 _09515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09249_ _09249_/A vssd1 vssd1 vccd1 vccd1 _11724_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _12260_/A vssd1 vssd1 vccd1 vccd1 _12260_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_119_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11247__S1 _10943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11211_ _19359_/Q _18973_/Q _19423_/Q _18542_/Q _11083_/S _11164_/X vssd1 vssd1 vccd1
+ vccd1 _11212_/B sky130_fd_sc_hd__mux4_1
XFILLER_147_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14134__S _14142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12191_ _18311_/A _17334_/B _12190_/X vssd1 vssd1 vccd1 vccd1 _12191_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11142_ _19456_/Q _19294_/Q _18703_/Q _18473_/Q _11224_/S _11330_/A vssd1 vssd1 vccd1
+ vccd1 _11142_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput76 _12175_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[14] sky130_fd_sc_hd__buf_2
Xoutput87 _12436_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[24] sky130_fd_sc_hd__buf_2
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11059__A _11059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15754__A _15808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15950_ _15950_/A vssd1 vssd1 vccd1 vccd1 _19401_/D sky130_fd_sc_hd__clkbuf_1
X_11073_ _11125_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11073_/X sky130_fd_sc_hd__or2_1
Xoutput98 _11907_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10758__S0 _09647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14901_ _14901_/A vssd1 vssd1 vccd1 vccd1 _18994_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input30_A io_dbus_rdata[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _10024_/A vssd1 vssd1 vccd1 vccd1 _11032_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09752__A _09752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15881_ _15903_/A vssd1 vssd1 vccd1 vccd1 _15890_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17460__A0 _17832_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__S _11493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17620_ _17524_/X _17606_/Y _17617_/X _17619_/X vssd1 vssd1 vccd1 vccd1 _17620_/X
+ sky130_fd_sc_hd__a211o_1
X_14832_ input41/X vssd1 vssd1 vccd1 vccd1 _14832_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19981_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17551_ _12674_/B _17533_/X _17544_/X _17548_/X _17646_/A vssd1 vssd1 vccd1 vccd1
+ _17551_/X sky130_fd_sc_hd__a41o_1
X_14763_ _14763_/A vssd1 vssd1 vccd1 vccd1 _18936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11975_ _19583_/Q _11974_/A _11912_/B _19585_/Q vssd1 vssd1 vccd1 vccd1 _11976_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA_output117_A _12654_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16502_ _19665_/Q _19664_/Q _19666_/Q _16664_/A vssd1 vssd1 vccd1 vccd1 _16673_/A
+ sky130_fd_sc_hd__and4_1
X_13714_ _14653_/A vssd1 vssd1 vccd1 vccd1 _13714_/X sky130_fd_sc_hd__clkbuf_2
X_17482_ _17581_/S vssd1 vssd1 vccd1 vccd1 _17674_/S sky130_fd_sc_hd__clkbuf_2
X_10926_ _19492_/Q _18904_/Q _18941_/Q _18515_/Q _10909_/S _09660_/A vssd1 vssd1 vccd1
+ vccd1 _10926_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14694_ _18901_/Q _14388_/X _14702_/S vssd1 vssd1 vccd1 vccd1 _14695_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19221_ _19573_/CLK _19221_/D vssd1 vssd1 vccd1 vccd1 _19221_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10930__S0 _11493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16433_ _13487_/X _19573_/Q _16437_/S vssd1 vssd1 vccd1 vccd1 _16434_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10857_ _19365_/Q _18979_/Q _19429_/Q _18548_/Q _10777_/A _10010_/X vssd1 vssd1 vccd1
+ vccd1 _10858_/B sky130_fd_sc_hd__mux4_1
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13645_ _13645_/A vssd1 vssd1 vccd1 vccd1 _18514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19152_ _19906_/CLK _19152_/D vssd1 vssd1 vccd1 vccd1 _19152_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16364_ _15839_/X _16363_/Y _16364_/S vssd1 vssd1 vccd1 vccd1 _16364_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _09693_/A _10785_/Y _10787_/Y _09737_/A vssd1 vssd1 vccd1 vccd1 _10788_/X
+ sky130_fd_sc_hd__o31a_1
X_13576_ _16268_/A vssd1 vssd1 vccd1 vccd1 _16364_/S sky130_fd_sc_hd__buf_2
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _18100_/X _18102_/X _17619_/A vssd1 vssd1 vccd1 vccd1 _18103_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15315_ _19167_/Q _15215_/X _15323_/S vssd1 vssd1 vccd1 vccd1 _15316_/A sky130_fd_sc_hd__mux2_1
X_19083_ _19308_/CLK _19083_/D vssd1 vssd1 vccd1 vccd1 _19083_/Q sky130_fd_sc_hd__dfxtp_1
X_12527_ _18090_/A _12527_/B vssd1 vssd1 vccd1 vccd1 _12531_/A sky130_fd_sc_hd__xor2_1
XFILLER_157_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16295_ _16301_/A _16301_/C vssd1 vssd1 vccd1 vccd1 _16295_/Y sky130_fd_sc_hd__xnor2_1
X_18034_ _17815_/A _18036_/B _17998_/A _18033_/Y vssd1 vssd1 vccd1 vccd1 _18034_/X
+ sky130_fd_sc_hd__o211a_1
X_15246_ _15246_/A vssd1 vssd1 vccd1 vccd1 _19144_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09927__A _09927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12458_ _12458_/A _12458_/B vssd1 vssd1 vccd1 vccd1 _12482_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11409_ _11406_/Y _10728_/A _11407_/A vssd1 vssd1 vccd1 vccd1 _11409_/Y sky130_fd_sc_hd__a21oi_1
X_15177_ _19120_/Q vssd1 vssd1 vccd1 vccd1 _15178_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__14044__S _14046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12389_ _12335_/A _12335_/B _12358_/A _12356_/A _12330_/A vssd1 vssd1 vccd1 vccd1
+ _12390_/B sky130_fd_sc_hd__a221o_1
XFILLER_67_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15829__A1 _15828_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14128_ _14128_/A vssd1 vssd1 vccd1 vccd1 _18689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19985_ _19985_/CLK _19985_/D vssd1 vssd1 vccd1 vccd1 _19985_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17863__B _17866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14979__S _14983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10771__C1 _09717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13883__S _13889_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15664__A _15808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13304__A2 _13173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14059_ _14059_/A vssd1 vssd1 vccd1 vccd1 _14068_/S sky130_fd_sc_hd__buf_4
X_18936_ _19487_/CLK _18936_/D vssd1 vssd1 vccd1 vccd1 _18936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09662__A _09662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18867_ _18973_/CLK _18867_/D vssd1 vssd1 vccd1 vccd1 _18867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17818_ _17865_/S _17817_/X _17723_/X vssd1 vssd1 vccd1 vccd1 _17818_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10601__A _11411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18798_ _19487_/CLK _18798_/D vssd1 vssd1 vccd1 vccd1 _18798_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13068__B2 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17749_ _17749_/A _17749_/B vssd1 vssd1 vccd1 vccd1 _17749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16926__C _16926_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19419_ _19952_/CLK _19419_/D vssd1 vssd1 vccd1 vccd1 _19419_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15765__A0 _19911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17506__A1 _17702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11477__S1 _10074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__A1 _09979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10048__A _10048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14889__S _14889_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15574__A _15574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09936_ _09936_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _09936_/Y sky130_fd_sc_hd__nor2_1
XFILLER_104_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09572__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ _18820_/Q _19155_/Q _10218_/S vssd1 vssd1 vccd1 vccd1 _09868_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10514__C1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _09699_/A _09797_/X _09696_/X vssd1 vssd1 vccd1 vccd1 _09798_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_136_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14918__A _14974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15513__S _15515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11760_ _19959_/Q _11348_/A _11809_/A vssd1 vssd1 vccd1 vccd1 _17429_/A sky130_fd_sc_hd__mux2_2
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10912__S0 _11493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10711_ _09680_/A _10710_/X _10043_/X vssd1 vssd1 vccd1 vccd1 _10711_/X sky130_fd_sc_hd__o21a_1
XFILLER_41_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11691_ _09307_/B _09215_/A _09215_/B _11619_/A _09275_/X vssd1 vssd1 vccd1 vccd1
+ _11693_/B sky130_fd_sc_hd__o2111ai_2
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14129__S _14131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _11452_/A _10639_/Y _10641_/Y _10757_/A vssd1 vssd1 vccd1 vccd1 _10642_/X
+ sky130_fd_sc_hd__o211a_1
X_13430_ _19917_/Q _12921_/X _13430_/S vssd1 vssd1 vccd1 vccd1 _13430_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13968__S _13972_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__A1 _10757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ _16313_/A _13362_/B vssd1 vssd1 vccd1 vccd1 _13363_/B sky130_fd_sc_hd__nor2_1
X_10573_ _19467_/Q _19305_/Q _18714_/Q _18484_/Q _11428_/S _09814_/A vssd1 vssd1 vccd1
+ vccd1 _10574_/B sky130_fd_sc_hd__mux4_1
XFILLER_154_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15100_ _15100_/A vssd1 vssd1 vccd1 vccd1 _19082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09747__A _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12312_ _12309_/Y _12311_/X _12583_/S vssd1 vssd1 vccd1 vccd1 _12312_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16080_ _13149_/X _19459_/Q _16084_/S vssd1 vssd1 vccd1 vccd1 _16081_/A sky130_fd_sc_hd__mux2_1
X_13292_ _13292_/A _13292_/B vssd1 vssd1 vccd1 vccd1 _15247_/A sky130_fd_sc_hd__and2_4
XFILLER_170_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15031_ _19052_/Q _14430_/X _15033_/S vssd1 vssd1 vccd1 vccd1 _15032_/A sky130_fd_sc_hd__mux2_1
X_12243_ _11749_/B _12234_/Y _12241_/X _12242_/Y vssd1 vssd1 vccd1 vccd1 _12243_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10392__S _10392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10979__S0 _11224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12604__C _18009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ _12174_/A _12174_/B vssd1 vssd1 vccd1 vccd1 _12175_/A sky130_fd_sc_hd__xnor2_4
XFILLER_96_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11125_ _11125_/A _11125_/B vssd1 vssd1 vccd1 vccd1 _11125_/X sky130_fd_sc_hd__or2_1
X_19770_ _19817_/CLK _19770_/D vssd1 vssd1 vccd1 vccd1 _19770_/Q sky130_fd_sc_hd__dfxtp_1
X_16982_ _19752_/Q _19751_/Q _16984_/D vssd1 vssd1 vccd1 vccd1 _16983_/C sky130_fd_sc_hd__and3_1
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12901__A _18460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18721_ _19476_/CLK _18721_/D vssd1 vssd1 vccd1 vccd1 _18721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09482__A _11202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ _11114_/S vssd1 vssd1 vccd1 vccd1 _11057_/S sky130_fd_sc_hd__clkbuf_4
X_15933_ _15933_/A vssd1 vssd1 vccd1 vccd1 _19393_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10505__C1 _09740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12620__B _12620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10007_ _10007_/A vssd1 vssd1 vccd1 vccd1 _11225_/A sky130_fd_sc_hd__clkbuf_4
X_18652_ _19051_/CLK _18652_/D vssd1 vssd1 vccd1 vccd1 _18652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15864_ _13149_/X _19363_/Q _15868_/S vssd1 vssd1 vccd1 vccd1 _15865_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17603_ _17603_/A vssd1 vssd1 vccd1 vccd1 _17604_/B sky130_fd_sc_hd__inv_2
X_14815_ _18960_/Q _14459_/X _14819_/S vssd1 vssd1 vccd1 vccd1 _14816_/A sky130_fd_sc_hd__mux2_1
X_18583_ _19302_/CLK _18583_/D vssd1 vssd1 vccd1 vccd1 _18583_/Q sky130_fd_sc_hd__dfxtp_1
X_15795_ _15814_/A _17220_/A vssd1 vssd1 vccd1 vccd1 _15795_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17534_ _17538_/A _17534_/B _17538_/C vssd1 vssd1 vccd1 vccd1 _17813_/A sky130_fd_sc_hd__or3_1
XFILLER_45_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14746_ _18925_/Q _14465_/X _14746_/S vssd1 vssd1 vccd1 vccd1 _14747_/A sky130_fd_sc_hd__mux2_1
X_11958_ _19823_/Q _11958_/B vssd1 vssd1 vccd1 vccd1 _11958_/X sky130_fd_sc_hd__or2_1
XFILLER_91_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17465_ _17866_/B _18001_/B _17465_/S vssd1 vssd1 vccd1 vccd1 _17465_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _18803_/Q _19138_/Q _10909_/S vssd1 vssd1 vccd1 vccd1 _10910_/B sky130_fd_sc_hd__mux2_1
X_14677_ _14677_/A vssd1 vssd1 vccd1 vccd1 _18895_/D sky130_fd_sc_hd__clkbuf_1
X_11889_ _12032_/A vssd1 vssd1 vccd1 vccd1 _12214_/A sky130_fd_sc_hd__buf_2
X_19204_ _19204_/CLK _19204_/D vssd1 vssd1 vccd1 vccd1 _19204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16416_ _16416_/A vssd1 vssd1 vccd1 vccd1 _19565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13628_ _13628_/A vssd1 vssd1 vccd1 vccd1 _18510_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11459__S1 _10703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17396_ _11673_/A _17396_/B _17396_/C _17396_/D vssd1 vssd1 vccd1 vccd1 _17396_/X
+ sky130_fd_sc_hd__and4b_1
XANTENNA__09977__A1 _09989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19135_ _19201_/CLK _19135_/D vssd1 vssd1 vccd1 vccd1 _19135_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13878__S _13878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16347_ _16347_/A _16347_/B _16347_/C vssd1 vssd1 vccd1 vccd1 _16353_/B sky130_fd_sc_hd__or3_1
X_13559_ _13559_/A vssd1 vssd1 vccd1 vccd1 _18500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10131__S1 _10718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11784__A1 _19516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19066_ _19389_/CLK _19066_/D vssd1 vssd1 vccd1 vccd1 _19066_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09657__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ _16278_/A _16282_/C vssd1 vssd1 vccd1 vccd1 _16278_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_145_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18017_ _12362_/Y _18007_/X _18016_/X _17778_/X vssd1 vssd1 vccd1 vccd1 _18017_/X
+ sky130_fd_sc_hd__a211o_1
X_15229_ _19139_/Q _15228_/X _15229_/S vssd1 vssd1 vccd1 vccd1 _15230_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09824__S1 _09899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19968_ _19971_/CLK _19968_/D vssd1 vssd1 vccd1 vccd1 _19968_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09721_ _19129_/Q _18895_/Q _19577_/Q _19225_/Q _09655_/X _09788_/A vssd1 vssd1 vccd1
+ vccd1 _09722_/B sky130_fd_sc_hd__mux4_1
X_18919_ _19507_/CLK _18919_/D vssd1 vssd1 vccd1 vccd1 _18919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19899_ _19914_/CLK _19899_/D vssd1 vssd1 vccd1 vccd1 _19899_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09652_ _10270_/S vssd1 vssd1 vccd1 vccd1 _09653_/A sky130_fd_sc_hd__buf_4
XFILLER_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09583_ _11199_/A vssd1 vssd1 vccd1 vccd1 _11012_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16429__S _16437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13642__A _15222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17114__A _17122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17727__A1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17768__B _17772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13788__S _13797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10983__C1 _09736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13089__A _15212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09286__B _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10506__A _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10940__S _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12721__A _17247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09919_ _10156_/A _09916_/X _09918_/X _09580_/A vssd1 vssd1 vccd1 vccd1 _09919_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10189__S1 _10219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20039_ _20052_/CLK _20039_/D vssd1 vssd1 vccd1 vccd1 _20039_/Q sky130_fd_sc_hd__dfxtp_1
X_12930_ _18127_/A vssd1 vssd1 vccd1 vccd1 _17808_/S sky130_fd_sc_hd__buf_4
XFILLER_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _13204_/A vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11138__S0 _10017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14599_/X _18871_/Q _14606_/S vssd1 vssd1 vccd1 vccd1 _14601_/A sky130_fd_sc_hd__mux2_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11812_ _11812_/A _17431_/A vssd1 vssd1 vccd1 vccd1 _11813_/B sky130_fd_sc_hd__nor2_1
X_15580_ _15580_/A vssd1 vssd1 vccd1 vccd1 _19285_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12686_/Y _15764_/A _12791_/X vssd1 vssd1 vccd1 vccd1 _19807_/D sky130_fd_sc_hd__o21ai_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _13790_/X _18844_/Q _14535_/S vssd1 vssd1 vccd1 vccd1 _14532_/A sky130_fd_sc_hd__mux2_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _12029_/C _11976_/B vssd1 vssd1 vccd1 vccd1 _11867_/A sky130_fd_sc_hd__nand2_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _13572_/X _19850_/Q _17258_/S vssd1 vssd1 vccd1 vccd1 _17251_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14666_/A vssd1 vssd1 vccd1 vccd1 _14462_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11674_ _12595_/B _11729_/A _12596_/B vssd1 vssd1 vccd1 vccd1 _11693_/C sky130_fd_sc_hd__o21bai_1
XFILLER_169_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16201_ _16201_/A vssd1 vssd1 vccd1 vccd1 _19513_/D sky130_fd_sc_hd__clkbuf_1
X_13413_ _18491_/Q _13412_/X _13434_/S vssd1 vssd1 vccd1 vccd1 _13414_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10625_ _10826_/S vssd1 vssd1 vccd1 vccd1 _10625_/X sky130_fd_sc_hd__clkbuf_4
X_17181_ _15724_/X _17167_/X _17180_/X _17171_/X vssd1 vssd1 vccd1 vccd1 _19827_/D
+ sky130_fd_sc_hd__o211a_1
X_14393_ _18801_/Q _14392_/X _14402_/S vssd1 vssd1 vccd1 vccd1 _14394_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11310__S0 _11114_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12963__B1 _11411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16132_ _13557_/X _19483_/Q _16132_/S vssd1 vssd1 vccd1 vccd1 _16133_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15198__B _15198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10556_ _10556_/A _10556_/B vssd1 vssd1 vccd1 vccd1 _11565_/A sky130_fd_sc_hd__nor2_1
X_13344_ _19869_/Q _12913_/X _13343_/X _19836_/Q vssd1 vssd1 vccd1 vccd1 _13344_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16063_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16132_/S sky130_fd_sc_hd__buf_4
X_10487_ _19501_/Q _18913_/Q _18950_/Q _18524_/Q _10390_/S _10333_/A vssd1 vssd1 vccd1
+ vccd1 _10487_/X sky130_fd_sc_hd__mux4_1
X_13275_ _13337_/A _13270_/X _13274_/Y _13324_/A vssd1 vssd1 vccd1 vccd1 _13276_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_136_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15014_ _19044_/Q _14404_/X _15022_/S vssd1 vssd1 vccd1 vccd1 _15015_/A sky130_fd_sc_hd__mux2_1
X_12226_ _17945_/B _12226_/B vssd1 vssd1 vccd1 vccd1 _12228_/A sky130_fd_sc_hd__xnor2_4
XFILLER_151_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12191__A1 _18311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19822_ _19859_/CLK _19822_/D vssd1 vssd1 vccd1 vccd1 _19822_/Q sky130_fd_sc_hd__dfxtp_2
X_12157_ _19830_/Q _19829_/Q _12157_/C vssd1 vssd1 vccd1 vccd1 _12217_/C sky130_fd_sc_hd__and3_1
XFILLER_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12631__A _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11108_ _09745_/A _11095_/Y _11106_/X _09752_/A _11107_/Y vssd1 vssd1 vccd1 vccd1
+ _12637_/B sky130_fd_sc_hd__o32a_4
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19753_ _19756_/CLK _19753_/D vssd1 vssd1 vccd1 vccd1 _19753_/Q sky130_fd_sc_hd__dfxtp_1
X_16965_ _19747_/Q _19746_/Q _16965_/C _16965_/D vssd1 vssd1 vccd1 vccd1 _16975_/D
+ sky130_fd_sc_hd__and4_1
X_12088_ _12119_/B _12088_/B _12153_/A _12088_/D vssd1 vssd1 vccd1 vccd1 _12088_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_110_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11377__S0 _10073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15942__A _15988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18704_ _19551_/CLK _18704_/D vssd1 vssd1 vccd1 vccd1 _18704_/Q sky130_fd_sc_hd__dfxtp_1
X_11039_ _11046_/A _11034_/X _11038_/X vssd1 vssd1 vccd1 vccd1 _11039_/Y sky130_fd_sc_hd__o21ai_1
X_15916_ _13557_/X _19387_/Q _15916_/S vssd1 vssd1 vccd1 vccd1 _15917_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10151__A _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19684_ _19720_/CLK _19684_/D vssd1 vssd1 vccd1 vccd1 _19684_/Q sky130_fd_sc_hd__dfxtp_1
X_16896_ _19730_/Q _19729_/Q _19728_/Q _16896_/D vssd1 vssd1 vccd1 vccd1 _16906_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09940__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18635_ _19258_/CLK _18635_/D vssd1 vssd1 vccd1 vccd1 _18635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15847_ _15903_/A vssd1 vssd1 vccd1 vccd1 _15916_/S sky130_fd_sc_hd__buf_4
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18566_ _19317_/CLK _18566_/D vssd1 vssd1 vccd1 vccd1 _18566_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _19913_/Q _15708_/X _16315_/B vssd1 vssd1 vccd1 vccd1 _15778_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17709__A1 _11816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17517_ _17545_/B vssd1 vssd1 vccd1 vccd1 _17721_/B sky130_fd_sc_hd__inv_2
X_14729_ _18917_/Q _14440_/X _14735_/S vssd1 vssd1 vccd1 vccd1 _14730_/A sky130_fd_sc_hd__mux2_1
X_18497_ _19480_/CLK _18497_/D vssd1 vssd1 vccd1 vccd1 _18497_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14992__S _15000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10352__S1 _10326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17448_ _17937_/A _17949_/A _17460_/S vssd1 vssd1 vccd1 vccd1 _17448_/X sky130_fd_sc_hd__mux2_1
X_17379_ _17379_/A _17379_/B _17379_/C _17379_/D vssd1 vssd1 vccd1 vccd1 _17392_/C
+ sky130_fd_sc_hd__or4_2
XANTENNA__18134__A1 _19960_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19118_ _19566_/CLK _19118_/D vssd1 vssd1 vccd1 vccd1 _19118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19049_ _19049_/CLK _19049_/D vssd1 vssd1 vccd1 vccd1 _19049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17808__S _17808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16948__A _19744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11157__A _19897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _09999_/A vssd1 vssd1 vccd1 vccd1 _10043_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09886__B1 _09696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09850__A _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09635_ _10500_/A vssd1 vssd1 vccd1 vccd1 _10403_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16159__S _16167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__A _19900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09566_ _09526_/X _09542_/X _09565_/X vssd1 vssd1 vccd1 vccd1 _09566_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09497_ _10937_/S vssd1 vssd1 vccd1 vccd1 _10872_/S sky130_fd_sc_hd__buf_2
XANTENNA__10343__S1 _10333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18125__A1 _12620_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ _10403_/Y _10405_/Y _10407_/Y _10409_/Y _09719_/A vssd1 vssd1 vccd1 vccd1
+ _10410_/X sky130_fd_sc_hd__o221a_1
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11390_ _18776_/Q _19047_/Q _19271_/Q _19015_/Q _10048_/A _10037_/A vssd1 vssd1 vccd1
+ vccd1 _11390_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10341_ _10589_/S vssd1 vssd1 vccd1 vccd1 _10494_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_152_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ _13351_/A vssd1 vssd1 vccd1 vccd1 _13060_/X sky130_fd_sc_hd__clkbuf_4
X_10272_ _09929_/X _10269_/Y _10271_/Y _10264_/A vssd1 vssd1 vccd1 vccd1 _10272_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12011_ _17176_/A _12034_/C vssd1 vssd1 vccd1 vccd1 _12011_/X sky130_fd_sc_hd__or2_1
XFILLER_105_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14142__S _14142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16858__A _16946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16750_ _16775_/A _16755_/C vssd1 vssd1 vccd1 vccd1 _16750_/Y sky130_fd_sc_hd__nor2_1
X_13962_ _13962_/A vssd1 vssd1 vccd1 vccd1 _18617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15701_ _18444_/Q _15701_/B vssd1 vssd1 vccd1 vccd1 _15701_/X sky130_fd_sc_hd__or2_1
XANTENNA__09760__A _12593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12913_ _12992_/A vssd1 vssd1 vccd1 vccd1 _12913_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16681_ _16680_/A _16680_/C _19668_/Q vssd1 vssd1 vccd1 vccd1 _16682_/C sky130_fd_sc_hd__a21oi_1
X_13893_ _13893_/A vssd1 vssd1 vccd1 vccd1 _18586_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16069__S _16073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18420_ _18426_/A _18420_/B vssd1 vssd1 vccd1 vccd1 _20047_/D sky130_fd_sc_hd__nor2_1
X_15632_ _15632_/A vssd1 vssd1 vccd1 vccd1 _19308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _19335_/Q _13245_/A _13099_/A _19525_/Q _12843_/X vssd1 vssd1 vccd1 vccd1
+ _12844_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _09328_/D _16811_/A _14825_/X input34/X vssd1 vssd1 vccd1 vccd1 _18352_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15574_/A vssd1 vssd1 vccd1 vccd1 _15572_/S sky130_fd_sc_hd__buf_2
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12989_/A vssd1 vssd1 vccd1 vccd1 _12775_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _15799_/Y _19874_/Q _17302_/S vssd1 vssd1 vccd1 vccd1 _17303_/A sky130_fd_sc_hd__mux2_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14514_ _14514_/A vssd1 vssd1 vccd1 vccd1 _18836_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _12606_/D _12946_/X _18281_/X _12825_/X vssd1 vssd1 vccd1 vccd1 _19993_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11726_ _17325_/A _17325_/B vssd1 vssd1 vccd1 vccd1 _12604_/A sky130_fd_sc_hd__nor2_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _19247_/Q _15267_/X _15500_/S vssd1 vssd1 vccd1 vccd1 _15495_/A sky130_fd_sc_hd__mux2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13189__A0 _19902_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17233_ _17228_/Y _17229_/X _17231_/X _17232_/X vssd1 vssd1 vccd1 vccd1 _19843_/D
+ sky130_fd_sc_hd__o211a_1
X_14445_ _14445_/A vssd1 vssd1 vccd1 vccd1 _18817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11657_ _11656_/X _17379_/A _11657_/S vssd1 vssd1 vccd1 vccd1 _11658_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14317__S _14319_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18116__A1 _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13221__S _13278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15002__A _15059_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12936__B1 _11302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10608_ _10824_/S vssd1 vssd1 vccd1 vccd1 _10608_/X sky130_fd_sc_hd__buf_4
XANTENNA__10098__S0 _11372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17164_ _19822_/Q _17164_/B vssd1 vssd1 vccd1 vccd1 _17164_/X sky130_fd_sc_hd__or2_1
XFILLER_167_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14376_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14376_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11588_ _11575_/Y _11577_/X _11578_/Y _11579_/Y _11587_/X vssd1 vssd1 vccd1 vccd1
+ _11588_/X sky130_fd_sc_hd__a221o_1
X_16115_ _13423_/X _19475_/Q _16117_/S vssd1 vssd1 vccd1 vccd1 _16116_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ _19911_/Q _12787_/B _13553_/S vssd1 vssd1 vccd1 vccd1 _13327_/X sky130_fd_sc_hd__mux2_1
X_10539_ _18779_/Q _19050_/Q _19274_/Q _19018_/Q _10533_/S _09665_/A vssd1 vssd1 vccd1
+ vccd1 _10539_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17095_ _17095_/A _19794_/Q _17095_/C vssd1 vssd1 vccd1 vccd1 _17097_/B sky130_fd_sc_hd__and3_1
X_16046_ _16046_/A vssd1 vssd1 vccd1 vccd1 _19444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13258_ _11656_/X _13256_/X _13257_/X vssd1 vssd1 vccd1 vccd1 _15241_/A sky130_fd_sc_hd__o21a_4
XFILLER_171_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12209_ _12338_/A _12338_/C vssd1 vssd1 vccd1 vccd1 _12209_/X sky130_fd_sc_hd__xor2_1
XFILLER_124_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13189_ _19902_/Q _15716_/B _13371_/A vssd1 vssd1 vccd1 vccd1 _13189_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19805_ _19805_/CLK _19805_/D vssd1 vssd1 vccd1 vccd1 _19805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14987__S _14987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17997_ _18001_/A _18001_/B _18077_/S vssd1 vssd1 vccd1 vccd1 _17998_/B sky130_fd_sc_hd__mux2_1
X_19736_ _19737_/CLK _19736_/D vssd1 vssd1 vccd1 vccd1 _19736_/Q sky130_fd_sc_hd__dfxtp_2
X_16948_ _19744_/Q vssd1 vssd1 vccd1 vccd1 _16957_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18052__A0 _19917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09963__S0 _10811_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16879_ _16921_/B _16883_/D _19724_/Q vssd1 vssd1 vccd1 vccd1 _16881_/B sky130_fd_sc_hd__a21oi_1
X_19667_ _19671_/CLK _19667_/D vssd1 vssd1 vccd1 vccd1 _19667_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_10_clock_A _19998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10573__S1 _09814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09420_ _09420_/A vssd1 vssd1 vccd1 vccd1 _17914_/A sky130_fd_sc_hd__clkbuf_2
X_18618_ _19049_/CLK _18618_/D vssd1 vssd1 vccd1 vccd1 _18618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19598_ _19601_/CLK _19598_/D vssd1 vssd1 vccd1 vccd1 _19598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09351_ _09349_/B _09347_/Y _13353_/A vssd1 vssd1 vccd1 vccd1 _11877_/A sky130_fd_sc_hd__a21o_1
X_18549_ _19430_/CLK _18549_/D vssd1 vssd1 vccd1 vccd1 _18549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09282_ _15198_/B _11640_/A vssd1 vssd1 vccd1 vccd1 _09282_/X sky130_fd_sc_hd__and2_1
XFILLER_100_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14227__S _14235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18107__A1 _19922_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11440__A _11440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15847__A _15903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16678__A _16678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14198__A _14209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10564__S1 _09814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09618_ _09618_/A vssd1 vssd1 vccd1 vccd1 _09619_/A sky130_fd_sc_hd__buf_2
XFILLER_83_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10890_ _19460_/Q _19298_/Q _18707_/Q _18477_/Q _09967_/A _09513_/A vssd1 vssd1 vccd1
+ vccd1 _10890_/X sky130_fd_sc_hd__mux4_1
X_09549_ _10294_/A vssd1 vssd1 vccd1 vccd1 _10368_/A sky130_fd_sc_hd__buf_2
XFILLER_34_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18346__A1 _17338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ _19607_/Q vssd1 vssd1 vccd1 vccd1 _12561_/A sky130_fd_sc_hd__buf_2
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _18665_/Q _19256_/Q _19418_/Q _18633_/Q _11384_/S _10105_/A vssd1 vssd1 vccd1
+ vccd1 _11511_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12491_ _19843_/Q _12491_/B vssd1 vssd1 vccd1 vccd1 _12545_/C sky130_fd_sc_hd__and2_1
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14230_ _14230_/A vssd1 vssd1 vccd1 vccd1 _18732_/D sky130_fd_sc_hd__clkbuf_1
X_11442_ _19481_/Q _19319_/Q _18728_/Q _18498_/Q _11372_/S _10813_/A vssd1 vssd1 vccd1
+ vccd1 _11443_/B sky130_fd_sc_hd__mux4_1
XFILLER_165_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11373_ _10825_/A _11372_/X _10613_/A vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14161_ _13761_/X _18702_/Q _14163_/S vssd1 vssd1 vccd1 vccd1 _14162_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10324_ _10544_/A vssd1 vssd1 vccd1 vccd1 _10436_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input60_A io_ibus_inst[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ _13112_/A vssd1 vssd1 vccd1 vccd1 _18474_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09755__A _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14092_ _18673_/Q _13639_/X _14098_/S vssd1 vssd1 vccd1 vccd1 _14093_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13277__A _15244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10255_ _19505_/Q _18917_/Q _18954_/Q _18528_/Q _09902_/S _09822_/A vssd1 vssd1 vccd1
+ vccd1 _10256_/B sky130_fd_sc_hd__mux4_1
X_13043_ _19326_/Q _12864_/X _12756_/A _19516_/Q _13042_/X vssd1 vssd1 vccd1 vccd1
+ _13043_/X sky130_fd_sc_hd__a221o_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17920_ _17533_/X _17912_/Y _17919_/X _18054_/A vssd1 vssd1 vccd1 vccd1 _17920_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17851_ _17853_/A _17853_/B vssd1 vssd1 vccd1 vccd1 _17851_/X sky130_fd_sc_hd__and2_1
X_10186_ _10188_/A _10185_/X _09696_/X vssd1 vssd1 vccd1 vccd1 _10186_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10413__B _12656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output147_A _16471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16802_ _19705_/Q _16799_/B _16801_/Y vssd1 vssd1 vccd1 vccd1 _19705_/D sky130_fd_sc_hd__o21a_1
X_17782_ _17782_/A vssd1 vssd1 vccd1 vccd1 _17782_/Y sky130_fd_sc_hd__inv_2
X_14994_ _19035_/Q _14376_/X _15000_/S vssd1 vssd1 vccd1 vccd1 _14995_/A sky130_fd_sc_hd__mux2_1
X_16733_ _16737_/B _16737_/C _16723_/X vssd1 vssd1 vccd1 vccd1 _16733_/Y sky130_fd_sc_hd__a21oi_1
X_19521_ _19542_/CLK _19521_/D vssd1 vssd1 vccd1 vccd1 _19521_/Q sky130_fd_sc_hd__dfxtp_2
X_13945_ _13945_/A vssd1 vssd1 vccd1 vccd1 _18609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19452_ _19671_/CLK _19452_/D vssd1 vssd1 vccd1 vccd1 _19452_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_184_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16664_ _16664_/A vssd1 vssd1 vccd1 vccd1 _16670_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13876_ _13777_/X _18579_/Q _13878_/S vssd1 vssd1 vccd1 vccd1 _13877_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15615_ _15615_/A vssd1 vssd1 vccd1 vccd1 _19300_/D sky130_fd_sc_hd__clkbuf_1
X_18403_ _18435_/A _18403_/B vssd1 vssd1 vccd1 vccd1 _20037_/D sky130_fd_sc_hd__nor2_1
XFILLER_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19383_ _19511_/CLK _19383_/D vssd1 vssd1 vccd1 vccd1 _19383_/Q sky130_fd_sc_hd__dfxtp_1
X_12827_ _12884_/A vssd1 vssd1 vccd1 vccd1 _16635_/A sky130_fd_sc_hd__clkbuf_2
X_16595_ _16820_/A vssd1 vssd1 vccd1 vccd1 _16783_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15431__S _15439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17212__A _17229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18334_ _12688_/B _18323_/X _18333_/X _18329_/X vssd1 vssd1 vccd1 vccd1 _20013_/D
+ sky130_fd_sc_hd__o211a_1
X_15546_ _19270_/Q _15238_/X _15550_/S vssd1 vssd1 vccd1 vccd1 _15547_/A sky130_fd_sc_hd__mux2_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12758_/A vssd1 vssd1 vccd1 vccd1 _13562_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16348__B1 _16347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12621__A2 _12620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11709_ _11856_/S _12632_/B _11708_/Y vssd1 vssd1 vccd1 vccd1 _11898_/D sky130_fd_sc_hd__o21a_1
X_18265_ _18265_/A vssd1 vssd1 vccd1 vccd1 _19986_/D sky130_fd_sc_hd__clkbuf_1
X_15477_ _15477_/A vssd1 vssd1 vccd1 vccd1 _19239_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12356__A _12356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12689_ _20015_/Q _12689_/B _12689_/C _09389_/A vssd1 vssd1 vccd1 vccd1 _12837_/B
+ sky130_fd_sc_hd__or4b_4
XANTENNA__11260__A _11260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17216_ _15784_/X _17212_/X _17214_/X _17215_/X vssd1 vssd1 vccd1 vccd1 _19838_/D
+ sky130_fd_sc_hd__o211a_1
X_14428_ _18812_/Q _14427_/X _14434_/S vssd1 vssd1 vccd1 vccd1 _14429_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18196_ _19956_/Q _19988_/Q _18196_/S vssd1 vssd1 vccd1 vccd1 _18197_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17866__B _17866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11188__A2 _11176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17147_ _17149_/A _17346_/B _17149_/C vssd1 vssd1 vccd1 vccd1 _17230_/A sky130_fd_sc_hd__nor3_2
X_14359_ _18790_/Q _13727_/X _14363_/S vssd1 vssd1 vccd1 vccd1 _14360_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10491__S0 _10390_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17078_ _17079_/A _17079_/C _17077_/Y vssd1 vssd1 vccd1 vccd1 _19787_/D sky130_fd_sc_hd__o21a_1
XFILLER_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16029_ _16029_/A vssd1 vssd1 vccd1 vccd1 _19436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10604__A _10604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__C1 _10994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__B2 _19905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19719_ _19720_/CLK _19719_/D vssd1 vssd1 vccd1 vccd1 _19719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16587__B1 _16577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09403_ _09358_/X _09401_/Y _09404_/B vssd1 vssd1 vccd1 vccd1 _09403_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16437__S _16437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15341__S _15345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13650__A _15228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17122__A _17122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _20020_/Q vssd1 vssd1 vccd1 vccd1 _16808_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16339__B1 _12444_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09265_ _11532_/A _11730_/B _11730_/C vssd1 vssd1 vccd1 vccd1 _09265_/X sky130_fd_sc_hd__or3_2
XANTENNA__11820__B1 _11816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17551__A2 _17533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11170__A _11170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09196_ _09196_/A vssd1 vssd1 vccd1 vccd1 _09269_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_140_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16172__S _16178_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09575__A _09975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17792__A _17792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__B _14074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10040_ _10040_/A vssd1 vssd1 vccd1 vccd1 _10700_/S sky130_fd_sc_hd__buf_4
XANTENNA__10234__S0 _10175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14842__A2_N _16315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13825__A _14650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11991_ _12194_/A _12104_/A vssd1 vssd1 vccd1 vccd1 _11992_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11990__D _17792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _15289_/A vssd1 vssd1 vccd1 vccd1 _14666_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10942_ _09955_/A _10940_/X _10941_/X vssd1 vssd1 vccd1 vccd1 _10942_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16578__B1 _16577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ _18518_/Q _13660_/X _13673_/S vssd1 vssd1 vccd1 vccd1 _13662_/A sky130_fd_sc_hd__mux2_1
X_10873_ _09513_/A _10872_/X _10955_/A vssd1 vssd1 vccd1 vccd1 _10873_/X sky130_fd_sc_hd__a21o_1
X_15400_ _14612_/X _19205_/Q _15406_/S vssd1 vssd1 vccd1 vccd1 _15401_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13560__A _13560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _19988_/Q _12593_/Y _12612_/S vssd1 vssd1 vccd1 vccd1 _12614_/B sky130_fd_sc_hd__mux2_2
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _13069_/X _19549_/Q _16382_/S vssd1 vssd1 vccd1 vccd1 _16381_/A sky130_fd_sc_hd__mux2_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _13592_/A _13592_/B vssd1 vssd1 vccd1 vccd1 _13592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15331_ _15331_/A vssd1 vssd1 vccd1 vccd1 _19174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12543_ _12538_/Y _12541_/X _12542_/Y vssd1 vssd1 vccd1 vccd1 _12543_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18050_ _18083_/A _18050_/B vssd1 vssd1 vccd1 vccd1 _18050_/X sky130_fd_sc_hd__or2_1
X_15262_ _15262_/A vssd1 vssd1 vccd1 vccd1 _19149_/D sky130_fd_sc_hd__clkbuf_1
X_12474_ _12474_/A vssd1 vssd1 vccd1 vccd1 _12474_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17001_ _17052_/A vssd1 vssd1 vccd1 vccd1 _17046_/A sky130_fd_sc_hd__buf_2
X_14213_ _14213_/A vssd1 vssd1 vccd1 vccd1 _18725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ _11537_/A _12667_/B vssd1 vssd1 vccd1 vccd1 _11425_/Y sky130_fd_sc_hd__nor2_1
X_15193_ _19128_/Q vssd1 vssd1 vccd1 vccd1 _15194_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_165_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ _18697_/Q _13739_/X _14146_/S vssd1 vssd1 vccd1 vccd1 _14145_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ _11579_/A _11356_/B vssd1 vssd1 vccd1 vccd1 _11580_/C sky130_fd_sc_hd__nand2_1
XFILLER_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ _10307_/A vssd1 vssd1 vccd1 vccd1 _10307_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18952_ _19053_/CLK _18952_/D vssd1 vssd1 vccd1 vccd1 _18952_/Q sky130_fd_sc_hd__dfxtp_1
X_14075_ _16062_/A _16371_/B vssd1 vssd1 vccd1 vccd1 _16809_/C sky130_fd_sc_hd__or2_4
XFILLER_112_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11287_ _11096_/A _11286_/X _18830_/Q vssd1 vssd1 vccd1 vccd1 _11287_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10225__S0 _09653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13026_ _19739_/Q _12912_/X _13025_/X _12917_/X vssd1 vssd1 vccd1 vccd1 _13026_/X
+ sky130_fd_sc_hd__a211o_2
X_17903_ _17899_/B _17903_/B vssd1 vssd1 vccd1 vccd1 _17904_/D sky130_fd_sc_hd__and2b_1
XFILLER_140_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10238_ _09750_/X _10227_/X _10236_/X _09757_/X _10237_/Y vssd1 vssd1 vccd1 vccd1
+ _12660_/B sky130_fd_sc_hd__o32a_4
X_18883_ _19311_/CLK _18883_/D vssd1 vssd1 vccd1 vccd1 _18883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15426__S _15428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10169_ _09479_/X _10164_/X _10166_/X _10168_/X _10205_/A vssd1 vssd1 vccd1 vccd1
+ _10169_/X sky130_fd_sc_hd__a221o_1
X_17834_ _17785_/X _17831_/X _17833_/Y _17794_/X vssd1 vssd1 vccd1 vccd1 _17834_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14977_ _19028_/Q _14456_/X _14983_/S vssd1 vssd1 vccd1 vccd1 _14978_/A sky130_fd_sc_hd__mux2_1
X_17765_ _17827_/A vssd1 vssd1 vccd1 vccd1 _17765_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19504_ _19504_/CLK _19504_/D vssd1 vssd1 vccd1 vccd1 _19504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13928_ _18295_/A _15373_/B _14151_/B vssd1 vssd1 vccd1 vccd1 _13985_/A sky130_fd_sc_hd__nor3_4
X_16716_ _16717_/B _16717_/C _19677_/Q vssd1 vssd1 vccd1 vccd1 _16718_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13173__C _19888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17696_ _17600_/X _17695_/Y _17530_/A vssd1 vssd1 vccd1 vccd1 _17696_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_90_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19435_ _19500_/CLK _19435_/D vssd1 vssd1 vccd1 vccd1 _19435_/Q sky130_fd_sc_hd__dfxtp_1
X_16647_ _16672_/A _16647_/B _16647_/C vssd1 vssd1 vccd1 vccd1 _19656_/D sky130_fd_sc_hd__nor3_1
X_13859_ _13746_/X _18571_/Q _13867_/S vssd1 vssd1 vccd1 vccd1 _13860_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19366_ _19366_/CLK _19366_/D vssd1 vssd1 vccd1 vccd1 _19366_/Q sky130_fd_sc_hd__dfxtp_1
X_16578_ _19633_/Q _16582_/C _16577_/X vssd1 vssd1 vccd1 vccd1 _16578_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__15792__A1 _19915_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11802__A0 _20044_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18317_ _18341_/A vssd1 vssd1 vccd1 vccd1 _18317_/X sky130_fd_sc_hd__clkbuf_2
X_15529_ _15529_/A vssd1 vssd1 vccd1 vccd1 _19262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19297_ _19553_/CLK _19297_/D vssd1 vssd1 vccd1 vccd1 _19297_/Q sky130_fd_sc_hd__dfxtp_1
X_18248_ _18248_/A vssd1 vssd1 vccd1 vccd1 _19978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15397__A _15443_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18179_ _16332_/A _19980_/Q _18181_/S vssd1 vssd1 vccd1 vccd1 _18180_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14505__S _14513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12814__A _12853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09952_ _10825_/A _09952_/B vssd1 vssd1 vccd1 vccd1 _09952_/X sky130_fd_sc_hd__and2_1
XFILLER_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12015__A2_N _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _10229_/A _09883_/B vssd1 vssd1 vccd1 vccd1 _09883_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10767__S1 _10030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14240__S _14246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09909__S0 _10244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10844__B2 _19902_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16167__S _16167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14476__A _14476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09317_ _18331_/A _19999_/Q _19887_/Q _09315_/X _09316_/X vssd1 vssd1 vccd1 vccd1
+ _09320_/C sky130_fd_sc_hd__o2111ai_1
XFILLER_139_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17787__A _18009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _09275_/C _09248_/B _11730_/B vssd1 vssd1 vccd1 vccd1 _17378_/B sky130_fd_sc_hd__or3_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_132_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ _20025_/Q vssd1 vssd1 vccd1 vccd1 _09191_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_5_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11210_ _09610_/A _11199_/X _11209_/X _09618_/A _19895_/Q vssd1 vssd1 vccd1 vccd1
+ _11348_/A sky130_fd_sc_hd__a32o_4
XFILLER_108_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12190_ _12190_/A vssd1 vssd1 vccd1 vccd1 _12190_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15838__A2 _13533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ _11141_/A _11141_/B vssd1 vssd1 vccd1 vccd1 _11141_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18411__A _18412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11072_ _19361_/Q _18975_/Q _19425_/Q _18544_/Q _11000_/S _10083_/A vssd1 vssd1 vccd1
+ vccd1 _11073_/B sky130_fd_sc_hd__mux4_1
Xoutput77 _12204_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[15] sky130_fd_sc_hd__buf_2
Xoutput88 _12463_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[25] sky130_fd_sc_hd__buf_2
XFILLER_110_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput99 _11940_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[6] sky130_fd_sc_hd__buf_2
XFILLER_103_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14900_ _14653_/X _18994_/Q _14900_/S vssd1 vssd1 vccd1 vccd1 _14901_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10758__S1 _10030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _11283_/A vssd1 vssd1 vccd1 vccd1 _10024_/A sky130_fd_sc_hd__buf_2
XFILLER_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_1_clock clkbuf_1_0_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_15880_ _15880_/A vssd1 vssd1 vccd1 vccd1 _19370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input23_A io_dbus_rdata[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17460__A1 _12385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ _14831_/A vssd1 vssd1 vccd1 vccd1 _14831_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17550_ _17940_/A vssd1 vssd1 vccd1 vccd1 _17646_/A sky130_fd_sc_hd__clkbuf_2
X_14762_ _18936_/Q _14382_/X _14764_/S vssd1 vssd1 vccd1 vccd1 _14763_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11974_ _11974_/A _19585_/Q _12240_/B vssd1 vssd1 vccd1 vccd1 _12027_/C sky130_fd_sc_hd__and3_1
XFILLER_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16501_ _19661_/Q _19663_/Q _19662_/Q _16656_/A vssd1 vssd1 vccd1 vccd1 _16664_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_56_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_57_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13713_ _15276_/A vssd1 vssd1 vccd1 vccd1 _14653_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17481_ _17479_/X _17480_/X _17486_/S vssd1 vssd1 vccd1 vccd1 _17481_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10925_ _10929_/A _10925_/B vssd1 vssd1 vccd1 vccd1 _10925_/Y sky130_fd_sc_hd__nor2_1
X_14693_ _14750_/S vssd1 vssd1 vccd1 vccd1 _14702_/S sky130_fd_sc_hd__buf_2
XFILLER_60_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19220_ _19401_/CLK _19220_/D vssd1 vssd1 vccd1 vccd1 _19220_/Q sky130_fd_sc_hd__dfxtp_1
X_16432_ _16432_/A vssd1 vssd1 vccd1 vccd1 _19572_/D sky130_fd_sc_hd__clkbuf_1
X_13644_ _18514_/Q _13643_/X _13652_/S vssd1 vssd1 vccd1 vccd1 _13645_/A sky130_fd_sc_hd__mux2_1
X_10856_ _10000_/X _10846_/Y _10851_/X _10855_/Y _09738_/A vssd1 vssd1 vccd1 vccd1
+ _10856_/X sky130_fd_sc_hd__o311a_1
XFILLER_16_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19151_ _19412_/CLK _19151_/D vssd1 vssd1 vccd1 vccd1 _19151_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16363_ _16367_/B _16363_/B vssd1 vssd1 vccd1 vccd1 _16363_/Y sky130_fd_sc_hd__nand2_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13575_/A vssd1 vssd1 vccd1 vccd1 _18502_/D sky130_fd_sc_hd__clkbuf_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10790_/A _10787_/B vssd1 vssd1 vccd1 vccd1 _10787_/Y sky130_fd_sc_hd__nor2_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18102_ _18098_/B _18097_/B _17794_/X _18101_/Y vssd1 vssd1 vccd1 vccd1 _18102_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15314_ _15371_/S vssd1 vssd1 vccd1 vccd1 _15323_/S sky130_fd_sc_hd__buf_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19082_ _19306_/CLK _19082_/D vssd1 vssd1 vccd1 vccd1 _19082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12526_ _17538_/A _18079_/A _12499_/B vssd1 vssd1 vccd1 vccd1 _12527_/B sky130_fd_sc_hd__a21o_1
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10694__S0 _10690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16294_ _16294_/A vssd1 vssd1 vccd1 vccd1 _19530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18033_ _18033_/A _18033_/B vssd1 vssd1 vccd1 vccd1 _18033_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15245_ _19144_/Q _15244_/X _15245_/S vssd1 vssd1 vccd1 vccd1 _15246_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12457_ _12457_/A _18058_/B vssd1 vssd1 vccd1 vccd1 _12458_/B sky130_fd_sc_hd__or2_1
XFILLER_173_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12634__A _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output91_A _12538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _11408_/A vssd1 vssd1 vccd1 vccd1 _11408_/Y sky130_fd_sc_hd__inv_2
X_15176_ _15176_/A vssd1 vssd1 vccd1 vccd1 _19119_/D sky130_fd_sc_hd__clkbuf_1
X_12388_ _12388_/A _12388_/B vssd1 vssd1 vccd1 vccd1 _12391_/A sky130_fd_sc_hd__nor2_2
XFILLER_67_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12760__A1 _19813_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14127_ _18689_/Q _13706_/X _14131_/S vssd1 vssd1 vccd1 vccd1 _14128_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11339_ _19484_/Q _18896_/Q _18933_/Q _18507_/Q _11030_/A _09658_/A vssd1 vssd1 vccd1
+ vccd1 _11339_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19984_ _19986_/CLK _19984_/D vssd1 vssd1 vccd1 vccd1 _19984_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18321__A _18321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14058_ _14058_/A vssd1 vssd1 vccd1 vccd1 _18659_/D sky130_fd_sc_hd__clkbuf_1
X_18935_ _19486_/CLK _18935_/D vssd1 vssd1 vccd1 vccd1 _18935_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13304__A3 _09349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13009_ _15197_/A vssd1 vssd1 vccd1 vccd1 _13009_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14060__S _14068_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18866_ _19196_/CLK _18866_/D vssd1 vssd1 vccd1 vccd1 _18866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17817_ _17820_/A _17820_/B vssd1 vssd1 vccd1 vccd1 _17817_/X sky130_fd_sc_hd__and2_1
XANTENNA__10601__B _12651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18797_ _19484_/CLK _18797_/D vssd1 vssd1 vccd1 vccd1 _18797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17748_ _17746_/Y _17747_/X _17748_/S vssd1 vssd1 vccd1 vccd1 _17748_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17679_ _17602_/S _17677_/X _17678_/X vssd1 vssd1 vccd1 vccd1 _17679_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19418_ _19418_/CLK _19418_/D vssd1 vssd1 vccd1 vccd1 _19418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19349_ _19844_/CLK _19349_/D vssd1 vssd1 vccd1 vccd1 _19349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16714__B1 _16667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13528__B1 _12810_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14235__S _14235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_132_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19487_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09853__A _09926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09935_ _19380_/Q _18994_/Q _19444_/Q _18563_/Q _10218_/S _09929_/X vssd1 vssd1 vccd1
+ vccd1 _09936_/B sky130_fd_sc_hd__mux4_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10999__A _10999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15066__S _15072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09866_ _10270_/S vssd1 vssd1 vccd1 vccd1 _10218_/S sky130_fd_sc_hd__clkbuf_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_147_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19666_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _19512_/Q _18924_/Q _18961_/Q _18535_/Q _09724_/S _09688_/A vssd1 vssd1 vccd1
+ vccd1 _09797_/X sky130_fd_sc_hd__mux4_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15590__A _15646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_9_0_clock clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_54_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _18775_/Q _19046_/Q _19270_/Q _19014_/Q _10753_/S _10014_/A vssd1 vssd1 vccd1
+ vccd1 _10710_/X sky130_fd_sc_hd__mux4_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _17381_/A _11690_/B _11694_/A _11690_/D vssd1 vssd1 vccd1 vccd1 _11690_/X
+ sky130_fd_sc_hd__and4_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12438__B _19602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10641_ _11452_/A _10641_/B vssd1 vssd1 vccd1 vccd1 _10641_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14827__A1_N _18311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10676__S0 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ _19945_/Q vssd1 vssd1 vccd1 vccd1 _16313_/A sky130_fd_sc_hd__clkbuf_2
X_10572_ _18650_/Q _19241_/Q _19403_/Q _18618_/Q _10382_/A _09815_/A vssd1 vssd1 vccd1
+ vccd1 _10572_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15749__B _18452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12311_ _12339_/C _12365_/D vssd1 vssd1 vccd1 vccd1 _12311_/X sky130_fd_sc_hd__xor2_1
XFILLER_155_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16181__A1 _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ _13282_/Y _13283_/X _13290_/X _13337_/A _13351_/A vssd1 vssd1 vccd1 vccd1
+ _13292_/B sky130_fd_sc_hd__a221o_1
XFILLER_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15030_ _15030_/A vssd1 vssd1 vccd1 vccd1 _19051_/D sky130_fd_sc_hd__clkbuf_1
X_12242_ _19530_/Q _11782_/X _12026_/X vssd1 vssd1 vccd1 vccd1 _12242_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10979__S1 _11330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ _12111_/A _12111_/B _12147_/A _12172_/Y vssd1 vssd1 vccd1 vccd1 _12174_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_123_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11124_ _19360_/Q _18974_/Q _19424_/Q _18543_/Q _11004_/S _11065_/X vssd1 vssd1 vccd1
+ vccd1 _11125_/B sky130_fd_sc_hd__mux4_1
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16981_ _19752_/Q _16981_/B vssd1 vssd1 vccd1 vccd1 _16983_/B sky130_fd_sc_hd__nor2_1
XFILLER_150_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12901__B _12901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18720_ _19570_/CLK _18720_/D vssd1 vssd1 vccd1 vccd1 _18720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11055_ _11125_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11055_/X sky130_fd_sc_hd__or2_1
X_15932_ _19393_/Q _15215_/X _15940_/S vssd1 vssd1 vccd1 vccd1 _15933_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10006_ _10006_/A vssd1 vssd1 vccd1 vccd1 _10007_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18651_ _19501_/CLK _18651_/D vssd1 vssd1 vccd1 vccd1 _18651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15863_ _15863_/A vssd1 vssd1 vccd1 vccd1 _19362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14814_ _14814_/A vssd1 vssd1 vccd1 vccd1 _18959_/D sky130_fd_sc_hd__clkbuf_1
X_17602_ _17527_/B _17601_/X _17602_/S vssd1 vssd1 vccd1 vccd1 _17602_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18582_ _19431_/CLK _18582_/D vssd1 vssd1 vccd1 vccd1 _18582_/Q sky130_fd_sc_hd__dfxtp_1
X_15794_ _15794_/A vssd1 vssd1 vccd1 vccd1 _19346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14745_ _14745_/A vssd1 vssd1 vccd1 vccd1 _18924_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17533_ _17533_/A vssd1 vssd1 vccd1 vccd1 _17533_/X sky130_fd_sc_hd__buf_2
X_11957_ _11957_/A _11957_/B vssd1 vssd1 vccd1 vccd1 _11957_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17464_ _19968_/Q _12076_/A _17464_/S vssd1 vssd1 vccd1 vccd1 _17866_/B sky130_fd_sc_hd__mux2_4
X_10908_ _10908_/A vssd1 vssd1 vccd1 vccd1 _10908_/Y sky130_fd_sc_hd__inv_2
X_14676_ _14675_/X _18895_/Q _14676_/S vssd1 vssd1 vccd1 vccd1 _14677_/A sky130_fd_sc_hd__mux2_1
X_11888_ _16208_/S vssd1 vssd1 vccd1 vccd1 _12032_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16415_ _13357_/X _19565_/Q _16415_/S vssd1 vssd1 vccd1 vccd1 _16416_/A sky130_fd_sc_hd__mux2_1
X_19203_ _19203_/CLK _19203_/D vssd1 vssd1 vccd1 vccd1 _19203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13627_ _18510_/Q _13626_/X _13631_/S vssd1 vssd1 vccd1 vccd1 _13628_/A sky130_fd_sc_hd__mux2_1
X_10839_ _19461_/Q _19299_/Q _18708_/Q _18478_/Q _09984_/X _09970_/X vssd1 vssd1 vccd1
+ vccd1 _10840_/B sky130_fd_sc_hd__mux4_1
XFILLER_20_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17395_ _17395_/A _17395_/B vssd1 vssd1 vccd1 vccd1 _17396_/D sky130_fd_sc_hd__nor2_1
XANTENNA__14844__A _18299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18316__A _18316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17220__A _17220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19134_ _19292_/CLK _19134_/D vssd1 vssd1 vccd1 vccd1 _19134_/Q sky130_fd_sc_hd__dfxtp_1
X_16346_ _16346_/A vssd1 vssd1 vccd1 vccd1 _19540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13558_ _18500_/Q _13557_/X _13558_/S vssd1 vssd1 vccd1 vccd1 _13559_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12981__A1 _18465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12509_ _12509_/A vssd1 vssd1 vccd1 vccd1 _12509_/Y sky130_fd_sc_hd__inv_8
X_19065_ _19129_/CLK _19065_/D vssd1 vssd1 vccd1 vccd1 _19065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16172__A1 _14628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16277_ _16277_/A vssd1 vssd1 vccd1 vccd1 _19527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13489_ _13489_/A vssd1 vssd1 vccd1 vccd1 _18496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18016_ _17928_/X _17848_/Y _18015_/X _17953_/X vssd1 vssd1 vccd1 vccd1 _18016_/X
+ sky130_fd_sc_hd__o211a_1
X_15228_ _15228_/A vssd1 vssd1 vccd1 vccd1 _15228_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13894__S _13900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15159_ _19111_/Q vssd1 vssd1 vccd1 vccd1 _15160_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__11092__S0 _11035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16475__A2 _12494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19967_ _19971_/CLK _19967_/D vssd1 vssd1 vccd1 vccd1 _19967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19511_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09720_ _09673_/Y _09697_/Y _09699_/Y _09713_/Y _09719_/X vssd1 vssd1 vccd1 vccd1
+ _09720_/X sky130_fd_sc_hd__o221a_1
XANTENNA__13195__A _15228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18918_ _19508_/CLK _18918_/D vssd1 vssd1 vccd1 vccd1 _18918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19898_ _19966_/CLK _19898_/D vssd1 vssd1 vccd1 vccd1 _19898_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_110_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09651_ _09651_/A vssd1 vssd1 vccd1 vccd1 _10270_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_110_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18849_ _19308_/CLK _18849_/D vssd1 vssd1 vccd1 vccd1 _18849_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15614__S _15622_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09582_ _18969_/Q vssd1 vssd1 vccd1 vccd1 _11199_/A sky130_fd_sc_hd__buf_4
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_79_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19573_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12539__A _19606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17727__A2 _17729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14754__A _14810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12972__A1 _18459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16163__A1 _14615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19987_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09583__A _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10830__S0 _10811_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12721__B _12837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09918_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09918_/X sky130_fd_sc_hd__or2_1
XANTENNA__11618__A _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12488__A0 _12485_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20038_ _20052_/CLK _20038_/D vssd1 vssd1 vccd1 vccd1 _20038_/Q sky130_fd_sc_hd__dfxtp_1
X_09849_ _10591_/S vssd1 vssd1 vccd1 vccd1 _10337_/A sky130_fd_sc_hd__buf_2
XANTENNA__18422__A1_N _18340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12860_ _16528_/A _19772_/Q _17129_/S _12859_/X vssd1 vssd1 vccd1 vccd1 _19772_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11138__S1 _10917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11812_/A _17431_/A vssd1 vssd1 vccd1 vccd1 _11813_/A sky130_fd_sc_hd__and2_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12791_ _16875_/A _12791_/B _19807_/Q vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__or3b_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12449__A _18336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14530_/A vssd1 vssd1 vccd1 vccd1 _18843_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11742_ _11910_/A vssd1 vssd1 vccd1 vccd1 _11976_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17959__B _17960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14461_/A vssd1 vssd1 vccd1 vccd1 _18822_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__A2_N _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11673_ _11673_/A _17379_/C _11673_/C _11672_/X vssd1 vssd1 vccd1 vccd1 _11901_/B
+ sky130_fd_sc_hd__or4b_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16200_ _19513_/Q _14669_/A _16200_/S vssd1 vssd1 vccd1 vccd1 _16201_/A sky130_fd_sc_hd__mux2_1
X_13412_ _15270_/A vssd1 vssd1 vccd1 vccd1 _13412_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10624_ _11443_/A vssd1 vssd1 vccd1 vccd1 _11438_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09758__A _19924_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17180_ _17180_/A _17180_/B vssd1 vssd1 vccd1 vccd1 _17180_/X sky130_fd_sc_hd__or2_1
X_14392_ _14596_/A vssd1 vssd1 vccd1 vccd1 _14392_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _16131_/A vssd1 vssd1 vccd1 vccd1 _19482_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11310__S1 _11260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12963__A1 _18452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13343_ _13343_/A vssd1 vssd1 vccd1 vccd1 _13343_/X sky130_fd_sc_hd__clkbuf_2
X_10555_ _10555_/A _12653_/B vssd1 vssd1 vccd1 vccd1 _10556_/B sky130_fd_sc_hd__nor2_1
XANTENNA__16154__A1 _14602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16062_ _16062_/A _16062_/B vssd1 vssd1 vccd1 vccd1 _16119_/A sky130_fd_sc_hd__or2_4
X_13274_ _13297_/C _13274_/B vssd1 vssd1 vccd1 vccd1 _13274_/Y sky130_fd_sc_hd__nor2_1
X_10486_ _10486_/A _10486_/B vssd1 vssd1 vccd1 vccd1 _10486_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15013_ _15059_/S vssd1 vssd1 vccd1 vccd1 _15022_/S sky130_fd_sc_hd__buf_2
XFILLER_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12225_ _12252_/A _12225_/B vssd1 vssd1 vccd1 vccd1 _12226_/B sky130_fd_sc_hd__nor2_2
XANTENNA__11074__S0 _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19821_ _19852_/CLK _19821_/D vssd1 vssd1 vccd1 vccd1 _19821_/Q sky130_fd_sc_hd__dfxtp_1
X_12156_ _17187_/A _12157_/C _19830_/Q vssd1 vssd1 vccd1 vccd1 _12156_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12631__B _12631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11107_ _19898_/Q vssd1 vssd1 vccd1 vccd1 _11107_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19752_ _19756_/CLK _19752_/D vssd1 vssd1 vccd1 vccd1 _19752_/Q sky130_fd_sc_hd__dfxtp_1
X_16964_ _16964_/A _16964_/B vssd1 vssd1 vccd1 vccd1 _16965_/D sky130_fd_sc_hd__and2_1
X_12087_ _12086_/A _12086_/C _19589_/Q vssd1 vssd1 vccd1 vccd1 _12088_/D sky130_fd_sc_hd__a21o_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11377__S1 _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18703_ _19666_/CLK _18703_/D vssd1 vssd1 vccd1 vccd1 _18703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15915_ _15915_/A vssd1 vssd1 vccd1 vccd1 _19386_/D sky130_fd_sc_hd__clkbuf_1
X_11038_ _11141_/A _11037_/X _09703_/A vssd1 vssd1 vccd1 vccd1 _11038_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19683_ _19720_/CLK _19683_/D vssd1 vssd1 vccd1 vccd1 _19683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16895_ _16923_/B _16900_/D _19730_/Q vssd1 vssd1 vccd1 vccd1 _16897_/B sky130_fd_sc_hd__a21oi_1
XFILLER_76_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17215__A _18289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18634_ _19952_/CLK _18634_/D vssd1 vssd1 vccd1 vccd1 _18634_/Q sky130_fd_sc_hd__dfxtp_1
X_15846_ _16134_/A _15990_/B vssd1 vssd1 vccd1 vccd1 _15903_/A sky130_fd_sc_hd__or2_4
XFILLER_94_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18565_ _19092_/CLK _18565_/D vssd1 vssd1 vccd1 vccd1 _18565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _12989_/A vssd1 vssd1 vccd1 vccd1 _12989_/X sky130_fd_sc_hd__clkbuf_2
X_15777_ _16364_/S _17209_/A vssd1 vssd1 vccd1 vccd1 _16315_/B sky130_fd_sc_hd__nor2_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17516_ _17473_/X _17513_/Y _17729_/A vssd1 vssd1 vccd1 vccd1 _17516_/X sky130_fd_sc_hd__mux2_1
X_14728_ _14728_/A vssd1 vssd1 vccd1 vccd1 _18916_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10888__S0 _09983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18496_ _19317_/CLK _18496_/D vssd1 vssd1 vccd1 vccd1 _18496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13889__S _13889_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14659_ _14659_/A vssd1 vssd1 vccd1 vccd1 _18889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17447_ _17447_/A vssd1 vssd1 vccd1 vccd1 _17937_/A sky130_fd_sc_hd__buf_2
XANTENNA__16393__A1 _19555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09668__A _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17378_ _17378_/A _17378_/B vssd1 vssd1 vccd1 vccd1 _17379_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11757__A2 _12633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19117_ _19565_/CLK _19117_/D vssd1 vssd1 vccd1 vccd1 _19117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16145__A1 _14589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16329_ _16369_/S vssd1 vssd1 vccd1 vccd1 _16365_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19048_ _19495_/CLK _19048_/D vssd1 vssd1 vccd1 vccd1 _19048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_179_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14513__S _14513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10717__B1 _10056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13129__S _13196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09703_ _09703_/A vssd1 vssd1 vccd1 vccd1 _09999_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09634_ _10544_/A vssd1 vssd1 vccd1 vccd1 _10500_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09565_ _10161_/A _09551_/X _09567_/A vssd1 vssd1 vccd1 vccd1 _09565_/X sky130_fd_sc_hd__a21o_1
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11445__A1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ _11191_/S vssd1 vssd1 vccd1 vccd1 _10937_/S sky130_fd_sc_hd__buf_4
XFILLER_168_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14484__A _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09578__A _10307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11620__B _11910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10517__A _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10340_ _10588_/A vssd1 vssd1 vccd1 vccd1 _10486_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10271_ _10271_/A _10271_/B vssd1 vssd1 vccd1 vccd1 _10271_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12732__A _18453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12010_ _19825_/Q vssd1 vssd1 vccd1 vccd1 _17176_/A sky130_fd_sc_hd__buf_2
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11381__B1 hold15/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11348__A _11348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13961_ _18617_/Q _13672_/X _13961_/S vssd1 vssd1 vccd1 vccd1 _13962_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12912_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12912_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15700_ _15700_/A vssd1 vssd1 vccd1 vccd1 _15700_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16680_ _16680_/A _19668_/Q _16680_/C vssd1 vssd1 vccd1 vccd1 _16682_/B sky130_fd_sc_hd__and3_1
XFILLER_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09760__B _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ _13799_/X _18586_/Q _13900_/S vssd1 vssd1 vccd1 vccd1 _13893_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15631_ _14634_/X _19308_/Q _15633_/S vssd1 vssd1 vccd1 vccd1 _15632_/A sky130_fd_sc_hd__mux2_1
X_12843_ _19772_/Q _12893_/B vssd1 vssd1 vccd1 vccd1 _12843_/X sky130_fd_sc_hd__and2_1
XFILLER_62_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18376__A1_N _18288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_opt_4_0_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11436__A1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15562_ _15562_/A vssd1 vssd1 vccd1 vccd1 _19277_/D sky130_fd_sc_hd__clkbuf_1
X_18350_ _16808_/A _18302_/B _18349_/X _18341_/X vssd1 vssd1 vccd1 vccd1 _20020_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _15700_/A vssd1 vssd1 vccd1 vccd1 _13587_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18364__A2 _14476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
X_17301_ _17301_/A vssd1 vssd1 vccd1 vccd1 _19873_/D sky130_fd_sc_hd__clkbuf_1
X_14513_ _13764_/X _18836_/Q _14513_/S vssd1 vssd1 vccd1 vccd1 _14514_/A sky130_fd_sc_hd__mux2_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11725_ _11729_/A _17378_/A _12598_/D vssd1 vssd1 vccd1 vccd1 _11733_/A sky130_fd_sc_hd__o21ai_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _15493_/A vssd1 vssd1 vccd1 vccd1 _19246_/D sky130_fd_sc_hd__clkbuf_1
X_18281_ _19993_/Q _18281_/B vssd1 vssd1 vccd1 vccd1 _18281_/X sky130_fd_sc_hd__or2_1
XFILLER_159_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13189__A1 _15716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14444_ _18817_/Q _14443_/X _14450_/S vssd1 vssd1 vccd1 vccd1 _14445_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17232_ _18289_/A vssd1 vssd1 vccd1 vccd1 _17232_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11656_ _13324_/A vssd1 vssd1 vccd1 vccd1 _11656_/X sky130_fd_sc_hd__buf_2
XFILLER_156_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10607_ _10734_/A _10605_/X _10613_/A vssd1 vssd1 vccd1 vccd1 _10607_/X sky130_fd_sc_hd__a21o_1
X_17163_ _17160_/Y _17153_/X _17162_/Y _17142_/X vssd1 vssd1 vccd1 vccd1 _19821_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10098__S1 _09515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14375_ _14375_/A vssd1 vssd1 vccd1 vccd1 _18795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11587_ _11579_/B _11580_/Y _11582_/X _11586_/X vssd1 vssd1 vccd1 vccd1 _11587_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16114_ _16114_/A vssd1 vssd1 vccd1 vccd1 _19474_/D sky130_fd_sc_hd__clkbuf_1
X_13326_ _16301_/B _13335_/C vssd1 vssd1 vccd1 vccd1 _13326_/X sky130_fd_sc_hd__xor2_1
X_10538_ _18587_/Q _18848_/Q _18747_/Q _19082_/Q _10266_/A _10592_/A vssd1 vssd1 vccd1
+ vccd1 _10538_/X sky130_fd_sc_hd__mux4_1
X_17094_ _17095_/A _17095_/C _17093_/Y vssd1 vssd1 vccd1 vccd1 _19793_/D sky130_fd_sc_hd__o21a_1
XFILLER_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_180_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16045_ _13433_/X _19444_/Q _16045_/S vssd1 vssd1 vccd1 vccd1 _16046_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13738__A _15295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13257_ input5/X _13172_/X _13175_/X vssd1 vssd1 vccd1 vccd1 _13257_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11047__S0 _10018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ _18780_/Q _19051_/Q _19275_/Q _19019_/Q _10382_/X _10462_/X vssd1 vssd1 vccd1
+ vccd1 _10469_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14333__S _14341_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12642__A _12651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12208_ _14477_/B vssd1 vssd1 vccd1 vccd1 _12208_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10175__A1 _19153_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13188_ _19651_/Q _12887_/A _12889_/A _19783_/Q _13187_/X vssd1 vssd1 vccd1 vccd1
+ _15716_/B sky130_fd_sc_hd__a221o_2
XFILLER_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19804_ _19804_/CLK _19804_/D vssd1 vssd1 vccd1 vccd1 _19804_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15953__A _15975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _12252_/A _12139_/B vssd1 vssd1 vccd1 vccd1 _12140_/B sky130_fd_sc_hd__nor2_1
XFILLER_111_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17996_ _18001_/A _18001_/B vssd1 vssd1 vccd1 vccd1 _18000_/B sky130_fd_sc_hd__and2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09317__B1 _19887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19735_ _19737_/CLK _19735_/D vssd1 vssd1 vccd1 vccd1 _19735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16947_ _16958_/A _16945_/B _16946_/Y vssd1 vssd1 vccd1 vccd1 _19743_/D sky130_fd_sc_hd__o21a_1
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19666_ _19666_/CLK _19666_/D vssd1 vssd1 vccd1 vccd1 _19666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09963__S1 _09515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16878_ _16898_/A vssd1 vssd1 vccd1 vccd1 _16897_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18617_ _19431_/CLK _18617_/D vssd1 vssd1 vccd1 vccd1 _18617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15829_ _19921_/Q _15828_/X _15840_/S vssd1 vssd1 vccd1 vccd1 _15829_/X sky130_fd_sc_hd__mux2_1
X_19597_ _19601_/CLK _19597_/D vssd1 vssd1 vccd1 vccd1 _19597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09350_ _09350_/A vssd1 vssd1 vccd1 vccd1 _13353_/A sky130_fd_sc_hd__buf_4
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12624__B1 _16303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18548_ _19555_/CLK _18548_/D vssd1 vssd1 vccd1 vccd1 _18548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10635__C1 _09603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11978__A2 _11972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09281_ _20040_/Q _20039_/Q _20038_/Q _20037_/Q vssd1 vssd1 vccd1 vccd1 _11640_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_61_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18479_ _19430_/CLK _18479_/D vssd1 vssd1 vccd1 vccd1 _18479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11721__A _12475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18107__A2 _17558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17315__A0 _15839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10337__A _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15339__S _15345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11168__A _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09617_ _09617_/A vssd1 vssd1 vccd1 vccd1 _09618_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09548_ _10734_/A vssd1 vssd1 vccd1 vccd1 _10294_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09479_ _09479_/A vssd1 vssd1 vccd1 vccd1 _09479_/X sky130_fd_sc_hd__buf_2
XANTENNA__13322__S _13358_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _11510_/A _11510_/B vssd1 vssd1 vccd1 vccd1 _11510_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12490_ _12208_/X _12488_/X _12489_/X vssd1 vssd1 vccd1 vccd1 _12490_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ _18664_/Q _19255_/Q _19417_/Q _18632_/Q _10625_/X _10604_/A vssd1 vssd1 vccd1
+ vccd1 _11441_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14160_ _14160_/A vssd1 vssd1 vccd1 vccd1 _18701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11372_ _18680_/Q _19175_/Q _11372_/S vssd1 vssd1 vccd1 vccd1 _11372_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09890__S0 _09872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13111_ _18474_/Q _13109_/X _13196_/S vssd1 vssd1 vccd1 vccd1 _13112_/A sky130_fd_sc_hd__mux2_1
X_10323_ _10323_/A vssd1 vssd1 vccd1 vccd1 _10323_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15249__S _15261_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14091_ _14091_/A vssd1 vssd1 vccd1 vccd1 _18672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12146__A2 _17884_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13042_ _18504_/Q _13077_/B vssd1 vssd1 vccd1 vccd1 _13042_/X sky130_fd_sc_hd__and2_1
XANTENNA_input53_A io_ibus_inst[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ _10254_/A _10254_/B vssd1 vssd1 vccd1 vccd1 _10254_/X sky130_fd_sc_hd__or2_1
XANTENNA__17972__B _17973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13992__S _13994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17850_ _11625_/B _17853_/B _17748_/S _17849_/X vssd1 vssd1 vccd1 vccd1 _17850_/X
+ sky130_fd_sc_hd__o211a_1
X_10185_ _19507_/Q _18919_/Q _18956_/Q _18530_/Q _09881_/X _10219_/A vssd1 vssd1 vccd1
+ vccd1 _10185_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16293__A0 _19530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09771__A _10205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16801_ _19705_/Q _16799_/B _16768_/X vssd1 vssd1 vccd1 vccd1 _16801_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17781_ _17827_/A vssd1 vssd1 vccd1 vccd1 _17781_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14993_ _14993_/A vssd1 vssd1 vccd1 vccd1 _19034_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14389__A _14472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13293__A _15247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19520_ _19837_/CLK _19520_/D vssd1 vssd1 vccd1 vccd1 _19520_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_75_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16732_ _19681_/Q _16728_/C _16731_/Y vssd1 vssd1 vccd1 vccd1 _19681_/D sky130_fd_sc_hd__o21a_1
XANTENNA__11201__S0 _11306_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__A1 _17379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13944_ _18609_/Q _13639_/X _13950_/S vssd1 vssd1 vccd1 vccd1 _13945_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_127_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10865__C1 _10063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19451_ _19577_/CLK _19451_/D vssd1 vssd1 vccd1 vccd1 _19451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16663_ _16672_/A _16663_/B _16663_/C vssd1 vssd1 vccd1 vccd1 _19662_/D sky130_fd_sc_hd__nor3_1
XFILLER_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13875_ _13875_/A vssd1 vssd1 vccd1 vccd1 _18578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18402_ _18435_/A _18402_/B vssd1 vssd1 vccd1 vccd1 _20036_/D sky130_fd_sc_hd__nor2_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15614_ _14608_/X _19300_/Q _15622_/S vssd1 vssd1 vccd1 vccd1 _15615_/A sky130_fd_sc_hd__mux2_1
X_12826_ _12795_/X _12796_/X _12822_/X _12825_/X vssd1 vssd1 vccd1 vccd1 _19806_/D
+ sky130_fd_sc_hd__a22o_1
X_19382_ _19510_/CLK _19382_/D vssd1 vssd1 vccd1 vccd1 _19382_/Q sky130_fd_sc_hd__dfxtp_1
X_16594_ _19638_/Q _16597_/C _16593_/Y vssd1 vssd1 vccd1 vccd1 _19638_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18333_ _18333_/A _18333_/B vssd1 vssd1 vccd1 vccd1 _18333_/X sky130_fd_sc_hd__or2_1
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15545_ _15545_/A vssd1 vssd1 vccd1 vccd1 _19269_/D sky130_fd_sc_hd__clkbuf_1
X_12757_ _13099_/A vssd1 vssd1 vccd1 vccd1 _12758_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16348__A1 _16347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12637__A _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15013__A _15059_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ _11704_/X _11706_/X _11707_/X _11894_/A vssd1 vssd1 vccd1 vccd1 _11708_/Y
+ sky130_fd_sc_hd__o211ai_2
X_15476_ _19239_/Q _15241_/X _15478_/S vssd1 vssd1 vccd1 vccd1 _15477_/A sky130_fd_sc_hd__mux2_1
X_18264_ _19986_/Q _12561_/A _18264_/S vssd1 vssd1 vccd1 vccd1 _18265_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12688_ _12688_/A _12688_/B vssd1 vssd1 vccd1 vccd1 _12689_/C sky130_fd_sc_hd__or2_1
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14427_ _14631_/A vssd1 vssd1 vccd1 vccd1 _14427_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17215_ _18289_/A vssd1 vssd1 vccd1 vccd1 _17215_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11639_ _11789_/A _11639_/B _11639_/C _11641_/C vssd1 vssd1 vccd1 vccd1 _11639_/X
+ sky130_fd_sc_hd__or4_1
X_18195_ _18195_/A vssd1 vssd1 vccd1 vccd1 _19955_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18324__A _18324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11188__A3 _11186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14358_ _14358_/A vssd1 vssd1 vccd1 vccd1 _18789_/D sky130_fd_sc_hd__clkbuf_1
X_17146_ _17146_/A _17146_/B vssd1 vssd1 vccd1 vccd1 _17149_/C sky130_fd_sc_hd__nand2_1
XFILLER_7_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13309_ _15251_/A vssd1 vssd1 vccd1 vccd1 _13309_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17077_ _17079_/A _17079_/C _17059_/X vssd1 vssd1 vccd1 vccd1 _17077_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10491__S1 _10333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14289_ _14289_/A vssd1 vssd1 vccd1 vccd1 _18759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16028_ _13309_/X _19436_/Q _16034_/S vssd1 vssd1 vccd1 vccd1 _16029_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14998__S _15000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__A2 _10687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11896__B2 _18336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__A _11464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16284__B1 _12444_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14299__A _14367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17979_ _17560_/A _17971_/Y _17978_/X _17966_/Y vssd1 vssd1 vccd1 vccd1 _17979_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_66_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19718_ _19718_/CLK _19718_/D vssd1 vssd1 vccd1 vccd1 _19718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10856__C1 _09738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19649_ _19782_/CLK _19649_/D vssd1 vssd1 vccd1 vccd1 _19649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15622__S _15622_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09402_ _19885_/Q _19884_/Q vssd1 vssd1 vccd1 vccd1 _09404_/B sky130_fd_sc_hd__nor2_1
X_09333_ _16816_/C _17346_/A vssd1 vssd1 vccd1 vccd1 _12857_/A sky130_fd_sc_hd__and2_1
XANTENNA__13270__A0 _19907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14238__S _14246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09264_ _11634_/B _09264_/B vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__nand2_2
XFILLER_166_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09195_ _09298_/A vssd1 vssd1 vccd1 vccd1 _11704_/A sky130_fd_sc_hd__inv_12
XFILLER_147_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13573__A1 _11890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10387__B2 _19912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17792__B _17792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10234__S1 _09858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16275__A0 _15738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_103_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11990_ _11990_/A _17772_/A _11990_/C _17792_/A vssd1 vssd1 vccd1 vccd1 _12104_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_91_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10941_ _11116_/A vssd1 vssd1 vccd1 vccd1 _10941_/X sky130_fd_sc_hd__buf_2
XFILLER_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13660_ _14612_/A vssd1 vssd1 vccd1 vccd1 _13660_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10872_ _18803_/Q _19138_/Q _10872_/S vssd1 vssd1 vccd1 vccd1 _10872_/X sky130_fd_sc_hd__mux2_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12611_ _12611_/A _12611_/B _12610_/X vssd1 vssd1 vccd1 vccd1 _12612_/S sky130_fd_sc_hd__or3b_2
XFILLER_25_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13591_ _13591_/A _13591_/B vssd1 vssd1 vccd1 vccd1 _13592_/B sky130_fd_sc_hd__nand2_2
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15330_ _19174_/Q _15238_/X _15334_/S vssd1 vssd1 vccd1 vccd1 _15331_/A sky130_fd_sc_hd__mux2_1
X_12542_ _19542_/Q _12122_/X _16303_/A vssd1 vssd1 vccd1 vccd1 _12542_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_157_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ _19149_/Q _15260_/X _15261_/S vssd1 vssd1 vccd1 vccd1 _15262_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15768__A _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12473_ _12473_/A vssd1 vssd1 vccd1 vccd1 _12473_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14212_ _13835_/X _18725_/Q _14218_/S vssd1 vssd1 vccd1 vccd1 _14213_/A sky130_fd_sc_hd__mux2_1
X_17000_ _17005_/C _17003_/C _16999_/Y vssd1 vssd1 vccd1 vccd1 _19757_/D sky130_fd_sc_hd__o21a_1
XANTENNA__12367__A2 _12362_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _11540_/A _11424_/B _11539_/A _11548_/C vssd1 vssd1 vccd1 vccd1 _11536_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13564__A1 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15192_ _15192_/A vssd1 vssd1 vccd1 vccd1 _19127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14143_ _14143_/A vssd1 vssd1 vccd1 vccd1 _18696_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_53_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ _11355_/A _12643_/A vssd1 vssd1 vccd1 vccd1 _11356_/B sky130_fd_sc_hd__or2_1
XFILLER_4_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10306_ _18783_/Q _19054_/Q _19278_/Q _19022_/Q _10302_/X _09817_/A vssd1 vssd1 vccd1
+ vccd1 _10306_/X sky130_fd_sc_hd__mux4_1
X_18951_ _19502_/CLK _18951_/D vssd1 vssd1 vccd1 vccd1 _18951_/Q sky130_fd_sc_hd__dfxtp_1
X_14074_ _14074_/A _14074_/B vssd1 vssd1 vccd1 vccd1 _16371_/B sky130_fd_sc_hd__or2_1
XFILLER_3_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11286_ _18572_/Q _18833_/Q _18732_/Q _19067_/Q _11280_/S _11179_/A vssd1 vssd1 vccd1
+ vccd1 _11286_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13025_ _18503_/Q _13546_/B _12707_/X _19325_/Q _13024_/X vssd1 vssd1 vccd1 vccd1
+ _13025_/X sky130_fd_sc_hd__a221o_1
XFILLER_79_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17902_ _17976_/A _17902_/B vssd1 vssd1 vccd1 vccd1 _17904_/C sky130_fd_sc_hd__nor2_1
X_10237_ _19915_/Q vssd1 vssd1 vccd1 vccd1 _10237_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11878__A1 _13172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18882_ _19564_/CLK _18882_/D vssd1 vssd1 vccd1 vccd1 _18882_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10225__S1 _09927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17833_ _17791_/X _17829_/Y _17832_/Y vssd1 vssd1 vccd1 vccd1 _17833_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10168_ _09567_/A _10167_/X _09580_/X vssd1 vssd1 vccd1 vccd1 _10168_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10440__A _10440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17764_ _17761_/X _17763_/X _17805_/S vssd1 vssd1 vccd1 vccd1 _17764_/X sky130_fd_sc_hd__mux2_2
X_14976_ _14976_/A vssd1 vssd1 vccd1 vccd1 _19027_/D sky130_fd_sc_hd__clkbuf_1
X_10099_ _19479_/Q _19317_/Q _18726_/Q _18496_/Q _11483_/S _10618_/A vssd1 vssd1 vccd1
+ vccd1 _10100_/B sky130_fd_sc_hd__mux4_1
XFILLER_47_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19503_ _19503_/CLK _19503_/D vssd1 vssd1 vccd1 vccd1 _19503_/Q sky130_fd_sc_hd__dfxtp_1
X_16715_ _16717_/B _16717_/C _16714_/Y vssd1 vssd1 vccd1 vccd1 _19676_/D sky130_fd_sc_hd__o21a_1
XFILLER_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13927_ _13927_/A vssd1 vssd1 vccd1 vccd1 _18602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13173__D input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17695_ _17702_/A _17693_/X _17694_/X vssd1 vssd1 vccd1 vccd1 _17695_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_19_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18319__A _18319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14847__A _14915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13751__A _13832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19434_ _19575_/CLK _19434_/D vssd1 vssd1 vccd1 vccd1 _19434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16646_ _16645_/A _16645_/C _19656_/Q vssd1 vssd1 vccd1 vccd1 _16647_/C sky130_fd_sc_hd__a21oi_1
X_13858_ _13926_/S vssd1 vssd1 vccd1 vccd1 _13867_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_16_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12809_ _19613_/Q _13142_/B _12801_/X _12808_/X vssd1 vssd1 vccd1 vccd1 _12813_/A
+ sky130_fd_sc_hd__o22a_2
XANTENNA__13252__A0 hold15/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19365_ _19555_/CLK _19365_/D vssd1 vssd1 vccd1 vccd1 _19365_/Q sky130_fd_sc_hd__dfxtp_1
X_16577_ _18281_/B vssd1 vssd1 vccd1 vccd1 _16577_/X sky130_fd_sc_hd__buf_2
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13789_ _13789_/A vssd1 vssd1 vccd1 vccd1 _18550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18316_ _18316_/A _18333_/B vssd1 vssd1 vccd1 vccd1 _18316_/X sky130_fd_sc_hd__or2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ _19262_/Q _15212_/X _15528_/S vssd1 vssd1 vccd1 vccd1 _15529_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11802__A1 _18319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_19296_ _19552_/CLK _19296_/D vssd1 vssd1 vccd1 vccd1 _19296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15678__A _16268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18247_ _19978_/Q _19599_/Q _18253_/S vssd1 vssd1 vccd1 vccd1 _18248_/A sky130_fd_sc_hd__mux2_1
X_15459_ _19231_/Q _15215_/X _15467_/S vssd1 vssd1 vccd1 vccd1 _15460_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13555__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18178_ _18178_/A vssd1 vssd1 vccd1 vccd1 _19947_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12814__B _12814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17129_ _19810_/Q _17128_/X _17129_/S vssd1 vssd1 vccd1 vccd1 _17130_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10615__A _10691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13307__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09951_ _18693_/Q _19188_/Q _10826_/S vssd1 vssd1 vccd1 vccd1 _09952_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09882_ _19381_/Q _18995_/Q _19445_/Q _18564_/Q _09881_/X _09874_/X vssd1 vssd1 vccd1
+ vccd1 _09883_/B sky130_fd_sc_hd__mux4_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16257__A0 _15724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10350__A _11464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09909__S1 _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17133__A _18413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10496__S _10496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10057__B1 _10056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ _20045_/Q _14074_/A vssd1 vssd1 vccd1 vccd1 _09316_/X sky130_fd_sc_hd__or2b_1
XFILLER_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09247_ _11523_/A _09269_/B _09266_/B vssd1 vssd1 vccd1 vccd1 _09263_/A sky130_fd_sc_hd__or3_1
XFILLER_166_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16183__S _16189_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14492__A input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09586__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09178_ _09271_/C vssd1 vssd1 vccd1 vccd1 _11785_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11140_ _18639_/Q _19230_/Q _19392_/Q _18607_/Q _11035_/X _11168_/A vssd1 vssd1 vccd1
+ vccd1 _11141_/B sky130_fd_sc_hd__mux4_1
XFILLER_162_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_clock clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_122_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10780__A1 _10030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput78 _12234_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[16] sky130_fd_sc_hd__buf_2
X_11071_ _09472_/A _11055_/X _11063_/X _11070_/X _11199_/A vssd1 vssd1 vccd1 vccd1
+ _11071_/X sky130_fd_sc_hd__a311o_1
XANTENNA__14431__S _14434_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12740__A _12853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput89 _12485_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[26] sky130_fd_sc_hd__buf_2
X_10022_ _18828_/Q vssd1 vssd1 vccd1 vccd1 _11283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14830_ _18401_/A vssd1 vssd1 vccd1 vccd1 _18359_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input16_A io_dbus_rdata[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14761_ _14761_/A vssd1 vssd1 vccd1 vccd1 _18935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11973_ _19585_/Q _12218_/A vssd1 vssd1 vccd1 vccd1 _11986_/A sky130_fd_sc_hd__or2_1
XFILLER_91_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16500_ _19659_/Q _19658_/Q _19660_/Q _16648_/A vssd1 vssd1 vccd1 vccd1 _16656_/A
+ sky130_fd_sc_hd__and4_1
X_13712_ _13712_/A vssd1 vssd1 vccd1 vccd1 _18530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10924_ _19364_/Q _18978_/Q _19428_/Q _18547_/Q _11493_/S _10910_/A vssd1 vssd1 vccd1
+ vccd1 _10925_/B sky130_fd_sc_hd__mux4_1
X_17480_ _12356_/A _17853_/B _17504_/S vssd1 vssd1 vccd1 vccd1 _17480_/X sky130_fd_sc_hd__mux2_1
X_14692_ _14692_/A vssd1 vssd1 vccd1 vccd1 _18900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13068__A1_N _13060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ _13471_/X _19572_/Q _16437_/S vssd1 vssd1 vccd1 vccd1 _16432_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10855_ _10052_/X _10852_/X _10854_/X vssd1 vssd1 vccd1 vccd1 _10855_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13643_ _14599_/A vssd1 vssd1 vccd1 vccd1 _13643_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19150_ _19409_/CLK _19150_/D vssd1 vssd1 vccd1 vccd1 _19150_/Q sky130_fd_sc_hd__dfxtp_1
X_13574_ _13573_/X _18502_/Q _13598_/S vssd1 vssd1 vccd1 vccd1 _13575_/A sky130_fd_sc_hd__mux2_1
X_16362_ _16361_/A _16361_/C _19955_/Q vssd1 vssd1 vccd1 vccd1 _16363_/B sky130_fd_sc_hd__o21ai_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _18773_/Q _19044_/Q _19268_/Q _19012_/Q _10048_/A _10037_/A vssd1 vssd1 vccd1
+ vccd1 _10787_/B sky130_fd_sc_hd__mux4_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _18121_/B _18101_/B vssd1 vssd1 vccd1 vccd1 _18101_/Y sky130_fd_sc_hd__nand2_1
X_12525_ _17525_/A vssd1 vssd1 vccd1 vccd1 _17538_/A sky130_fd_sc_hd__clkbuf_2
X_15313_ _15313_/A vssd1 vssd1 vccd1 vccd1 _19166_/D sky130_fd_sc_hd__clkbuf_1
X_19081_ _19305_/CLK _19081_/D vssd1 vssd1 vccd1 vccd1 _19081_/Q sky130_fd_sc_hd__dfxtp_1
X_16293_ _19530_/Q _16292_/X _16325_/S vssd1 vssd1 vccd1 vccd1 _16294_/A sky130_fd_sc_hd__mux2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10694__S1 _11371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16093__S _16095_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18032_ _18036_/A _18036_/B vssd1 vssd1 vccd1 vccd1 _18032_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15244_ _15244_/A vssd1 vssd1 vccd1 vccd1 _15244_/X sky130_fd_sc_hd__buf_2
X_12456_ _12457_/A _18058_/B vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__nand2_1
XFILLER_138_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12634__B _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ _11407_/A _11406_/Y vssd1 vssd1 vccd1 vccd1 _11408_/A sky130_fd_sc_hd__or2b_1
XFILLER_172_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15175_ _19119_/Q vssd1 vssd1 vccd1 vccd1 _15176_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12387_ _12387_/A _18023_/B vssd1 vssd1 vccd1 vccd1 _12388_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14126_ _14126_/A vssd1 vssd1 vccd1 vccd1 _18688_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output84_A _12362_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11338_ _11342_/A _11338_/B vssd1 vssd1 vccd1 vccd1 _11338_/Y sky130_fd_sc_hd__nor2_1
X_19983_ _19986_/CLK _19983_/D vssd1 vssd1 vccd1 vccd1 _19983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15437__S _15439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ _18659_/Q _13714_/X _14057_/S vssd1 vssd1 vccd1 vccd1 _14058_/A sky130_fd_sc_hd__mux2_1
X_18934_ _19485_/CLK _18934_/D vssd1 vssd1 vccd1 vccd1 _18934_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14341__S _14341_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12650__A _12650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ _11319_/A _11269_/B vssd1 vssd1 vccd1 vccd1 _11269_/X sky130_fd_sc_hd__or2_1
XFILLER_98_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13304__A4 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13008_ input1/X _12988_/X _13004_/X _13007_/X vssd1 vssd1 vccd1 vccd1 _15197_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_79_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18865_ _19727_/CLK _18865_/D vssd1 vssd1 vccd1 vccd1 _18865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17816_ _17849_/A _17820_/A _17814_/X _17815_/X vssd1 vssd1 vccd1 vccd1 _17816_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18796_ _19485_/CLK _18796_/D vssd1 vssd1 vccd1 vccd1 _18796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12276__A1 _10459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17747_ _17749_/A _17749_/B _18109_/S vssd1 vssd1 vccd1 vccd1 _17747_/X sky130_fd_sc_hd__mux2_1
X_14959_ _19020_/Q _14430_/X _14961_/S vssd1 vssd1 vccd1 vccd1 _14960_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14577__A _14676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17678_ _17677_/S _17527_/B _17587_/Y _17675_/S vssd1 vssd1 vccd1 vccd1 _17678_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14296__B _18297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19417_ _19417_/CLK _19417_/D vssd1 vssd1 vccd1 vccd1 _19417_/Q sky130_fd_sc_hd__dfxtp_1
X_16629_ _16629_/A _16629_/B _16629_/C vssd1 vssd1 vccd1 vccd1 _19650_/D sky130_fd_sc_hd__nor3_1
XANTENNA__12097__A _12097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19348_ _19876_/CLK _19348_/D vssd1 vssd1 vccd1 vccd1 _19348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19279_ _19409_/CLK _19279_/D vssd1 vssd1 vccd1 vccd1 _19279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17911__B1 _17910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14516__S _14524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13656__A _13744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14251__S _14257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09934_ _09891_/X _09923_/Y _09928_/X _09933_/Y _09741_/A vssd1 vssd1 vccd1 vccd1
+ _09934_/X sky130_fd_sc_hd__o311a_1
XFILLER_86_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09865_ _10271_/A vssd1 vssd1 vccd1 vccd1 _09868_/A sky130_fd_sc_hd__buf_2
XFILLER_131_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input8_A io_dbus_rdata[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16967__A _19748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11711__B1 _17581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _09800_/A _09796_/B vssd1 vssd1 vccd1 vccd1 _09796_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16178__S _16178_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14487__A input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _18809_/Q _19144_/Q _10640_/S vssd1 vssd1 vccd1 vccd1 _10641_/B sky130_fd_sc_hd__mux2_1
XFILLER_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10239__B _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10571_ _10571_/A _10571_/B vssd1 vssd1 vccd1 vccd1 _10571_/X sky130_fd_sc_hd__or2_1
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10676__S1 _09957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12310_ _19597_/Q vssd1 vssd1 vccd1 vccd1 _12339_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13290_ _19908_/Q _13289_/X _13430_/S vssd1 vssd1 vccd1 vccd1 _13290_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12241_ _12366_/A _12241_/B _12288_/C vssd1 vssd1 vccd1 vccd1 _12241_/X sky130_fd_sc_hd__or3_1
XFILLER_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12172_ _12172_/A _12172_/B vssd1 vssd1 vccd1 vccd1 _12172_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11123_ _10875_/X _11110_/X _11118_/X _11122_/X _11012_/A vssd1 vssd1 vccd1 vccd1
+ _11123_/X sky130_fd_sc_hd__a311o_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16980_ _19751_/Q _16984_/D _16979_/Y vssd1 vssd1 vccd1 vccd1 _19751_/D sky130_fd_sc_hd__o21a_1
XANTENNA__14161__S _14163_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12470__A _19842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11054_ _19103_/Q _18869_/Q _19551_/Q _19199_/Q _11237_/S _10083_/A vssd1 vssd1 vccd1
+ vccd1 _11055_/B sky130_fd_sc_hd__mux4_1
X_15931_ _15988_/S vssd1 vssd1 vccd1 vccd1 _15940_/S sky130_fd_sc_hd__buf_2
XFILLER_77_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10005_ _18828_/Q vssd1 vssd1 vccd1 vccd1 _10006_/A sky130_fd_sc_hd__clkbuf_4
X_18650_ _19049_/CLK _18650_/D vssd1 vssd1 vccd1 vccd1 _18650_/Q sky130_fd_sc_hd__dfxtp_1
X_15862_ _13128_/X _19362_/Q _15868_/S vssd1 vssd1 vccd1 vccd1 _15863_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17601_ _17505_/X _17527_/B _17601_/S vssd1 vssd1 vccd1 vccd1 _17601_/X sky130_fd_sc_hd__mux2_1
X_14813_ _18959_/Q _14456_/X _14819_/S vssd1 vssd1 vccd1 vccd1 _14814_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18581_ _19268_/CLK _18581_/D vssd1 vssd1 vccd1 vccd1 _18581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output122_A _12659_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15793_ _15792_/X _19346_/Q _15801_/S vssd1 vssd1 vccd1 vccd1 _15794_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17532_ _17794_/A vssd1 vssd1 vccd1 vccd1 _17533_/A sky130_fd_sc_hd__clkbuf_2
X_14744_ _18924_/Q _14462_/X _14746_/S vssd1 vssd1 vccd1 vccd1 _14745_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11956_ _11956_/A _11956_/B vssd1 vssd1 vccd1 vccd1 _11957_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17463_ _17853_/B _12356_/A _17465_/S vssd1 vssd1 vccd1 vccd1 _17463_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10907_ _18675_/Q _19170_/Q _11085_/A vssd1 vssd1 vccd1 vccd1 _10908_/A sky130_fd_sc_hd__mux2_1
X_14675_ _14675_/A vssd1 vssd1 vccd1 vccd1 _14675_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11887_ _17162_/A _11886_/X _11957_/A vssd1 vssd1 vccd1 vccd1 _11887_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19202_ _19203_/CLK _19202_/D vssd1 vssd1 vccd1 vccd1 _19202_/Q sky130_fd_sc_hd__dfxtp_1
X_16414_ _16414_/A vssd1 vssd1 vccd1 vccd1 _19564_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17501__A _17601_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10838_ _09989_/A _10837_/X _09964_/X vssd1 vssd1 vccd1 vccd1 _10838_/X sky130_fd_sc_hd__o21a_1
X_13626_ _14586_/A vssd1 vssd1 vccd1 vccd1 _13626_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17394_ _17394_/A _17394_/B _17394_/C vssd1 vssd1 vccd1 vccd1 _17396_/C sky130_fd_sc_hd__and3_1
XFILLER_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ _19391_/CLK _19133_/D vssd1 vssd1 vccd1 vccd1 _19133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16345_ _19540_/Q _16344_/X _16365_/S vssd1 vssd1 vccd1 vccd1 _16346_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11233__A2 _11219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769_ _19463_/Q _19301_/Q _18710_/Q _18480_/Q _11451_/S _10037_/X vssd1 vssd1 vccd1
+ vccd1 _10769_/X sky130_fd_sc_hd__mux4_2
X_13557_ _15298_/A vssd1 vssd1 vccd1 vccd1 _13557_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__13240__S _13278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _12520_/B _12508_/B vssd1 vssd1 vccd1 vccd1 _12509_/A sky130_fd_sc_hd__xnor2_2
X_19064_ _19288_/CLK _19064_/D vssd1 vssd1 vccd1 vccd1 _19064_/Q sky130_fd_sc_hd__dfxtp_1
X_13488_ _18496_/Q _13487_/X _13524_/S vssd1 vssd1 vccd1 vccd1 _13489_/A sky130_fd_sc_hd__mux2_1
X_16276_ _19527_/Q _16275_/X _16280_/S vssd1 vssd1 vccd1 vccd1 _16277_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18015_ _17765_/X _17847_/Y _18014_/X _17940_/X vssd1 vssd1 vccd1 vccd1 _18015_/X
+ sky130_fd_sc_hd__a211o_1
X_12439_ _12439_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _12439_/Y sky130_fd_sc_hd__nor2_2
X_15227_ _15227_/A vssd1 vssd1 vccd1 vccd1 _19138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09954__A _09954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15158_ _15158_/A vssd1 vssd1 vccd1 vccd1 _19110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11092__S1 _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14109_ _18681_/Q _13672_/X _14109_/S vssd1 vssd1 vccd1 vccd1 _14110_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13476__A _16347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15089_ _15089_/A vssd1 vssd1 vccd1 vccd1 _19077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19966_ _19966_/CLK _19966_/D vssd1 vssd1 vccd1 vccd1 _19966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15683__A1 _19897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18917_ _19504_/CLK _18917_/D vssd1 vssd1 vccd1 vccd1 _18917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12497__B2 _12496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19897_ _19963_/CLK _19897_/D vssd1 vssd1 vccd1 vccd1 _19897_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09650_ _10496_/S vssd1 vssd1 vccd1 vccd1 _09651_/A sky130_fd_sc_hd__buf_2
XFILLER_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18848_ _19306_/CLK _18848_/D vssd1 vssd1 vccd1 vccd1 _18848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_clock clock vssd1 vssd1 vccd1 vccd1 clkbuf_0_clock/X sky130_fd_sc_hd__clkbuf_16
XFILLER_83_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09581_ _09777_/A _09570_/X _09572_/X _09580_/X vssd1 vssd1 vccd1 vccd1 _09581_/X
+ sky130_fd_sc_hd__o211a_1
X_18779_ _19049_/CLK _18779_/D vssd1 vssd1 vccd1 vccd1 _18779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12249__B2 _11771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_175_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14100__A _14146_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17188__A1 _12874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14246__S _14246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13150__S _13196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_149_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17360__A1 _19887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09864__A _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10830__S1 _09970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09917_ _18659_/Q _19250_/Q _19412_/Q _18627_/Q _10245_/S _09899_/A vssd1 vssd1 vccd1
+ vccd1 _09918_/B sky130_fd_sc_hd__mux4_1
XFILLER_144_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20037_ _20052_/CLK _20037_/D vssd1 vssd1 vccd1 vccd1 _20037_/Q sky130_fd_sc_hd__dfxtp_1
X_09848_ _10264_/A vssd1 vssd1 vccd1 vccd1 _09860_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09773_/A _09778_/X _09580_/X vssd1 vssd1 vccd1 vccd1 _09779_/X sky130_fd_sc_hd__o21a_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _19960_/Q _11808_/X _11966_/A vssd1 vssd1 vccd1 vccd1 _17431_/A sky130_fd_sc_hd__mux2_2
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12884_/A vssd1 vssd1 vccd1 vccd1 _16875_/A sky130_fd_sc_hd__buf_4
XANTENNA__17179__A1 _15718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18376__B1 _18374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11741_ _11911_/A vssd1 vssd1 vccd1 vccd1 _12029_/C sky130_fd_sc_hd__clkbuf_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14460_ _18822_/Q _14459_/X _14466_/S vssd1 vssd1 vccd1 vccd1 _14461_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11672_ _11684_/A _09265_/X _11910_/A _09420_/A _17394_/A vssd1 vssd1 vccd1 vccd1
+ _11672_/X sky130_fd_sc_hd__o2111a_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10623_ _10623_/A _10623_/B _10623_/C vssd1 vssd1 vccd1 vccd1 _10623_/X sky130_fd_sc_hd__or3_2
X_13411_ _13398_/X _13409_/Y _13410_/Y vssd1 vssd1 vccd1 vccd1 _15270_/A sky130_fd_sc_hd__a21oi_4
X_14391_ _14391_/A vssd1 vssd1 vccd1 vccd1 _18800_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16130_ _13540_/X _19482_/Q _16132_/S vssd1 vssd1 vccd1 vccd1 _16131_/A sky130_fd_sc_hd__mux2_1
X_13342_ _13342_/A vssd1 vssd1 vccd1 vccd1 _13342_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ _10555_/A _12653_/B vssd1 vssd1 vccd1 vccd1 _10556_/A sky130_fd_sc_hd__and2_1
XFILLER_10_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13273_ _16278_/A _13271_/B _13038_/A vssd1 vssd1 vccd1 vccd1 _13274_/B sky130_fd_sc_hd__o21ai_1
X_16061_ _16061_/A vssd1 vssd1 vccd1 vccd1 _19451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10485_ _19373_/Q _18987_/Q _19437_/Q _18556_/Q _10439_/S _10397_/X vssd1 vssd1 vccd1
+ vccd1 _10486_/B sky130_fd_sc_hd__mux4_1
XFILLER_154_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12224_ _12196_/B _17933_/B vssd1 vssd1 vccd1 vccd1 _12225_/B sky130_fd_sc_hd__and2b_1
X_15012_ _15012_/A vssd1 vssd1 vccd1 vccd1 _19043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11074__S1 _10083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19820_ _19857_/CLK _19820_/D vssd1 vssd1 vccd1 vccd1 _19820_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_97_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12155_ _19527_/Q _12155_/B vssd1 vssd1 vccd1 vccd1 _12155_/X sky130_fd_sc_hd__or2_1
XFILLER_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11809__A _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_2_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_193_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _20048_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11106_ _11099_/Y _11101_/Y _11103_/Y _11105_/Y _10994_/X vssd1 vssd1 vccd1 vccd1
+ _11106_/X sky130_fd_sc_hd__o221a_2
X_19751_ _19756_/CLK _19751_/D vssd1 vssd1 vccd1 vccd1 _19751_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12479__A1 _10139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16963_ _19745_/Q _19744_/Q _19743_/Q _19742_/Q vssd1 vssd1 vccd1 vccd1 _16964_/B
+ sky130_fd_sc_hd__and4_1
X_12086_ _12086_/A _19589_/Q _12086_/C vssd1 vssd1 vccd1 vccd1 _12119_/B sky130_fd_sc_hd__and3_1
XFILLER_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09344__A1 _19894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18702_ _18836_/CLK _18702_/D vssd1 vssd1 vccd1 vccd1 _18702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15914_ _13540_/X _19386_/Q _15916_/S vssd1 vssd1 vccd1 vccd1 _15915_/A sky130_fd_sc_hd__mux2_1
X_11037_ _18769_/Q _19040_/Q _19264_/Q _19008_/Q _11035_/X _11168_/A vssd1 vssd1 vccd1
+ vccd1 _11037_/X sky130_fd_sc_hd__mux4_1
X_19682_ _19682_/CLK _19682_/D vssd1 vssd1 vccd1 vccd1 _19682_/Q sky130_fd_sc_hd__dfxtp_1
X_16894_ _16923_/B _16900_/D _16893_/X vssd1 vssd1 vccd1 vccd1 _19729_/D sky130_fd_sc_hd__o21ba_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18633_ _19556_/CLK _18633_/D vssd1 vssd1 vccd1 vccd1 _18633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15845_ _15845_/A vssd1 vssd1 vccd1 vccd1 _19355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18564_ _19449_/CLK _18564_/D vssd1 vssd1 vccd1 vccd1 _18564_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _18457_/Q _13577_/X _15775_/X vssd1 vssd1 vccd1 vccd1 _17209_/A sky130_fd_sc_hd__a21oi_2
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _12988_/A vssd1 vssd1 vccd1 vccd1 _12988_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12100__B1 _12376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17515_ _17888_/A vssd1 vssd1 vccd1 vccd1 _17729_/A sky130_fd_sc_hd__clkbuf_2
X_14727_ _18916_/Q _14436_/X _14735_/S vssd1 vssd1 vccd1 vccd1 _14728_/A sky130_fd_sc_hd__mux2_1
X_18495_ _19478_/CLK _18495_/D vssd1 vssd1 vccd1 vccd1 _18495_/Q sky130_fd_sc_hd__dfxtp_1
X_11939_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__or2_4
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10888__S1 _10084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15450__S _15456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_131_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19489_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17231__A _19843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10662__B1 _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17446_ _17914_/B _17960_/B _17460_/S vssd1 vssd1 vccd1 vccd1 _17446_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09949__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14658_ _14656_/X _18889_/Q _14670_/S vssd1 vssd1 vccd1 vccd1 _14659_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13609_ _14074_/B vssd1 vssd1 vccd1 vccd1 _18297_/A sky130_fd_sc_hd__inv_2
XANTENNA__14066__S _14068_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17377_ _17377_/A vssd1 vssd1 vccd1 vccd1 _19892_/D sky130_fd_sc_hd__clkbuf_1
X_14589_ _14589_/A vssd1 vssd1 vccd1 vccd1 _14589_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19116_ _19564_/CLK _19116_/D vssd1 vssd1 vccd1 vccd1 _19116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16328_ _16213_/X _16327_/Y _15795_/Y vssd1 vssd1 vccd1 vccd1 _16328_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_146_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19196_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19047_ _19366_/CLK _19047_/D vssd1 vssd1 vccd1 vccd1 _19047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16259_ _19524_/Q _16257_/X _16280_/S vssd1 vssd1 vccd1 vccd1 _16260_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12167__A0 _19971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10717__A1 _11399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10623__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19949_ _19981_/CLK _19949_/D vssd1 vssd1 vccd1 vccd1 _19949_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15625__S _15633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09702_ _10980_/A vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__buf_2
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09633_ _10339_/A vssd1 vssd1 vccd1 vccd1 _10544_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13419__A0 _19916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09564_ _09833_/A vssd1 vssd1 vccd1 vccd1 _09567_/A sky130_fd_sc_hd__buf_2
XFILLER_82_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10102__C1 _09602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09495_ _18965_/Q vssd1 vssd1 vccd1 vccd1 _11191_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17030__B1 _17021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17141__A _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14484__B _18408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10405__B1 _09696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10270_ _18816_/Q _19151_/Q _10270_/S vssd1 vssd1 vccd1 vccd1 _10271_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10169__C1 _10205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12732__B _13301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11348__B _12633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15535__S _15539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13960_ _13960_/A vssd1 vssd1 vccd1 vccd1 _18616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12911_ _12911_/A vssd1 vssd1 vccd1 vccd1 _12911_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10679__S _11429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13891_ _13913_/A vssd1 vssd1 vccd1 vccd1 _13900_/S sky130_fd_sc_hd__buf_2
XFILLER_47_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15630_ _15630_/A vssd1 vssd1 vccd1 vccd1 _19307_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12842_ _12842_/A vssd1 vssd1 vccd1 vccd1 _12842_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _19277_/Q _15260_/X _15561_/S vssd1 vssd1 vccd1 vccd1 _15562_/A sky130_fd_sc_hd__mux2_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _19808_/Q _12749_/X _12686_/Y _12772_/X vssd1 vssd1 vccd1 vccd1 _19808_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17220_/Y _19873_/Q _17302_/S vssd1 vssd1 vccd1 vccd1 _17301_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14512_/A vssd1 vssd1 vccd1 vccd1 _18835_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09769__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18280_ _19992_/Q _12825_/X _18279_/X _17243_/X vssd1 vssd1 vccd1 vccd1 _19992_/D
+ sky130_fd_sc_hd__o211a_1
X_11724_ _12610_/B _11724_/B _11724_/C _11724_/D vssd1 vssd1 vccd1 vccd1 _12598_/D
+ sky130_fd_sc_hd__or4_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _19246_/Q _15263_/X _15500_/S vssd1 vssd1 vccd1 vccd1 _15493_/A sky130_fd_sc_hd__mux2_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17231_ _19843_/Q _17240_/B vssd1 vssd1 vccd1 vccd1 _17231_/X sky130_fd_sc_hd__or2_1
X_14443_ _14647_/A vssd1 vssd1 vccd1 vccd1 _14443_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11811__B _17431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11655_ _18930_/Q vssd1 vssd1 vccd1 vccd1 _13324_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_63_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19092_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _10606_/A vssd1 vssd1 vccd1 vccd1 _10613_/A sky130_fd_sc_hd__clkbuf_2
X_17162_ _17162_/A _17197_/A vssd1 vssd1 vccd1 vccd1 _17162_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12936__A2 _09464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14374_ _18795_/Q _14369_/X _14386_/S vssd1 vssd1 vccd1 vccd1 _14375_/A sky130_fd_sc_hd__mux2_1
X_11586_ _11586_/A _11586_/B _11586_/C _11585_/X vssd1 vssd1 vccd1 vccd1 _11586_/X
+ sky130_fd_sc_hd__or4b_1
X_16113_ _13412_/X _19474_/Q _16117_/S vssd1 vssd1 vccd1 vccd1 _16114_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10537_ _10544_/A _10537_/B vssd1 vssd1 vccd1 vccd1 _10537_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_123_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13325_ _19943_/Q vssd1 vssd1 vccd1 vccd1 _16301_/B sky130_fd_sc_hd__clkbuf_2
X_17093_ _17095_/A _17095_/C _17059_/X vssd1 vssd1 vccd1 vccd1 _17093_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ _16044_/A vssd1 vssd1 vccd1 vccd1 _19443_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_78_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19317_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ _09842_/A _10465_/X _10467_/X vssd1 vssd1 vccd1 vccd1 _10468_/X sky130_fd_sc_hd__a21o_1
X_13256_ _13363_/A _13252_/X _13255_/X vssd1 vssd1 vccd1 vccd1 _13256_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__11047__S1 _10974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09565__A1 _10161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ _17338_/B _12378_/A _12207_/C _12207_/D vssd1 vssd1 vccd1 vccd1 _14477_/B
+ sky130_fd_sc_hd__nor4_4
X_13187_ _19715_/Q _13144_/S _12723_/A _19683_/Q _13186_/X vssd1 vssd1 vccd1 vccd1
+ _13187_/X sky130_fd_sc_hd__a221o_1
X_10399_ _10436_/A _10398_/X _09709_/A vssd1 vssd1 vccd1 vccd1 _10399_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19803_ _19803_/CLK _19803_/D vssd1 vssd1 vccd1 vccd1 _19803_/Q sky130_fd_sc_hd__dfxtp_1
X_12138_ _17884_/A _12195_/B vssd1 vssd1 vccd1 vccd1 _12139_/B sky130_fd_sc_hd__nor2_1
XFILLER_150_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18967__D _18967_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17995_ _17995_/A _17995_/B vssd1 vssd1 vccd1 vccd1 _17995_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11255__A1_N _12633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19734_ _19734_/CLK _19734_/D vssd1 vssd1 vccd1 vccd1 _19734_/Q sky130_fd_sc_hd__dfxtp_1
X_16946_ _16946_/A _16946_/B vssd1 vssd1 vccd1 vccd1 _16946_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17226__A _19842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12069_ _12069_/A vssd1 vssd1 vccd1 vccd1 _12376_/A sky130_fd_sc_hd__buf_2
XFILLER_78_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19665_ _19794_/CLK _19665_/D vssd1 vssd1 vccd1 vccd1 _19665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16877_ _16921_/B _16883_/D _16876_/X vssd1 vssd1 vccd1 vccd1 _19723_/D sky130_fd_sc_hd__o21ba_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18616_ _18845_/CLK _18616_/D vssd1 vssd1 vccd1 vccd1 _18616_/Q sky130_fd_sc_hd__dfxtp_1
X_15828_ _15818_/X _18465_/Q _15819_/Y _15827_/X vssd1 vssd1 vccd1 vccd1 _15828_/X
+ sky130_fd_sc_hd__a31o_2
Xclkbuf_leaf_16_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19608_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19596_ _19601_/CLK _19596_/D vssd1 vssd1 vccd1 vccd1 _19596_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_48_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18547_ _19555_/CLK _18547_/D vssd1 vssd1 vccd1 vccd1 _18547_/Q sky130_fd_sc_hd__dfxtp_1
X_15759_ _15759_/A vssd1 vssd1 vccd1 vccd1 _19340_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12624__A1 _19545_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__A _10039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09280_ _19996_/Q vssd1 vssd1 vccd1 vccd1 _15198_/B sky130_fd_sc_hd__clkinv_4
X_18478_ _19576_/CLK _18478_/D vssd1 vssd1 vccd1 vccd1 _18478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11721__B _18336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17429_ _17429_/A vssd1 vssd1 vccd1 vccd1 _17642_/B sky130_fd_sc_hd__buf_2
XFILLER_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12927__A2 _12908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11286__S1 _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13929__A _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14524__S _14524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13664__A _14615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17136__A input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__A0 _12309_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09616_ _09616_/A vssd1 vssd1 vccd1 vccd1 _09616_/X sky130_fd_sc_hd__buf_2
XFILLER_83_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09547_ _10825_/A vssd1 vssd1 vccd1 vccd1 _10734_/A sky130_fd_sc_hd__buf_4
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15090__S _15094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ _09820_/A vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10721__S0 _10644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _11440_/A _11440_/B vssd1 vssd1 vccd1 vccd1 _11440_/X sky130_fd_sc_hd__or2_1
XFILLER_11_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11371_ _11371_/A _11371_/B vssd1 vssd1 vccd1 vccd1 _11371_/X sky130_fd_sc_hd__and2_1
XANTENNA__14434__S _14434_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16215__A _16219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09890__S1 _09858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10322_ _10322_/A vssd1 vssd1 vccd1 vccd1 _10323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13110_ _13558_/S vssd1 vssd1 vccd1 vccd1 _13196_/S sky130_fd_sc_hd__buf_2
X_14090_ _18672_/Q _13634_/X _14098_/S vssd1 vssd1 vccd1 vccd1 _14091_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13041_ _19612_/Q vssd1 vssd1 vccd1 vccd1 _16518_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11359__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10253_ _19377_/Q _18991_/Q _19441_/Q _18560_/Q _09902_/S _10151_/A vssd1 vssd1 vccd1
+ vccd1 _10254_/B sky130_fd_sc_hd__mux4_1
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10184_ _10184_/A _10184_/B vssd1 vssd1 vccd1 vccd1 _10184_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18282__A2 _12946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input46_A io_ibus_inst[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16800_ _19704_/Q _16798_/B _16799_/Y vssd1 vssd1 vccd1 vccd1 _19704_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17046__A _17046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17780_ _19899_/Q _17758_/X _17779_/X vssd1 vssd1 vccd1 vccd1 _19899_/D sky130_fd_sc_hd__o21a_1
XFILLER_94_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14992_ _19034_/Q _14369_/X _15000_/S vssd1 vssd1 vccd1 vccd1 _14993_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16731_ _16731_/A _16737_/C vssd1 vssd1 vccd1 vccd1 _16731_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13943_ _13943_/A vssd1 vssd1 vccd1 vccd1 _18608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11201__S1 _09511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19450_ _19576_/CLK _19450_/D vssd1 vssd1 vccd1 vccd1 _19450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16662_ _16661_/A _16661_/C _19662_/Q vssd1 vssd1 vccd1 vccd1 _16663_/C sky130_fd_sc_hd__a21oi_1
XFILLER_62_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13874_ _13774_/X _18578_/Q _13878_/S vssd1 vssd1 vccd1 vccd1 _13875_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18401_ _18401_/A vssd1 vssd1 vccd1 vccd1 _18435_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15613_ _15659_/S vssd1 vssd1 vccd1 vccd1 _15622_/S sky130_fd_sc_hd__buf_6
X_19381_ _19571_/CLK _19381_/D vssd1 vssd1 vccd1 vccd1 _19381_/Q sky130_fd_sc_hd__dfxtp_1
X_12825_ _18323_/A vssd1 vssd1 vccd1 vccd1 _12825_/X sky130_fd_sc_hd__clkbuf_2
X_16593_ _16593_/A _16593_/B vssd1 vssd1 vccd1 vccd1 _16593_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18332_ _09394_/A _18323_/X _18331_/Y _18329_/X vssd1 vssd1 vccd1 vccd1 _20012_/D
+ sky130_fd_sc_hd__o211a_1
X_15544_ _19269_/Q _15235_/X _15550_/S vssd1 vssd1 vccd1 vccd1 _15545_/A sky130_fd_sc_hd__mux2_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12756_/A vssd1 vssd1 vccd1 vccd1 _13099_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12637__B _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _18263_/A vssd1 vssd1 vccd1 vccd1 _19985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _20029_/Q _11854_/B _11616_/A vssd1 vssd1 vccd1 vccd1 _11707_/X sky130_fd_sc_hd__o21a_1
X_15475_ _15475_/A vssd1 vssd1 vccd1 vccd1 _19238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12687_ _12687_/A vssd1 vssd1 vccd1 vccd1 _13142_/B sky130_fd_sc_hd__clkbuf_4
X_17214_ _19838_/Q _17226_/B vssd1 vssd1 vccd1 vccd1 _17214_/X sky130_fd_sc_hd__or2_1
X_14426_ _14426_/A vssd1 vssd1 vccd1 vccd1 _18811_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12909__A2 _16678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11638_ _11638_/A _11789_/B vssd1 vssd1 vccd1 vccd1 _11641_/C sky130_fd_sc_hd__or2_1
X_18194_ _19955_/Q _19987_/Q _18196_/S vssd1 vssd1 vccd1 vccd1 _18195_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13749__A _18293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17145_ _19816_/Q _17140_/X _17144_/Y vssd1 vssd1 vccd1 vccd1 _19816_/D sky130_fd_sc_hd__o21a_1
X_14357_ _18789_/Q _13723_/X _14363_/S vssd1 vssd1 vccd1 vccd1 _14358_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09946__B _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _11569_/A _11569_/B vssd1 vssd1 vccd1 vccd1 _11569_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12653__A _12657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13308_ _13060_/X _13299_/X _13302_/X _13307_/X vssd1 vssd1 vccd1 vccd1 _15251_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_171_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17076_ _19786_/Q _17072_/B _17075_/Y vssd1 vssd1 vccd1 vccd1 _19786_/D sky130_fd_sc_hd__o21a_1
X_14288_ _13841_/X _18759_/Q _14290_/S vssd1 vssd1 vccd1 vccd1 _14289_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16027_ _16027_/A vssd1 vssd1 vccd1 vccd1 _19435_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15964__A _15975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11269__A _11319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ _15238_/A vssd1 vssd1 vccd1 vccd1 _13239_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18340__A _18340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__B1 _16303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__A3 _10698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10901__A _11035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17978_ _18002_/A _17978_/B _17978_/C _17978_/D vssd1 vssd1 vccd1 vccd1 _17978_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_111_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19717_ _19721_/CLK _19717_/D vssd1 vssd1 vccd1 vccd1 _19717_/Q sky130_fd_sc_hd__dfxtp_1
X_16929_ _19739_/Q vssd1 vssd1 vccd1 vccd1 _16957_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19648_ _19783_/CLK _19648_/D vssd1 vssd1 vccd1 vccd1 _19648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09401_ _09377_/X _09401_/B _09401_/C vssd1 vssd1 vccd1 vccd1 _09401_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_53_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19579_ _19892_/CLK _19579_/D vssd1 vssd1 vccd1 vccd1 _19579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09332_ _09297_/Y _09322_/X _09325_/Y _09339_/A _12098_/A vssd1 vssd1 vccd1 vccd1
+ _17346_/A sky130_fd_sc_hd__a221o_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09263_ _09263_/A vssd1 vssd1 vccd1 vccd1 _11684_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09194_ _09275_/B _09269_/C _09275_/C vssd1 vssd1 vccd1 vccd1 _09298_/A sky130_fd_sc_hd__or3_4
XANTENNA__13659__A _15235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13573__A2 _13572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10387__A2 _10376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11179__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__A _10083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__A1 _10980_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11195__S0 _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ _18802_/Q _19137_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10871_ _11482_/A _10871_/B vssd1 vssd1 vccd1 vccd1 _10871_/X sky130_fd_sc_hd__and2_1
XFILLER_45_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_clock clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 _19998_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _12610_/A _12610_/B _12610_/C vssd1 vssd1 vccd1 vccd1 _12610_/X sky130_fd_sc_hd__or3_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13587_/X _13588_/X _13589_/Y _12770_/X _18439_/Q vssd1 vssd1 vccd1 vccd1
+ _13591_/B sky130_fd_sc_hd__a32o_4
XANTENNA__09465__B1 _09464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12541_ _11745_/X _12539_/Y _12581_/C _12120_/X vssd1 vssd1 vccd1 vccd1 _12541_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_129_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15260_ _15260_/A vssd1 vssd1 vccd1 vccd1 _15260_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15768__B _15768_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ _19603_/Q _12363_/X _12468_/X _12471_/Y vssd1 vssd1 vccd1 vccd1 _12472_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_8_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14211_ _14211_/A vssd1 vssd1 vccd1 vccd1 _18724_/D sky130_fd_sc_hd__clkbuf_1
X_11423_ _11552_/A _11554_/A _11552_/C _10241_/A _11422_/Y vssd1 vssd1 vccd1 vccd1
+ _11548_/C sky130_fd_sc_hd__a311o_1
X_15191_ _19127_/Q vssd1 vssd1 vccd1 vccd1 _15192_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_172_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14142_ _18696_/Q _13735_/X _14142_/S vssd1 vssd1 vccd1 vccd1 _14143_/A sky130_fd_sc_hd__mux2_1
X_11354_ _11160_/Y _11351_/X _11586_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11580_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ _10523_/A vssd1 vssd1 vccd1 vccd1 _10378_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18950_ _19501_/CLK _18950_/D vssd1 vssd1 vccd1 vccd1 _18950_/Q sky130_fd_sc_hd__dfxtp_1
X_11285_ _18764_/Q _19035_/Q _19259_/Q _19003_/Q _11329_/S _10978_/A vssd1 vssd1 vccd1
+ vccd1 _11285_/X sky130_fd_sc_hd__mux4_1
X_14073_ _14073_/A vssd1 vssd1 vccd1 vccd1 _18666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10236_ _10229_/Y _10231_/Y _10233_/Y _10235_/Y _09719_/X vssd1 vssd1 vccd1 vccd1
+ _10236_/X sky130_fd_sc_hd__o221a_2
XANTENNA__09782__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13024_ _19851_/Q _12842_/A _13343_/A _19818_/Q vssd1 vssd1 vccd1 vccd1 _13024_/X
+ sky130_fd_sc_hd__a22o_1
X_17901_ _17814_/X _17902_/B _17900_/X _17723_/A vssd1 vssd1 vccd1 vccd1 _17904_/B
+ sky130_fd_sc_hd__o211a_1
X_18881_ _19308_/CLK _18881_/D vssd1 vssd1 vccd1 vccd1 _18881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output152_A _12318_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17463__A0 _17853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17832_ _17832_/A _17832_/B vssd1 vssd1 vccd1 vccd1 _17832_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10167_ _18786_/Q _19057_/Q _19281_/Q _19025_/Q _09508_/A _10148_/X vssd1 vssd1 vccd1
+ vccd1 _10167_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17763_ _17762_/X _17602_/X _17930_/S vssd1 vssd1 vccd1 vccd1 _17763_/X sky130_fd_sc_hd__mux2_1
X_14975_ _19027_/Q _14452_/X _14983_/S vssd1 vssd1 vccd1 vccd1 _14976_/A sky130_fd_sc_hd__mux2_1
X_10098_ _18662_/Q _19253_/Q _19415_/Q _18630_/Q _11372_/S _09515_/A vssd1 vssd1 vccd1
+ vccd1 _10098_/X sky130_fd_sc_hd__mux4_1
XANTENNA__16816__A_N _16815_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19502_ _19502_/CLK _19502_/D vssd1 vssd1 vccd1 vccd1 _19502_/Q sky130_fd_sc_hd__dfxtp_1
X_16714_ _16717_/B _16717_/C _16667_/X vssd1 vssd1 vccd1 vccd1 _16714_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13926_ _13850_/X _18602_/Q _13926_/S vssd1 vssd1 vccd1 vccd1 _13927_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17694_ _17694_/A vssd1 vssd1 vccd1 vccd1 _17694_/X sky130_fd_sc_hd__clkbuf_2
X_19433_ _19497_/CLK _19433_/D vssd1 vssd1 vccd1 vccd1 _19433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16645_ _16645_/A _19656_/Q _16645_/C vssd1 vssd1 vccd1 vccd1 _16647_/B sky130_fd_sc_hd__and3_1
X_13857_ _13913_/A vssd1 vssd1 vccd1 vccd1 _13926_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__14339__S _14341_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12648__A _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15024__A _15046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ _19327_/Q _13154_/A _12696_/X _19820_/Q _12807_/X vssd1 vssd1 vccd1 vccd1
+ _12808_/X sky130_fd_sc_hd__a221o_1
X_19364_ _19555_/CLK _19364_/D vssd1 vssd1 vccd1 vccd1 _19364_/Q sky130_fd_sc_hd__dfxtp_1
X_16576_ _19632_/Q _16574_/B _16575_/Y vssd1 vssd1 vccd1 vccd1 _19632_/D sky130_fd_sc_hd__o21a_1
XANTENNA__13252__A1 _15736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13788_ _13787_/X _18550_/Q _13797_/S vssd1 vssd1 vccd1 vccd1 _13789_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18315_ _18335_/A vssd1 vssd1 vccd1 vccd1 _18333_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ _15527_/A vssd1 vssd1 vccd1 vccd1 _19261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12739_ _12739_/A vssd1 vssd1 vccd1 vccd1 _12853_/A sky130_fd_sc_hd__clkbuf_4
X_19295_ _19551_/CLK _19295_/D vssd1 vssd1 vccd1 vccd1 _19295_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09957__A _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18246_ _18246_/A vssd1 vssd1 vccd1 vccd1 _19977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ _15515_/S vssd1 vssd1 vccd1 vccd1 _15467_/S sky130_fd_sc_hd__buf_2
X_14409_ _18806_/Q _14408_/X _14418_/S vssd1 vssd1 vccd1 vccd1 _14410_/A sky130_fd_sc_hd__mux2_1
X_18177_ _19947_/Q _19979_/Q _18181_/S vssd1 vssd1 vccd1 vccd1 _18178_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15389_ _14596_/X _19200_/Q _15395_/S vssd1 vssd1 vccd1 vccd1 _15390_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17128_ _19806_/Q _12026_/X _12856_/B _17141_/A vssd1 vssd1 vccd1 vccd1 _17128_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17151__C1 _18412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09950_ _11481_/S vssd1 vssd1 vccd1 vccd1 _10826_/S sky130_fd_sc_hd__clkbuf_4
X_17059_ _17101_/A vssd1 vssd1 vccd1 vccd1 _17059_/X sky130_fd_sc_hd__buf_2
XANTENNA__14802__S _14808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ _10216_/S vssd1 vssd1 vccd1 vccd1 _09881_/X sky130_fd_sc_hd__clkbuf_4
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11177__S0 _11147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15633__S _15633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17757__A1 _19898_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10924__S0 _11493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09790__S0 _09724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14249__S _14257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10057__A1 _10052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16972__B _19748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09315_ _20000_/Q _20045_/Q vssd1 vssd1 vccd1 vccd1 _09315_/X sky130_fd_sc_hd__or2b_1
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10152__S1 _10196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09246_ _11634_/B vssd1 vssd1 vccd1 vccd1 _11675_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09177_ _20027_/Q vssd1 vssd1 vccd1 vccd1 _09271_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11070_ _11127_/A _11066_/X _11068_/X _11069_/X vssd1 vssd1 vccd1 vccd1 _11070_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput79 _12260_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[17] sky130_fd_sc_hd__buf_2
XFILLER_150_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10021_ _10021_/A vssd1 vssd1 vccd1 vccd1 _10021_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13328__S _13554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14760_ _18935_/Q _14379_/X _14764_/S vssd1 vssd1 vccd1 vccd1 _14761_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11972_ _11972_/A vssd1 vssd1 vccd1 vccd1 _11972_/Y sky130_fd_sc_hd__inv_4
X_13711_ _18530_/Q _13710_/X _13715_/S vssd1 vssd1 vccd1 vccd1 _13712_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10923_ _10043_/A _10905_/Y _10911_/X _10922_/Y _09737_/A vssd1 vssd1 vccd1 vccd1
+ _10923_/X sky130_fd_sc_hd__o311a_1
XANTENNA__14159__S _14163_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14691_ _18900_/Q _14385_/X _14691_/S vssd1 vssd1 vccd1 vccd1 _14692_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16430_ _16430_/A vssd1 vssd1 vccd1 vccd1 _19571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ _15222_/A vssd1 vssd1 vccd1 vccd1 _14599_/A sky130_fd_sc_hd__clkbuf_2
X_10854_ _10792_/A _10853_/X _10655_/A vssd1 vssd1 vccd1 vccd1 _10854_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13998__S _13998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15779__A _15808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16361_/A _19955_/Q _16361_/C vssd1 vssd1 vccd1 vccd1 _16367_/B sky130_fd_sc_hd__or3_1
XANTENNA__16374__S _16382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13573_ _11890_/X _13572_/X _11843_/B vssd1 vssd1 vccd1 vccd1 _13573_/X sky130_fd_sc_hd__a21bo_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10785_ _10792_/A _10785_/B vssd1 vssd1 vccd1 vccd1 _10785_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18100_ _17607_/X _18101_/B _18099_/X _17697_/X vssd1 vssd1 vccd1 vccd1 _18100_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12993__B1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15312_ _19166_/Q _15212_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _15313_/A sky130_fd_sc_hd__mux2_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19080_ _19560_/CLK _19080_/D vssd1 vssd1 vccd1 vccd1 _19080_/Q sky130_fd_sc_hd__dfxtp_1
X_12524_ _12473_/X _12667_/B _12474_/X _12523_/X vssd1 vssd1 vccd1 vccd1 _18090_/A
+ sky130_fd_sc_hd__a2bb2o_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16292_ _12741_/X _16291_/Y _16318_/S vssd1 vssd1 vccd1 vccd1 _16292_/X sky130_fd_sc_hd__mux2_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17920__A1 _17533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18031_ _18033_/B vssd1 vssd1 vccd1 vccd1 _18036_/A sky130_fd_sc_hd__inv_2
XFILLER_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15243_ _15243_/A vssd1 vssd1 vccd1 vccd1 _19143_/D sky130_fd_sc_hd__clkbuf_1
X_12455_ _12455_/A vssd1 vssd1 vccd1 vccd1 _18058_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11406_ _11406_/A _12649_/A vssd1 vssd1 vccd1 vccd1 _11406_/Y sky130_fd_sc_hd__nand2_1
X_15174_ _15174_/A vssd1 vssd1 vccd1 vccd1 _19118_/D sky130_fd_sc_hd__clkbuf_1
X_12386_ _12387_/A _18023_/B vssd1 vssd1 vccd1 vccd1 _12388_/A sky130_fd_sc_hd__and2_1
X_14125_ _18688_/Q _13702_/X _14131_/S vssd1 vssd1 vccd1 vccd1 _14126_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11337_ _19356_/Q _18970_/Q _19420_/Q _18539_/Q _11026_/S _11179_/X vssd1 vssd1 vccd1
+ vccd1 _11338_/B sky130_fd_sc_hd__mux4_1
XANTENNA__14622__S _14622_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19982_ _19986_/CLK _19982_/D vssd1 vssd1 vccd1 vccd1 _19982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14056_ _14056_/A vssd1 vssd1 vccd1 vccd1 _18658_/D sky130_fd_sc_hd__clkbuf_1
X_18933_ _19484_/CLK _18933_/D vssd1 vssd1 vccd1 vccd1 _18933_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output77_A _12204_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ _19357_/Q _18971_/Q _19421_/Q _18540_/Q _11262_/X _11113_/A vssd1 vssd1 vccd1
+ vccd1 _11269_/B sky130_fd_sc_hd__mux4_1
XFILLER_122_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12650__B _12651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _13174_/A vssd1 vssd1 vccd1 vccd1 _13007_/X sky130_fd_sc_hd__clkbuf_4
X_10219_ _10219_/A _10219_/B vssd1 vssd1 vccd1 vccd1 _10219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18864_ _19290_/CLK _18864_/D vssd1 vssd1 vccd1 vccd1 _18864_/Q sky130_fd_sc_hd__dfxtp_1
X_11199_ _11199_/A _11199_/B _11199_/C vssd1 vssd1 vccd1 vccd1 _11199_/X sky130_fd_sc_hd__or3_4
XFILLER_94_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17815_ _17815_/A _17820_/B vssd1 vssd1 vccd1 vccd1 _17815_/X sky130_fd_sc_hd__or2_1
X_18795_ _19484_/CLK _18795_/D vssd1 vssd1 vccd1 vccd1 _18795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14858__A _14915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17746_ _17749_/A _17749_/B vssd1 vssd1 vccd1 vccd1 _17746_/Y sky130_fd_sc_hd__nand2_1
X_14958_ _14958_/A vssd1 vssd1 vccd1 vccd1 _19019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _13825_/X _18594_/Q _13911_/S vssd1 vssd1 vccd1 vccd1 _13910_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17677_ _17586_/X _17589_/X _17677_/S vssd1 vssd1 vccd1 vccd1 _17677_/X sky130_fd_sc_hd__mux2_1
X_14889_ _14637_/X _18989_/Q _14889_/S vssd1 vssd1 vccd1 vccd1 _14890_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14296__C _18295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19416_ _19416_/CLK _19416_/D vssd1 vssd1 vccd1 vccd1 _19416_/Q sky130_fd_sc_hd__dfxtp_1
X_16628_ _16627_/A _16627_/C _19650_/Q vssd1 vssd1 vccd1 vccd1 _16629_/C sky130_fd_sc_hd__a21oi_1
XFILLER_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09524__S0 _09763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19347_ _19876_/CLK _19347_/D vssd1 vssd1 vccd1 vccd1 _19347_/Q sky130_fd_sc_hd__dfxtp_1
X_16559_ _16593_/A _16564_/C vssd1 vssd1 vccd1 vccd1 _16559_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14593__A _14676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12984__B1 _12593_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19278_ _19409_/CLK _19278_/D vssd1 vssd1 vccd1 vccd1 _19278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17911__A1 _11403_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18229_ _19970_/Q _12152_/A _18231_/S vssd1 vssd1 vccd1 vccd1 _18230_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_171_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12841__A _12992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09933_ _09936_/A _09930_/X _09932_/X vssd1 vssd1 vccd1 vccd1 _09933_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11398__S0 _10640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09864_ _09929_/A vssd1 vssd1 vccd1 vccd1 _10271_/A sky130_fd_sc_hd__buf_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _19384_/Q _18998_/Q _19448_/Q _18567_/Q _09726_/S _09730_/X vssd1 vssd1 vccd1
+ vccd1 _09796_/B sky130_fd_sc_hd__mux4_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13672__A _14621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15363__S _15367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_96_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16194__S _16200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14707__S _14713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18155__A1 _19969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10570_ _19499_/Q _18911_/Q _18948_/Q _18522_/Q _10560_/S _09815_/A vssd1 vssd1 vccd1
+ vccd1 _10571_/B sky130_fd_sc_hd__mux4_1
XFILLER_50_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ _20051_/Q _20050_/Q _20049_/Q vssd1 vssd1 vccd1 vccd1 _11730_/C sky130_fd_sc_hd__or3_1
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12240_ _19594_/Q _12240_/B _12240_/C vssd1 vssd1 vccd1 vccd1 _12288_/C sky130_fd_sc_hd__and3_1
XFILLER_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10738__C1 _09979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12171_ _12108_/A _12145_/A _12144_/A vssd1 vssd1 vccd1 vccd1 _12172_/B sky130_fd_sc_hd__a21oi_1
XFILLER_150_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11122_ _11117_/X _11119_/X _11121_/X _11069_/X vssd1 vssd1 vccd1 vccd1 _11122_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11389__S0 _10640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15930_ _15930_/A vssd1 vssd1 vccd1 vccd1 _19392_/D sky130_fd_sc_hd__clkbuf_1
X_11053_ _10961_/X _12639_/B _11052_/Y vssd1 vssd1 vccd1 vccd1 _11580_/A sky130_fd_sc_hd__o21bai_1
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10004_ _10847_/S vssd1 vssd1 vccd1 vccd1 _10777_/A sky130_fd_sc_hd__buf_4
XFILLER_103_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10061__S0 _10777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15861_ _15861_/A vssd1 vssd1 vccd1 vccd1 _19361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17600_ _17923_/S vssd1 vssd1 vccd1 vccd1 _17600_/X sky130_fd_sc_hd__clkbuf_2
X_14812_ _14812_/A vssd1 vssd1 vccd1 vccd1 _18958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18580_ _19288_/CLK _18580_/D vssd1 vssd1 vccd1 vccd1 _18580_/Q sky130_fd_sc_hd__dfxtp_1
X_15792_ _19915_/Q _15708_/X _16324_/A vssd1 vssd1 vccd1 vccd1 _15792_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12258__A2 _17949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17531_ _17542_/A _17721_/B _17538_/C vssd1 vssd1 vccd1 vccd1 _17794_/A sky130_fd_sc_hd__or3_1
XANTENNA__11466__B1 _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14743_ _14743_/A vssd1 vssd1 vccd1 vccd1 _18923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11955_ _11885_/B _11917_/Y _11953_/Y _11954_/Y vssd1 vssd1 vccd1 vccd1 _11956_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output115_A _12651_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__S _11306_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10906_ _11222_/S vssd1 vssd1 vccd1 vccd1 _11085_/A sky130_fd_sc_hd__clkbuf_4
X_17462_ _17462_/A vssd1 vssd1 vccd1 vccd1 _17853_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14674_ _14674_/A vssd1 vssd1 vccd1 vccd1 _18894_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13207__B2 _19524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11886_ _11917_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _11886_/X sky130_fd_sc_hd__xor2_1
XFILLER_33_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16413_ _13331_/X _19564_/Q _16415_/S vssd1 vssd1 vccd1 vccd1 _16414_/A sky130_fd_sc_hd__mux2_1
X_19201_ _19201_/CLK _19201_/D vssd1 vssd1 vccd1 vccd1 _19201_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11218__B1 _09703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13625_ _15209_/A vssd1 vssd1 vccd1 vccd1 _14586_/A sky130_fd_sc_hd__clkbuf_2
X_10837_ _19493_/Q _18905_/Q _18942_/Q _18516_/Q _09984_/X _09985_/X vssd1 vssd1 vccd1
+ vccd1 _10837_/X sky130_fd_sc_hd__mux4_2
X_17393_ _17393_/A _17393_/B vssd1 vssd1 vccd1 vccd1 _17397_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18146__A1 _19965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19132_ _19392_/CLK _19132_/D vssd1 vssd1 vccd1 vccd1 _19132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15302__A _15358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14844__C _14844_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16344_ _16213_/X _16343_/Y _15814_/Y vssd1 vssd1 vccd1 vccd1 _16344_/X sky130_fd_sc_hd__a21o_1
X_13556_ _13324_/X _13554_/X _13555_/X vssd1 vssd1 vccd1 vccd1 _15298_/A sky130_fd_sc_hd__o21a_1
X_10768_ _10768_/A _10768_/B vssd1 vssd1 vccd1 vccd1 _10768_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11233__A3 _11231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12645__B _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19063_ _19063_/CLK _19063_/D vssd1 vssd1 vccd1 vccd1 _19063_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10441__A1 _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ _12505_/Y _12485_/B _12506_/X vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__a21oi_1
XFILLER_173_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16275_ _15738_/X _16274_/Y _16318_/S vssd1 vssd1 vccd1 vccd1 _16275_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13487_ _15286_/A vssd1 vssd1 vccd1 vccd1 _13487_/X sky130_fd_sc_hd__buf_2
XFILLER_145_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10699_ _09613_/A _10687_/X _10698_/X _09996_/X _19905_/Q vssd1 vssd1 vccd1 vccd1
+ _10727_/A sky130_fd_sc_hd__a32o_4
X_18014_ _17612_/X _18011_/X _18013_/Y _17634_/X vssd1 vssd1 vccd1 vccd1 _18014_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15226_ _19138_/Q _15225_/X _15229_/S vssd1 vssd1 vccd1 vccd1 _15227_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12438_ _19601_/Q _19602_/Q _12438_/C vssd1 vssd1 vccd1 vccd1 _12465_/B sky130_fd_sc_hd__and3_1
XFILLER_173_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15448__S _15456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15157_ _19110_/Q vssd1 vssd1 vccd1 vccd1 _15158_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__17229__A _17229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12661__A _12663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12369_ _15840_/S vssd1 vssd1 vccd1 vccd1 _16303_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_5_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14108_ _14108_/A vssd1 vssd1 vccd1 vccd1 _18680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15088_ _14612_/X _19077_/Q _15094_/S vssd1 vssd1 vccd1 vccd1 _15089_/A sky130_fd_sc_hd__mux2_1
X_19965_ _19966_/CLK _19965_/D vssd1 vssd1 vccd1 vccd1 _19965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13143__B1 _13141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18916_ _19504_/CLK _18916_/D vssd1 vssd1 vccd1 vccd1 _18916_/Q sky130_fd_sc_hd__dfxtp_1
X_14039_ _14039_/A vssd1 vssd1 vccd1 vccd1 _18650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19896_ _19963_/CLK _19896_/D vssd1 vssd1 vccd1 vccd1 _19896_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14488__A1_N _17339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18847_ _19305_/CLK _18847_/D vssd1 vssd1 vccd1 vccd1 _18847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09580_ _09580_/A vssd1 vssd1 vccd1 vccd1 _09580_/X sky130_fd_sc_hd__buf_2
XFILLER_94_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18778_ _19049_/CLK _18778_/D vssd1 vssd1 vccd1 vccd1 _18778_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_118_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17729_ _17729_/A _17729_/B vssd1 vssd1 vccd1 vccd1 _17729_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10355__S1 _10440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10680__A1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14527__S _14535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15212__A _15212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12957__B1 _10727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13667__A _15241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14262__S _14268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11393__C1 _09738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12290__B _12395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09916_ _19476_/Q _19314_/Q _18723_/Q _18493_/Q _10244_/S _10148_/A vssd1 vssd1 vccd1
+ vccd1 _09916_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10091__A _10817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20036_ _20052_/CLK _20036_/D vssd1 vssd1 vccd1 vccd1 _20036_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09353__A2 _09345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ _09616_/X _09828_/X _09846_/X _09623_/X _19918_/Q vssd1 vssd1 vccd1 vccd1
+ _09947_/A sky130_fd_sc_hd__a32o_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16189__S _16189_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _19480_/Q _19318_/Q _18727_/Q _18497_/Q _09542_/S _09526_/X vssd1 vssd1 vccd1
+ vccd1 _09778_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13437__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18376__B2 _18375_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11740_/A vssd1 vssd1 vccd1 vccd1 _11740_/Y sky130_fd_sc_hd__clkinv_4
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11671_/A vssd1 vssd1 vccd1 vccd1 _11671_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18128__A1 _19957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12948__B1 _11082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13410_ input15/X _13353_/X _13354_/X vssd1 vssd1 vccd1 vccd1 _13410_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_168_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10622_ _11440_/A _10616_/X _10620_/X _10621_/X vssd1 vssd1 vccd1 vccd1 _10623_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14390_ _18800_/Q _14388_/X _14402_/S vssd1 vssd1 vccd1 vccd1 _14391_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10959__C1 _10949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13341_ _13341_/A vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _09749_/A _10542_/X _10551_/X _09756_/A _10552_/Y vssd1 vssd1 vccd1 vccd1
+ _12653_/B sky130_fd_sc_hd__o32a_4
XFILLER_10_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16060_ _13557_/X _19451_/Q _16060_/S vssd1 vssd1 vccd1 vccd1 _16061_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13272_ _19939_/Q vssd1 vssd1 vccd1 vccd1 _16278_/A sky130_fd_sc_hd__clkbuf_2
X_10484_ _09615_/A _10474_/X _10483_/X _09622_/A _19910_/Q vssd1 vssd1 vccd1 vccd1
+ _11562_/A sky130_fd_sc_hd__a32o_4
XFILLER_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15011_ _19043_/Q _14401_/X _15011_/S vssd1 vssd1 vccd1 vccd1 _15012_/A sky130_fd_sc_hd__mux2_1
X_12223_ _12272_/B vssd1 vssd1 vccd1 vccd1 _17945_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14172__S _14174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10282__S0 _10173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ _12116_/A _12148_/Y _12153_/X _11977_/X vssd1 vssd1 vccd1 vccd1 _12154_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_64_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ _10976_/X _11104_/X _10980_/X vssd1 vssd1 vccd1 vccd1 _11105_/Y sky130_fd_sc_hd__o21ai_1
X_19750_ _19756_/CLK _19750_/D vssd1 vssd1 vccd1 vccd1 _19750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14900__S _14900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16962_ _19747_/Q _16967_/C vssd1 vssd1 vccd1 vccd1 _16966_/B sky130_fd_sc_hd__nor2_1
X_12085_ _19589_/Q _12150_/B vssd1 vssd1 vccd1 vccd1 _12095_/A sky130_fd_sc_hd__or2_1
XFILLER_110_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18701_ _19196_/CLK _18701_/D vssd1 vssd1 vccd1 vccd1 _18701_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09344__A2 _09341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15913_ _15913_/A vssd1 vssd1 vccd1 vccd1 _19385_/D sky130_fd_sc_hd__clkbuf_1
X_11036_ _11283_/A vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__buf_4
X_19681_ _19769_/CLK _19681_/D vssd1 vssd1 vccd1 vccd1 _19681_/Q sky130_fd_sc_hd__dfxtp_1
X_16893_ _16923_/B _16923_/C _16896_/D _16875_/X vssd1 vssd1 vccd1 vccd1 _16893_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18632_ _19063_/CLK _18632_/D vssd1 vssd1 vccd1 vccd1 _18632_/Q sky130_fd_sc_hd__dfxtp_1
X_15844_ _15843_/X _19355_/Q _15844_/S vssd1 vssd1 vccd1 vccd1 _15845_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18563_ _19476_/CLK _18563_/D vssd1 vssd1 vccd1 vccd1 _18563_/Q sky130_fd_sc_hd__dfxtp_1
X_15775_ _18457_/Q _13370_/X _15774_/Y _13580_/X vssd1 vssd1 vccd1 vccd1 _15775_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12987_ _13173_/A _12986_/Y _18930_/Q _09325_/A vssd1 vssd1 vccd1 vccd1 _12988_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15731__S _15747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14737_/A vssd1 vssd1 vccd1 vccd1 _14735_/S sky130_fd_sc_hd__clkbuf_4
X_17514_ _17594_/A vssd1 vssd1 vccd1 vccd1 _17888_/A sky130_fd_sc_hd__clkbuf_2
X_18494_ _19481_/CLK _18494_/D vssd1 vssd1 vccd1 vccd1 _18494_/Q sky130_fd_sc_hd__dfxtp_1
X_11938_ _11938_/A _11938_/B vssd1 vssd1 vccd1 vccd1 _11939_/B sky130_fd_sc_hd__and2_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17445_ _17445_/A vssd1 vssd1 vccd1 vccd1 _17960_/B sky130_fd_sc_hd__buf_2
X_14657_ _14657_/A vssd1 vssd1 vccd1 vccd1 _14670_/S sky130_fd_sc_hd__buf_4
XFILLER_21_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11869_ _19580_/Q _19581_/Q _11792_/B _19582_/Q vssd1 vssd1 vccd1 vccd1 _11870_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12656__A _12657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12939__A0 _18319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ _14574_/A vssd1 vssd1 vccd1 vccd1 _13608_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17376_ _17376_/A _17376_/B vssd1 vssd1 vccd1 vccd1 _17377_/A sky130_fd_sc_hd__and2_1
XANTENNA__12403__A2 _12661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14588_ _14588_/A vssd1 vssd1 vccd1 vccd1 _18867_/D sky130_fd_sc_hd__clkbuf_1
X_19115_ _19470_/CLK _19115_/D vssd1 vssd1 vccd1 vccd1 _19115_/Q sky130_fd_sc_hd__dfxtp_1
X_16327_ _16332_/A _16332_/C vssd1 vssd1 vccd1 vccd1 _16327_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13539_ _13539_/A _13539_/B vssd1 vssd1 vccd1 vccd1 _15295_/A sky130_fd_sc_hd__nor2_2
XFILLER_118_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18343__A _18343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19046_ _19495_/CLK _19046_/D vssd1 vssd1 vccd1 vccd1 _19046_/Q sky130_fd_sc_hd__dfxtp_1
X_16258_ _16369_/S vssd1 vssd1 vccd1 vccd1 _16280_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12167__A1 _10672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13487__A _15286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15209_ _15209_/A vssd1 vssd1 vccd1 vccd1 _15209_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_44_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ _19508_/Q _14653_/A _16189_/S vssd1 vssd1 vccd1 vccd1 _16190_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10273__S0 _09926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15906__S _15912_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19948_ _19985_/CLK _19948_/D vssd1 vssd1 vccd1 vccd1 _19948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09904__S _09904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _18830_/Q vssd1 vssd1 vccd1 vccd1 _10980_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17406__B _17542_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19879_ _19879_/CLK _19879_/D vssd1 vssd1 vccd1 vccd1 _19879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09632_ _11460_/A vssd1 vssd1 vccd1 vccd1 _10339_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13419__A1 _12901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14111__A _14133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _10256_/A vssd1 vssd1 vccd1 vccd1 _09833_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12627__C1 _12026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18358__B2 _18357_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16369__A0 _19545_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09494_ _10166_/A vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14257__S _14257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11470__A _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11602__B1 _11598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12158__A1 _12855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15088__S _15094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12732__C _13301_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14720__S _14724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20019_ _20020_/CLK _20019_/D vssd1 vssd1 vccd1 vccd1 _20019_/Q sky130_fd_sc_hd__dfxtp_1
X_12910_ _12989_/A vssd1 vssd1 vccd1 vccd1 _13144_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13890_ _13890_/A vssd1 vssd1 vccd1 vccd1 _18585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12841_ _12992_/A vssd1 vssd1 vccd1 vccd1 _12842_/A sky130_fd_sc_hd__buf_2
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15560_/A vssd1 vssd1 vccd1 vccd1 _19276_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _17245_/S _12772_/B vssd1 vssd1 vccd1 vccd1 _12772_/X sky130_fd_sc_hd__and2_1
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _13761_/X _18835_/Q _14513_/S vssd1 vssd1 vccd1 vccd1 _14512_/A sky130_fd_sc_hd__mux2_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11723_ _18340_/A _11723_/B _20051_/Q vssd1 vssd1 vccd1 vccd1 _11724_/C sky130_fd_sc_hd__or3b_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _15502_/A vssd1 vssd1 vccd1 vccd1 _15500_/S sky130_fd_sc_hd__buf_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17230_/A vssd1 vssd1 vccd1 vccd1 _17240_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14442_/A vssd1 vssd1 vccd1 vccd1 _18816_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11654_/A vssd1 vssd1 vccd1 vccd1 _18928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ _18681_/Q _19176_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _10605_/X sky130_fd_sc_hd__mux2_1
X_17161_ _17229_/A vssd1 vssd1 vccd1 vccd1 _17197_/A sky130_fd_sc_hd__buf_2
XFILLER_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14373_ _14472_/S vssd1 vssd1 vccd1 vccd1 _14386_/S sky130_fd_sc_hd__buf_2
X_11585_ _10139_/X _10140_/B _11584_/X _11470_/Y vssd1 vssd1 vccd1 vccd1 _11585_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_10_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16382__S _16382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16112_ _16112_/A vssd1 vssd1 vccd1 vccd1 _19473_/D sky130_fd_sc_hd__clkbuf_1
X_13324_ _13324_/A vssd1 vssd1 vccd1 vccd1 _13324_/X sky130_fd_sc_hd__clkbuf_2
X_10536_ _19114_/Q _18880_/Q _19562_/Q _19210_/Q _10266_/A _10592_/A vssd1 vssd1 vccd1
+ vccd1 _10537_/B sky130_fd_sc_hd__mux4_1
XFILLER_156_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17092_ _19792_/Q _17089_/B _17091_/Y vssd1 vssd1 vccd1 vccd1 _19792_/D sky130_fd_sc_hd__o21a_1
XFILLER_127_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16043_ _13423_/X _19443_/Q _16045_/S vssd1 vssd1 vccd1 vccd1 _16044_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13255_ _13255_/A _13255_/B _13271_/B vssd1 vssd1 vccd1 vccd1 _13255_/X sky130_fd_sc_hd__or3_1
XFILLER_89_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _10294_/A _10466_/X _10523_/A vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10724__A _19905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12206_ _12584_/B vssd1 vssd1 vccd1 vccd1 _12206_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10255__S0 _09902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13186_ _19619_/Q _13204_/A _13185_/X vssd1 vssd1 vccd1 vccd1 _13186_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10398_ _18590_/Q _18851_/Q _18750_/Q _19085_/Q _10392_/S _10397_/X vssd1 vssd1 vccd1
+ vccd1 _10398_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19802_ _19803_/CLK _19802_/D vssd1 vssd1 vccd1 vccd1 _19802_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15726__S _15757_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ _12137_/A vssd1 vssd1 vccd1 vccd1 _12252_/A sky130_fd_sc_hd__buf_2
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17994_ _10411_/Y _17861_/X _17993_/X vssd1 vssd1 vccd1 vccd1 _19912_/D sky130_fd_sc_hd__a21oi_1
XFILLER_97_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09724__S _09724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19733_ _19734_/CLK _19733_/D vssd1 vssd1 vccd1 vccd1 _19733_/Q sky130_fd_sc_hd__dfxtp_1
X_16945_ _16958_/A _16945_/B vssd1 vssd1 vccd1 vccd1 _16946_/B sky130_fd_sc_hd__and2_1
X_12068_ _12045_/A _12044_/B _12137_/A vssd1 vssd1 vccd1 vccd1 _12074_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12321__B2 _12320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _19458_/Q _19296_/Q _18705_/Q _18475_/Q _11237_/S _10083_/A vssd1 vssd1 vccd1
+ vccd1 _11020_/B sky130_fd_sc_hd__mux4_1
X_19664_ _19794_/CLK _19664_/D vssd1 vssd1 vccd1 vccd1 _19664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16876_ _16921_/B _16921_/C _16880_/D _16875_/X vssd1 vssd1 vccd1 vccd1 _16876_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18615_ _19464_/CLK _18615_/D vssd1 vssd1 vccd1 vccd1 _18615_/Q sky130_fd_sc_hd__dfxtp_1
X_15827_ _18465_/Q _13502_/X _15826_/Y _13587_/A vssd1 vssd1 vccd1 vccd1 _15827_/X
+ sky130_fd_sc_hd__o211a_1
X_19595_ _19601_/CLK _19595_/D vssd1 vssd1 vccd1 vccd1 _19595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11507__S0 _11384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17242__A _19848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15758_ _15757_/X _19340_/Q _15772_/S vssd1 vssd1 vccd1 vccd1 _15759_/A sky130_fd_sc_hd__mux2_1
X_18546_ _19553_/CLK _18546_/D vssd1 vssd1 vccd1 vccd1 _18546_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14709_ _18908_/Q _14411_/X _14713_/S vssd1 vssd1 vccd1 vccd1 _14710_/A sky130_fd_sc_hd__mux2_1
X_15689_ _19898_/Q _15688_/X _15719_/S vssd1 vssd1 vccd1 vccd1 _15689_/X sky130_fd_sc_hd__mux2_1
X_18477_ _19552_/CLK _18477_/D vssd1 vssd1 vccd1 vccd1 _18477_/Q sky130_fd_sc_hd__dfxtp_1
X_17428_ _17417_/X _17425_/X _17685_/S vssd1 vssd1 vccd1 vccd1 _17428_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17359_ _11623_/Y _11621_/Y _11625_/X _18273_/S vssd1 vssd1 vccd1 vccd1 _17359_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19029_ _19285_/CLK _19029_/D vssd1 vssd1 vccd1 vccd1 _19029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13010__A _14074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14540__S _14546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09939__S0 _09653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09615_ _09615_/A vssd1 vssd1 vccd1 vccd1 _09616_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15371__S _15371_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13680__A _15251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17152__A _17152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ _11482_/A vssd1 vssd1 vccd1 vccd1 _10825_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ _10314_/A vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10721__S1 _10645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_192_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _20020_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12379__B2 _12378_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10485__S0 _10439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11370_ _18808_/Q _19143_/Q _11372_/S vssd1 vssd1 vccd1 vccd1 _11371_/B sky130_fd_sc_hd__mux2_1
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10321_ _09616_/A _10309_/X _10320_/X _09623_/A _19913_/Q vssd1 vssd1 vccd1 vccd1
+ _10363_/A sky130_fd_sc_hd__a32o_2
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13040_ _19676_/Q vssd1 vssd1 vccd1 vccd1 _16717_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10252_ _09820_/X _10243_/X _10247_/X _10251_/X _09588_/A vssd1 vssd1 vccd1 vccd1
+ _10252_/X sky130_fd_sc_hd__a311o_1
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11359__B _12647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10183_ _19379_/Q _18993_/Q _19443_/Q _18562_/Q _09723_/A _09868_/A vssd1 vssd1 vccd1
+ vccd1 _10184_/B sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_130_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19491_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17490__A1 _17488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input39_A io_ibus_inst[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ _15059_/S vssd1 vssd1 vccd1 vccd1 _15000_/S sky130_fd_sc_hd__buf_2
XFILLER_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12303__A1 _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16730_ _16740_/D vssd1 vssd1 vccd1 vccd1 _16737_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13942_ _18608_/Q _13634_/X _13950_/S vssd1 vssd1 vccd1 vccd1 _13943_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_145_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19290_/CLK sky130_fd_sc_hd__clkbuf_16
X_16661_ _16661_/A _19662_/Q _16661_/C vssd1 vssd1 vccd1 vccd1 _16663_/B sky130_fd_sc_hd__and3_1
X_13873_ _13873_/A vssd1 vssd1 vccd1 vccd1 _18577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15281__S hold9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18400_ _18426_/A _18400_/B vssd1 vssd1 vccd1 vccd1 _20035_/D sky130_fd_sc_hd__nor2_1
X_15612_ _15612_/A vssd1 vssd1 vccd1 vccd1 _19299_/D sky130_fd_sc_hd__clkbuf_1
X_12824_ _12824_/A vssd1 vssd1 vccd1 vccd1 _18323_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19380_ _19508_/CLK _19380_/D vssd1 vssd1 vccd1 vccd1 _19380_/Q sky130_fd_sc_hd__dfxtp_1
X_16592_ _19638_/Q _16597_/C vssd1 vssd1 vccd1 vccd1 _16593_/B sky130_fd_sc_hd__and2_1
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15543_ _15543_/A vssd1 vssd1 vccd1 vccd1 _19268_/D sky130_fd_sc_hd__clkbuf_1
X_18331_ _18331_/A _18331_/B vssd1 vssd1 vccd1 vccd1 _18331_/Y sky130_fd_sc_hd__nand2_1
X_12755_ _12755_/A vssd1 vssd1 vccd1 vccd1 _13560_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18262_ _19985_/Q _19606_/Q _18264_/S vssd1 vssd1 vccd1 vccd1 _18263_/A sky130_fd_sc_hd__mux2_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _20042_/Q _12935_/A _12937_/C vssd1 vssd1 vccd1 vccd1 _11706_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15474_ _19238_/Q _15238_/X _15478_/S vssd1 vssd1 vccd1 vccd1 _15475_/A sky130_fd_sc_hd__mux2_1
X_12686_ _17245_/S vssd1 vssd1 vccd1 vccd1 _12686_/Y sky130_fd_sc_hd__inv_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _18811_/Q _14424_/X _14434_/S vssd1 vssd1 vccd1 vccd1 _14426_/A sky130_fd_sc_hd__mux2_1
X_17213_ _17242_/B vssd1 vssd1 vccd1 vccd1 _17226_/B sky130_fd_sc_hd__clkbuf_1
X_11637_ _20031_/Q _20030_/Q _20029_/Q _18288_/A vssd1 vssd1 vccd1 vccd1 _11639_/C
+ sky130_fd_sc_hd__or4_1
X_18193_ _18193_/A vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__clkbuf_1
XFILLER_156_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16406__A _16428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__A _12976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17144_ _13596_/B _17140_/X _17101_/X vssd1 vssd1 vccd1 vccd1 _17144_/Y sky130_fd_sc_hd__a21oi_1
X_14356_ _14356_/A vssd1 vssd1 vccd1 vccd1 _18788_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13749__B _15198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ _11568_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11568_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12653__B _12653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13307_ input8/X _13303_/X _13306_/X vssd1 vssd1 vccd1 vccd1 _13307_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10519_ _10519_/A _10519_/B _10519_/C vssd1 vssd1 vccd1 vccd1 _10519_/X sky130_fd_sc_hd__or3_2
XFILLER_116_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17075_ _17108_/A _17079_/C vssd1 vssd1 vccd1 vccd1 _17075_/Y sky130_fd_sc_hd__nor2_1
X_14287_ _14287_/A vssd1 vssd1 vccd1 vccd1 _18758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11499_ _11510_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11499_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16026_ _13293_/X _19435_/Q _16034_/S vssd1 vssd1 vccd1 vccd1 _16027_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10228__S0 _09872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13238_ _11656_/X _13236_/X _13237_/X vssd1 vssd1 vccd1 vccd1 _15238_/A sky130_fd_sc_hd__o21a_4
XFILLER_143_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12542__A1 _19542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15456__S _15456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13169_ _19933_/Q vssd1 vssd1 vccd1 vccd1 _16248_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10553__B1 _09756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17977_ _17973_/B _17977_/B vssd1 vssd1 vccd1 vccd1 _17978_/D sky130_fd_sc_hd__and2b_1
XFILLER_84_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17671__S _17808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19716_ _19718_/CLK _19716_/D vssd1 vssd1 vccd1 vccd1 _19716_/Q sky130_fd_sc_hd__dfxtp_1
X_16928_ _19738_/Q _16955_/A _16927_/Y vssd1 vssd1 vccd1 vccd1 _19738_/D sky130_fd_sc_hd__o21a_1
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11716__C _17610_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10856__A1 _10000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19647_ _19783_/CLK _19647_/D vssd1 vssd1 vccd1 vccd1 _19647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16859_ _19718_/Q _16856_/C _16858_/Y vssd1 vssd1 vccd1 vccd1 _19718_/D sky130_fd_sc_hd__o21a_1
XFILLER_81_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14596__A _14596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09400_ _11833_/A _09394_/X _12810_/B _12687_/A _09399_/X vssd1 vssd1 vccd1 vccd1
+ _09401_/C sky130_fd_sc_hd__o311a_1
XFILLER_1_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19578_ _19592_/CLK _19578_/D vssd1 vssd1 vccd1 vccd1 _19578_/Q sky130_fd_sc_hd__dfxtp_1
X_09331_ _11690_/B _11616_/A vssd1 vssd1 vccd1 vccd1 _12098_/A sky130_fd_sc_hd__nand2_2
XANTENNA__11805__A0 _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18529_ _19377_/CLK _18529_/D vssd1 vssd1 vccd1 vccd1 _18529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11224__S _11224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ _09262_/A vssd1 vssd1 vccd1 vccd1 _17325_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14535__S _14535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ _09272_/A _09264_/B vssd1 vssd1 vccd1 vccd1 _09275_/C sky130_fd_sc_hd__or2_1
XFILLER_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09934__C1 _09741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13675__A _15247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_62_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19510_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17581__S _17581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11195__S1 _09511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_166_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10870_ _18675_/Q _19170_/Q _10872_/S vssd1 vssd1 vccd1 vccd1 _10871_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_77_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19417_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12738__B _18453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09529_ _09981_/A vssd1 vssd1 vccd1 vccd1 _09530_/A sky130_fd_sc_hd__buf_4
XANTENNA__09465__A1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12540_ _19606_/Q _12540_/B vssd1 vssd1 vccd1 vccd1 _12581_/C sky130_fd_sc_hd__and2_1
XFILLER_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _12314_/X _12469_/Y _12491_/B _12537_/A vssd1 vssd1 vccd1 vccd1 _12471_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16226__A _16226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14210_ _13831_/X _18724_/Q _14218_/S vssd1 vssd1 vccd1 vccd1 _14211_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11422_ _11550_/B vssd1 vssd1 vccd1 vccd1 _11422_/Y sky130_fd_sc_hd__inv_2
X_15190_ _15190_/A vssd1 vssd1 vccd1 vccd1 _19126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14141_ _14141_/A vssd1 vssd1 vccd1 vccd1 _18695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11353_ _10961_/X _12639_/B _11082_/X _12637_/B _11052_/Y vssd1 vssd1 vccd1 vccd1
+ _11586_/B sky130_fd_sc_hd__o221ai_1
XFILLER_152_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10783__B1 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19601_/CLK sky130_fd_sc_hd__clkbuf_16
X_10304_ _10380_/A _10304_/B vssd1 vssd1 vccd1 vccd1 _10304_/X sky130_fd_sc_hd__or2_1
XFILLER_3_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14072_ _18666_/Q _13743_/X _14072_/S vssd1 vssd1 vccd1 vccd1 _14073_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11284_ _11179_/X _11281_/Y _11283_/Y _11291_/A vssd1 vssd1 vccd1 vccd1 _11284_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12524__B2 _12523_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ _19775_/Q vssd1 vssd1 vccd1 vccd1 _17044_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17900_ _17945_/A _17903_/B _17607_/A _17899_/Y vssd1 vssd1 vccd1 vccd1 _17900_/X
+ sky130_fd_sc_hd__a211o_1
X_10235_ _09860_/A _10234_/X _09891_/X vssd1 vssd1 vccd1 vccd1 _10235_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17057__A _17066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18880_ _19306_/CLK _18880_/D vssd1 vssd1 vccd1 vccd1 _18880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17463__A1 _12356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17831_ _17829_/Y _17830_/X _18089_/S vssd1 vssd1 vccd1 vccd1 _17831_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10166_ _10166_/A _10166_/B vssd1 vssd1 vccd1 vccd1 _10166_/X sky130_fd_sc_hd__or2_1
XFILLER_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output145_A _12133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16896__A _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17491__S _17601_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17762_ _17660_/X _17658_/X _17800_/S vssd1 vssd1 vccd1 vccd1 _17762_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14974_ _14974_/A vssd1 vssd1 vccd1 vccd1 _14983_/S sky130_fd_sc_hd__buf_4
X_10097_ _10812_/S vssd1 vssd1 vccd1 vccd1 _11372_/S sky130_fd_sc_hd__buf_4
XFILLER_47_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19501_ _19501_/CLK _19501_/D vssd1 vssd1 vccd1 vccd1 _19501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10838__A1 _09989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16713_ _19675_/Q _16709_/C _16712_/Y vssd1 vssd1 vccd1 vccd1 _19675_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13925_ _13925_/A vssd1 vssd1 vccd1 vccd1 _18601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17693_ _17510_/B _17527_/B _17799_/S vssd1 vssd1 vccd1 vccd1 _17693_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12929__A _18138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13524__S _13524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19432_ _19464_/CLK _19432_/D vssd1 vssd1 vccd1 vccd1 _19432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13856_ _16134_/A _14502_/A vssd1 vssd1 vccd1 vccd1 _13913_/A sky130_fd_sc_hd__or2_4
X_16644_ _16645_/A _16645_/C _16643_/Y vssd1 vssd1 vccd1 vccd1 _19655_/D sky130_fd_sc_hd__o21a_1
XANTENNA__12648__B _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ _18505_/Q _13546_/B _13560_/A _19853_/Q _12806_/X vssd1 vssd1 vccd1 vccd1
+ _12807_/X sky130_fd_sc_hd__a221o_1
XFILLER_90_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19363_ _19553_/CLK _19363_/D vssd1 vssd1 vccd1 vccd1 _19363_/Q sky130_fd_sc_hd__dfxtp_1
X_13787_ _14612_/A vssd1 vssd1 vccd1 vccd1 _13787_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16575_ _16593_/A _16582_/C vssd1 vssd1 vccd1 vccd1 _16575_/Y sky130_fd_sc_hd__nor2_1
X_10999_ _10999_/A vssd1 vssd1 vccd1 vccd1 _11000_/S sky130_fd_sc_hd__buf_4
XFILLER_163_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18314_ _20005_/Q _18310_/X _18313_/Y _18303_/X vssd1 vssd1 vccd1 vccd1 _20005_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15526_ _19261_/Q _15209_/X _15528_/S vssd1 vssd1 vccd1 vccd1 _15527_/A sky130_fd_sc_hd__mux2_1
X_12738_ _15680_/A _18453_/Q vssd1 vssd1 vccd1 vccd1 _12738_/Y sky130_fd_sc_hd__nand2_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ _19794_/CLK _19294_/D vssd1 vssd1 vccd1 vccd1 _19294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15457_ _15457_/A vssd1 vssd1 vccd1 vccd1 _19230_/D sky130_fd_sc_hd__clkbuf_1
X_18245_ _19977_/Q _12340_/A _18253_/S vssd1 vssd1 vccd1 vccd1 _18246_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14355__S _14363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12669_ _12669_/A _12669_/B vssd1 vssd1 vccd1 vccd1 _12669_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__12664__A _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16136__A _16204_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14408_ _14612_/A vssd1 vssd1 vccd1 vccd1 _14408_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10449__S0 _10325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15388_ _15388_/A vssd1 vssd1 vccd1 vccd1 _19199_/D sky130_fd_sc_hd__clkbuf_1
X_18176_ _18176_/A vssd1 vssd1 vccd1 vccd1 _19946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11566__A2 _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14339_ _18781_/Q _13689_/X _14341_/S vssd1 vssd1 vccd1 vccd1 _14340_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15975__A _15975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17127_ _17127_/A vssd1 vssd1 vccd1 vccd1 _17141_/A sky130_fd_sc_hd__buf_2
XFILLER_143_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10184__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17058_ _19780_/Q _17055_/B _17057_/Y vssd1 vssd1 vccd1 vccd1 _19780_/D sky130_fd_sc_hd__o21a_1
XFILLER_131_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16009_ _16009_/A vssd1 vssd1 vccd1 vccd1 _19427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09880_ _09712_/A _09860_/Y _09869_/X _09879_/Y _09741_/X vssd1 vssd1 vccd1 vccd1
+ _09880_/X sky130_fd_sc_hd__o311a_1
XFILLER_131_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14090__S _14098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15914__S _15916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11177__S1 _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__B2 _10840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17757__A2 _09419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15215__A _15215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10924__S1 _10910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__S1 _09730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09314_ _12378_/A _19998_/Q vssd1 vssd1 vccd1 vccd1 _09320_/B sky130_fd_sc_hd__xor2_1
XFILLER_90_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10688__S0 _10614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__B2 _19896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09245_ _11730_/A _12595_/C _09249_/A vssd1 vssd1 vccd1 vccd1 _17382_/A sky130_fd_sc_hd__or3_1
XANTENNA__12574__A _12574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09176_ _11627_/B vssd1 vssd1 vccd1 vccd1 _11680_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10214__C1 _09605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_92_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12513__S _12562_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10020_ _18693_/Q _19188_/Q _11384_/S vssd1 vssd1 vccd1 vccd1 _10021_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12809__A2 _13142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10968__S _10968_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ _11971_/A _11971_/B vssd1 vssd1 vccd1 vccd1 _11972_/A sky130_fd_sc_hd__xor2_1
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12749__A _16939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13710_ _14650_/A vssd1 vssd1 vccd1 vccd1 _13710_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10922_ _10929_/A _10912_/X _10921_/X vssd1 vssd1 vccd1 vccd1 _10922_/Y sky130_fd_sc_hd__o21ai_1
X_14690_ _14690_/A vssd1 vssd1 vccd1 vccd1 _18899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13641_ _13641_/A vssd1 vssd1 vccd1 vccd1 _18513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10853_ _18580_/Q _18841_/Q _18740_/Q _19075_/Q _10048_/A _10037_/A vssd1 vssd1 vccd1
+ vccd1 _10853_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16360_/A vssd1 vssd1 vccd1 vccd1 _19543_/D sky130_fd_sc_hd__clkbuf_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _13568_/X _13569_/X _13571_/Y _12903_/X _18437_/Q vssd1 vssd1 vccd1 vccd1
+ _13572_/X sky130_fd_sc_hd__a32o_4
XANTENNA__12442__B1 _13591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ _18581_/Q _18842_/Q _18741_/Q _19076_/Q _10751_/S _10112_/A vssd1 vssd1 vccd1
+ vccd1 _10785_/B sky130_fd_sc_hd__mux4_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15311_ _15311_/A vssd1 vssd1 vccd1 vccd1 _19165_/D sky130_fd_sc_hd__clkbuf_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12523_ _18343_/A _12568_/B vssd1 vssd1 vccd1 vccd1 _12523_/X sky130_fd_sc_hd__or2_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16291_ _16301_/C _16291_/B vssd1 vssd1 vccd1 vccd1 _16291_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15242_ _19143_/Q _15241_/X _15245_/S vssd1 vssd1 vccd1 vccd1 _15243_/A sky130_fd_sc_hd__mux2_1
X_18030_ _19915_/Q _18019_/X _18029_/X vssd1 vssd1 vccd1 vccd1 _19915_/D sky130_fd_sc_hd__o21a_1
XFILLER_145_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12454_ _19982_/Q _09947_/A _12528_/S vssd1 vssd1 vccd1 vccd1 _12455_/A sky130_fd_sc_hd__mux2_4
XFILLER_138_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11405_ _11406_/A _12649_/A vssd1 vssd1 vccd1 vccd1 _11407_/A sky130_fd_sc_hd__nor2_1
X_15173_ _19118_/Q vssd1 vssd1 vccd1 vccd1 _15174_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__14903__S _14911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12385_ _12385_/A vssd1 vssd1 vccd1 vccd1 _18023_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14124_ _14124_/A vssd1 vssd1 vccd1 vccd1 _18687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11336_ _10980_/X _11326_/Y _11331_/X _11335_/Y _09735_/A vssd1 vssd1 vccd1 vccd1
+ _11336_/X sky130_fd_sc_hd__o311a_2
XFILLER_153_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19981_ _19981_/CLK _19981_/D vssd1 vssd1 vccd1 vccd1 _19981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14055_ _18658_/Q _13710_/X _14057_/S vssd1 vssd1 vccd1 vccd1 _14056_/A sky130_fd_sc_hd__mux2_1
X_18932_ _19892_/CLK _18932_/D vssd1 vssd1 vccd1 vccd1 _18932_/Q sky130_fd_sc_hd__dfxtp_1
X_11267_ _10875_/A _11257_/X _11261_/X _11266_/X _11199_/A vssd1 vssd1 vccd1 vccd1
+ _11267_/X sky130_fd_sc_hd__a311o_4
XFILLER_106_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13006_ _13305_/A vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10218_ _18817_/Q _19152_/Q _10218_/S vssd1 vssd1 vccd1 vccd1 _10219_/B sky130_fd_sc_hd__mux2_1
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18863_ _19480_/CLK _18863_/D vssd1 vssd1 vccd1 vccd1 _18863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11198_ _11204_/A _11195_/X _11197_/X _09574_/A vssd1 vssd1 vccd1 vccd1 _11199_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11181__B1 _10988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15734__S _15747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17814_ _17998_/A vssd1 vssd1 vccd1 vccd1 _17814_/X sky130_fd_sc_hd__buf_2
X_10149_ _19507_/Q _18919_/Q _18956_/Q _18530_/Q _10162_/S _10148_/X vssd1 vssd1 vccd1
+ vccd1 _10150_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18794_ _19954_/CLK _18794_/D vssd1 vssd1 vccd1 vccd1 _18794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17745_ _17600_/X _17744_/Y _17530_/A vssd1 vssd1 vccd1 vccd1 _17745_/Y sky130_fd_sc_hd__a21oi_2
X_14957_ _19019_/Q _14427_/X _14961_/S vssd1 vssd1 vccd1 vccd1 _14958_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12659__A _12663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15035__A _15046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ _13908_/A vssd1 vssd1 vccd1 vccd1 _18593_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11484__A1 _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17676_ _17676_/A vssd1 vssd1 vccd1 vccd1 _17676_/Y sky130_fd_sc_hd__inv_2
X_14888_ _14888_/A vssd1 vssd1 vccd1 vccd1 _18988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12378__B _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19415_ _19511_/CLK _19415_/D vssd1 vssd1 vccd1 vccd1 _19415_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16627_ _16627_/A _19650_/Q _16627_/C vssd1 vssd1 vccd1 vccd1 _16629_/B sky130_fd_sc_hd__and3_1
XFILLER_90_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13839_ _13838_/X _18566_/Q _13845_/S vssd1 vssd1 vccd1 vccd1 _13840_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09968__A _10675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19346_ _19844_/CLK _19346_/D vssd1 vssd1 vccd1 vccd1 _19346_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09524__S1 _09526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16558_ _19626_/Q _16558_/B vssd1 vssd1 vccd1 vccd1 _16564_/C sky130_fd_sc_hd__and2_1
XFILLER_148_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15509_ _19254_/Q _15289_/X _15511_/S vssd1 vssd1 vccd1 vccd1 _15510_/A sky130_fd_sc_hd__mux2_1
X_19277_ _19407_/CLK _19277_/D vssd1 vssd1 vccd1 vccd1 _19277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16489_ _12487_/A _12494_/A _12490_/Y _12494_/Y _12908_/X vssd1 vssd1 vccd1 vccd1
+ _19604_/D sky130_fd_sc_hd__a221oi_1
XANTENNA__17911__A2 _17861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18228_ _18228_/A vssd1 vssd1 vccd1 vccd1 _19969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_114_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18159_ _16278_/A _19971_/Q _18159_/S vssd1 vssd1 vccd1 vccd1 _18160_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14813__S _14819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09932_ _09884_/A _09931_/X _09891_/A vssd1 vssd1 vccd1 vccd1 _09932_/X sky130_fd_sc_hd__o21a_1
XFILLER_116_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11398__S1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20052_ _20052_/CLK _20052_/D vssd1 vssd1 vccd1 vccd1 _20052_/Q sky130_fd_sc_hd__dfxtp_1
X_09863_ _09863_/A vssd1 vssd1 vccd1 vccd1 _09863_/Y sky130_fd_sc_hd__inv_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09712_/X _09784_/Y _09789_/X _09793_/Y _09741_/X vssd1 vssd1 vccd1 vccd1
+ _09794_/X sky130_fd_sc_hd__o311a_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_39_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17160__A _17160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12975__A1 _18461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10817__A _10817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09228_ _11601_/A _09248_/B _09238_/A vssd1 vssd1 vccd1 vccd1 _09262_/A sky130_fd_sc_hd__or3_1
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10738__B1 _10737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16469__A2 _16449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ _12170_/A _12170_/B vssd1 vssd1 vccd1 vccd1 _12174_/A sky130_fd_sc_hd__and2_2
XFILLER_162_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ _11317_/A _11121_/B vssd1 vssd1 vccd1 vccd1 _11121_/X sky130_fd_sc_hd__or2_1
XANTENNA__10552__A _19909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11389__S1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11052_ _10961_/X _12639_/B _11352_/A _12638_/B vssd1 vssd1 vccd1 vccd1 _11052_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_107_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10003_ _10909_/S vssd1 vssd1 vccd1 vccd1 _10847_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__10061__S1 _10010_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15860_ _13109_/X _19361_/Q _15868_/S vssd1 vssd1 vccd1 vccd1 _15861_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input21_A io_dbus_rdata[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ _18958_/Q _14452_/X _14819_/S vssd1 vssd1 vccd1 vccd1 _14812_/A sky130_fd_sc_hd__mux2_1
X_15791_ _15806_/A _17217_/A vssd1 vssd1 vccd1 vccd1 _16324_/A sky130_fd_sc_hd__nor2_1
XFILLER_18_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11383__A _11383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11466__A1 _11460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17530_ _17530_/A _17929_/A vssd1 vssd1 vccd1 vccd1 _17530_/Y sky130_fd_sc_hd__nor2_1
X_14742_ _18923_/Q _14459_/X _14746_/S vssd1 vssd1 vccd1 vccd1 _14743_/A sky130_fd_sc_hd__mux2_1
X_11954_ _19822_/Q _13597_/A vssd1 vssd1 vccd1 vccd1 _11954_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10905_ _10929_/A _10905_/B vssd1 vssd1 vccd1 vccd1 _10905_/Y sky130_fd_sc_hd__nor2_1
X_17461_ _17458_/X _17460_/X _17500_/S vssd1 vssd1 vccd1 vccd1 _17461_/X sky130_fd_sc_hd__mux2_1
X_14673_ _14672_/X _18894_/Q _14676_/S vssd1 vssd1 vccd1 vccd1 _14674_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11885_ _11917_/B _11885_/B vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output108_A _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19200_ _19200_/CLK _19200_/D vssd1 vssd1 vccd1 vccd1 _19200_/Q sky130_fd_sc_hd__dfxtp_1
X_16412_ _16412_/A vssd1 vssd1 vccd1 vccd1 _19563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13624_ _13624_/A vssd1 vssd1 vccd1 vccd1 _18509_/D sky130_fd_sc_hd__clkbuf_1
X_10836_ _10840_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _10836_/X sky130_fd_sc_hd__or2_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17392_ _17392_/A _17392_/B _17392_/C _17392_/D vssd1 vssd1 vccd1 vccd1 _17542_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_13_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19131_ _19258_/CLK _19131_/D vssd1 vssd1 vccd1 vccd1 _19131_/Q sky130_fd_sc_hd__dfxtp_1
X_16343_ _16347_/A _16347_/C vssd1 vssd1 vccd1 vccd1 _16343_/Y sky130_fd_sc_hd__xnor2_2
X_13555_ input25/X _13303_/X _13306_/X vssd1 vssd1 vccd1 vccd1 _13555_/X sky130_fd_sc_hd__a21o_1
XFILLER_160_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ _18646_/Q _19237_/Q _19399_/Q _18614_/Q _10644_/X _10030_/A vssd1 vssd1 vccd1
+ vccd1 _10768_/B sky130_fd_sc_hd__mux4_1
XFILLER_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10727__A _10727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ _12481_/A _18068_/B vssd1 vssd1 vccd1 vccd1 _12506_/X sky130_fd_sc_hd__and2b_1
X_19062_ _19574_/CLK _19062_/D vssd1 vssd1 vccd1 vccd1 _19062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16274_ _16282_/C _16274_/B vssd1 vssd1 vccd1 vccd1 _16274_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13486_ _13007_/X _13474_/Y _13485_/X vssd1 vssd1 vccd1 vccd1 _15286_/A sky130_fd_sc_hd__o21ai_4
XFILLER_157_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10698_ _10689_/X _10693_/X _10695_/X _10697_/X _09603_/A vssd1 vssd1 vccd1 vccd1
+ _10698_/X sky130_fd_sc_hd__a221o_4
X_18013_ _17771_/X _18008_/Y _18012_/Y vssd1 vssd1 vccd1 vccd1 _18013_/Y sky130_fd_sc_hd__a21oi_1
X_15225_ _15225_/A vssd1 vssd1 vccd1 vccd1 _15225_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12437_ _12416_/A _12438_/C _19602_/Q vssd1 vssd1 vccd1 vccd1 _12439_/A sky130_fd_sc_hd__a21oi_1
XFILLER_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13391__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15156_ _15156_/A vssd1 vssd1 vccd1 vccd1 _19109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12368_ _12444_/A vssd1 vssd1 vccd1 vccd1 _15840_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12661__B _12661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14107_ _18680_/Q _13668_/X _14109_/S vssd1 vssd1 vccd1 vccd1 _14108_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11319_ _11319_/A _11319_/B vssd1 vssd1 vccd1 vccd1 _11319_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10462__A _10462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15087_ _15087_/A vssd1 vssd1 vccd1 vccd1 _19076_/D sky130_fd_sc_hd__clkbuf_1
X_19964_ _19966_/CLK _19964_/D vssd1 vssd1 vccd1 vccd1 _19964_/Q sky130_fd_sc_hd__dfxtp_1
X_12299_ _12188_/X _12656_/B _12298_/Y vssd1 vssd1 vccd1 vccd1 _17989_/B sky130_fd_sc_hd__a21o_2
XFILLER_113_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09347__B1 _19888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18915_ _19053_/CLK _18915_/D vssd1 vssd1 vccd1 vccd1 _18915_/Q sky130_fd_sc_hd__dfxtp_1
X_14038_ _18650_/Q _13676_/X _14046_/S vssd1 vssd1 vccd1 vccd1 _14039_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19895_ _19895_/CLK _19895_/D vssd1 vssd1 vccd1 vccd1 _19895_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__14869__A _14915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18846_ _19302_/CLK _18846_/D vssd1 vssd1 vccd1 vccd1 _18846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18777_ _18777_/CLK _18777_/D vssd1 vssd1 vccd1 vccd1 _18777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15989_ _15989_/A vssd1 vssd1 vccd1 vccd1 _19419_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15840__A0 _19923_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11457__A1 _11460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17728_ _17607_/X _17724_/Y _17727_/X vssd1 vssd1 vccd1 vccd1 _17728_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17899__B _17899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17659_ _17657_/X _17658_/X _17760_/S vssd1 vssd1 vccd1 vccd1 _17845_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14808__S _14808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11209__A1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19329_ _19859_/CLK _19329_/D vssd1 vssd1 vccd1 vccd1 _19329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16148__A1 _14592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10637__A _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14159__A0 _13758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13013__A _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12709__B2 _19530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10815__S0 _10617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11468__A _19922_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09915_ _10147_/A _09915_/B vssd1 vssd1 vccd1 vccd1 _09915_/X sky130_fd_sc_hd__or2_1
XFILLER_120_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09846_ _09479_/A _09831_/X _09833_/X _09845_/X _09605_/X vssd1 vssd1 vccd1 vccd1
+ _09846_/X sky130_fd_sc_hd__a311o_1
X_20035_ _20049_/CLK _20035_/D vssd1 vssd1 vccd1 vccd1 _20035_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11696__A1 _20041_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11240__S0 _11129_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09777_/X sky130_fd_sc_hd__or2_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__A2 _17412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14718__S _14724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _19578_/Q _16444_/C vssd1 vssd1 vccd1 vccd1 _11671_/A sky130_fd_sc_hd__and2_4
XFILLER_168_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10621_ _10621_/A vssd1 vssd1 vccd1 vccd1 _10621_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13340_ _19725_/Q vssd1 vssd1 vccd1 vccd1 _16922_/C sky130_fd_sc_hd__clkbuf_2
X_10552_ _19909_/Q vssd1 vssd1 vccd1 vccd1 _10552_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13858__A _13926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13271_ _19939_/Q _13271_/B vssd1 vssd1 vccd1 vccd1 _13297_/C sky130_fd_sc_hd__and2_1
X_10483_ _10314_/X _10476_/X _10478_/X _10482_/X _09604_/A vssd1 vssd1 vccd1 vccd1
+ _10483_/X sky130_fd_sc_hd__a311o_1
XFILLER_136_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15010_ _15010_/A vssd1 vssd1 vccd1 vccd1 _19042_/D sky130_fd_sc_hd__clkbuf_1
X_12222_ _12188_/X _12653_/B _12221_/Y vssd1 vssd1 vccd1 vccd1 _12272_/B sky130_fd_sc_hd__a21o_1
XANTENNA__17639__A1 _18118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10806__S0 _10081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input69_A io_irq_uart_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18300__A2 _18291_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12153_ _12153_/A _12153_/B _12153_/C _12153_/D vssd1 vssd1 vccd1 vccd1 _12153_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_64_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10282__S1 _09887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16311__A1 _19533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11104_ _18640_/Q _19231_/Q _19393_/Q _18608_/Q _11224_/S _10917_/A vssd1 vssd1 vccd1
+ vccd1 _11104_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16961_ _16967_/C _16961_/B vssd1 vssd1 vccd1 vccd1 _19746_/D sky130_fd_sc_hd__nor2_1
X_12084_ _12084_/A vssd1 vssd1 vccd1 vccd1 _12084_/Y sky130_fd_sc_hd__inv_6
XFILLER_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18700_ _19727_/CLK _18700_/D vssd1 vssd1 vccd1 vccd1 _18700_/Q sky130_fd_sc_hd__dfxtp_1
X_15912_ _13523_/X _19385_/Q _15912_/S vssd1 vssd1 vccd1 vccd1 _15913_/A sky130_fd_sc_hd__mux2_1
X_11035_ _11035_/A vssd1 vssd1 vccd1 vccd1 _11035_/X sky130_fd_sc_hd__buf_4
XFILLER_77_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18064__A1 _19918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19680_ _19769_/CLK _19680_/D vssd1 vssd1 vccd1 vccd1 _19680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16892_ _16897_/A _16892_/B _16900_/D vssd1 vssd1 vccd1 vccd1 _19728_/D sky130_fd_sc_hd__nor3_1
XFILLER_65_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18631_ _19512_/CLK _18631_/D vssd1 vssd1 vccd1 vccd1 _18631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15843_ _19924_/Q _12127_/A _13604_/B vssd1 vssd1 vccd1 vccd1 _15843_/X sky130_fd_sc_hd__a21o_1
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18562_ _19313_/CLK _18562_/D vssd1 vssd1 vccd1 vccd1 _18562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _15818_/A _18457_/Q vssd1 vssd1 vccd1 vccd1 _15774_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12986_ _13173_/B vssd1 vssd1 vccd1 vccd1 _12986_/Y sky130_fd_sc_hd__inv_2
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12100__A2 _12319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17513_ _17513_/A vssd1 vssd1 vccd1 vccd1 _17513_/Y sky130_fd_sc_hd__inv_2
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _14725_/A vssd1 vssd1 vccd1 vccd1 _18915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _19508_/CLK _18493_/D vssd1 vssd1 vccd1 vccd1 _18493_/Q sky130_fd_sc_hd__dfxtp_1
X_11937_ _11938_/A _11938_/B vssd1 vssd1 vccd1 vccd1 _11939_/A sky130_fd_sc_hd__nor2_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12937__A _18316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _17444_/A vssd1 vssd1 vccd1 vccd1 _17914_/B sky130_fd_sc_hd__buf_2
X_14656_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14656_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11868_ _19581_/Q _19582_/Q _11868_/C vssd1 vssd1 vccd1 vccd1 _11912_/B sky130_fd_sc_hd__and3_1
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12656__B _12656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18119__A2 _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12939__A1 _11808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10819_ _09475_/A _10810_/X _10814_/X _10818_/X _10834_/A vssd1 vssd1 vccd1 vccd1
+ _10819_/X sky130_fd_sc_hd__a311o_2
X_13607_ _15197_/A vssd1 vssd1 vccd1 vccd1 _14574_/A sky130_fd_sc_hd__buf_2
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17375_ _11704_/A _12824_/A _17358_/A _19892_/Q vssd1 vssd1 vccd1 vccd1 _17376_/B
+ sky130_fd_sc_hd__a22o_1
X_11799_ _11771_/X _11796_/X _11798_/X vssd1 vssd1 vccd1 vccd1 _11799_/X sky130_fd_sc_hd__a21o_4
X_14587_ _14586_/X _18867_/Q _14590_/S vssd1 vssd1 vccd1 vccd1 _14588_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10821__A_N _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19114_ _19306_/CLK _19114_/D vssd1 vssd1 vccd1 vccd1 _19114_/Q sky130_fd_sc_hd__dfxtp_1
X_16326_ _16326_/A vssd1 vssd1 vccd1 vccd1 _19536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13538_ _13337_/X _13534_/X _13537_/X vssd1 vssd1 vccd1 vccd1 _13539_/B sky130_fd_sc_hd__a21oi_2
XFILLER_158_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19045_ _19369_/CLK _19045_/D vssd1 vssd1 vccd1 vccd1 _19045_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13768__A _13851_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14363__S _14363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16257_ _15724_/X _16256_/Y _16262_/S vssd1 vssd1 vccd1 vccd1 _16257_/X sky130_fd_sc_hd__mux2_1
X_13469_ _13054_/A _13468_/X _13036_/X vssd1 vssd1 vccd1 vccd1 _13469_/X sky130_fd_sc_hd__o21a_1
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15208_ _15208_/A vssd1 vssd1 vccd1 vccd1 _19132_/D sky130_fd_sc_hd__clkbuf_1
X_16188_ _16188_/A vssd1 vssd1 vccd1 vccd1 _19507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11914__A2 _11907_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10192__A _19916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15139_ _19101_/Q vssd1 vssd1 vccd1 vccd1 _15140_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_142_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09981__A _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19947_ _19981_/CLK _19947_/D vssd1 vssd1 vccd1 vccd1 _19947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14599__A _14599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ _19483_/Q _19321_/Q _18730_/Q _18500_/Q _09655_/X _09788_/A vssd1 vssd1 vccd1
+ vccd1 _09700_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13707__S _13715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19878_ _19879_/CLK _19878_/D vssd1 vssd1 vccd1 vccd1 _19878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09631_ _10794_/A vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__buf_4
XANTENNA__12321__A1_N _12376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18829_ _19794_/CLK _18829_/D vssd1 vssd1 vccd1 vccd1 _18829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09562_ _09918_/A vssd1 vssd1 vccd1 vccd1 _10256_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09493_ _10156_/A vssd1 vssd1 vccd1 vccd1 _10166_/A sky130_fd_sc_hd__buf_2
XANTENNA__10102__A1 _09979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14538__S _14546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11470__B _12668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15369__S _15371_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14273__S _14279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13355__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10169__A1 _09479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11461__S0 _10649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11213__S0 _10968_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20018_ _20018_/CLK _20018_/D vssd1 vssd1 vccd1 vccd1 _20018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09829_ _10243_/A vssd1 vssd1 vccd1 vccd1 _10207_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15832__S _18466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12840_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12840_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12735_/X _12765_/X _12768_/Y _12770_/X _18454_/Q vssd1 vssd1 vccd1 vccd1
+ _12772_/B sky130_fd_sc_hd__a32o_4
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11722_ _20048_/Q vssd1 vssd1 vccd1 vccd1 _18340_/A sky130_fd_sc_hd__clkbuf_4
X_14510_ _14510_/A vssd1 vssd1 vccd1 vccd1 _18834_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15490_/A vssd1 vssd1 vccd1 vccd1 _19245_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _18816_/Q _14440_/X _14450_/S vssd1 vssd1 vccd1 vccd1 _14442_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _18928_/Q _11652_/X _11657_/S vssd1 vssd1 vccd1 vccd1 _11654_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13043__B1 _12756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ _10604_/A _10604_/B vssd1 vssd1 vccd1 vccd1 _10604_/X sky130_fd_sc_hd__and2_1
XANTENNA__09798__B1 _09696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14372_ _14453_/A vssd1 vssd1 vccd1 vccd1 _14472_/S sky130_fd_sc_hd__buf_6
X_17160_ _17160_/A vssd1 vssd1 vccd1 vccd1 _17160_/Y sky130_fd_sc_hd__inv_2
X_11584_ _11584_/A _11584_/B vssd1 vssd1 vccd1 vccd1 _11584_/X sky130_fd_sc_hd__and2_1
XFILLER_31_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16111_ _13393_/X _19473_/Q _16117_/S vssd1 vssd1 vccd1 vccd1 _16112_/A sky130_fd_sc_hd__mux2_1
X_13323_ _13323_/A vssd1 vssd1 vccd1 vccd1 _18486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10535_ _10534_/A _10531_/Y _10534_/Y _10339_/A vssd1 vssd1 vccd1 vccd1 _10535_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14183__S _14185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17091_ _17108_/A _17095_/C vssd1 vssd1 vccd1 vccd1 _17091_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12492__A _12492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16042_ _16042_/A vssd1 vssd1 vccd1 vccd1 _19442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_clock_A _19998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13254_ _19937_/Q _19938_/Q _13254_/C vssd1 vssd1 vccd1 vccd1 _13271_/B sky130_fd_sc_hd__and3_1
X_10466_ _18684_/Q _19179_/Q _10466_/S vssd1 vssd1 vccd1 vccd1 _10466_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12205_ _19593_/Q vssd1 vssd1 vccd1 vccd1 _12338_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10255__S1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10216__S _10216_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13185_ _19747_/Q _12912_/X _13184_/X _12917_/X vssd1 vssd1 vccd1 vccd1 _13185_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14911__S _14911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ _10592_/A vssd1 vssd1 vccd1 vccd1 _10397_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__16296__A0 _12772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19801_ _19803_/CLK _19801_/D vssd1 vssd1 vccd1 vccd1 _19801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12136_ _12136_/A vssd1 vssd1 vccd1 vccd1 _17903_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17993_ _12309_/A _17844_/X _17992_/X _17858_/X vssd1 vssd1 vccd1 vccd1 _17993_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19732_ _19734_/CLK _19732_/D vssd1 vssd1 vccd1 vccd1 _19732_/Q sky130_fd_sc_hd__dfxtp_1
X_16944_ _16941_/Y _16939_/C _16943_/X vssd1 vssd1 vccd1 vccd1 _19742_/D sky130_fd_sc_hd__a21oi_1
X_12067_ _12247_/A _12062_/X _12065_/X _12066_/X vssd1 vssd1 vccd1 vccd1 _16465_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_49_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11018_ _11274_/A vssd1 vssd1 vccd1 vccd1 _11125_/A sky130_fd_sc_hd__clkbuf_2
X_19663_ _19794_/CLK _19663_/D vssd1 vssd1 vccd1 vccd1 _19663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16875_ _16875_/A vssd1 vssd1 vccd1 vccd1 _16875_/X sky130_fd_sc_hd__buf_2
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18614_ _18777_/CLK _18614_/D vssd1 vssd1 vccd1 vccd1 _18614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15826_ _15837_/A _18465_/Q vssd1 vssd1 vccd1 vccd1 _15826_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19594_ _19594_/CLK _19594_/D vssd1 vssd1 vccd1 vccd1 _19594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18545_ _19552_/CLK _18545_/D vssd1 vssd1 vccd1 vccd1 _18545_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17242__B _17242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15757_ _19909_/Q _12741_/X _15757_/S vssd1 vssd1 vccd1 vccd1 _15757_/X sky130_fd_sc_hd__mux2_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12667__A _12669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12969_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17548__B1 _17976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14708_ _14708_/A vssd1 vssd1 vccd1 vccd1 _18907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18476_ _19553_/CLK _18476_/D vssd1 vssd1 vccd1 vccd1 _18476_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15688_ _13568_/X _15686_/X _15687_/Y _12903_/X _18442_/Q vssd1 vssd1 vccd1 vccd1
+ _15688_/X sky130_fd_sc_hd__a32o_4
XANTENNA__16220__B1 _16219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17427_ _17677_/S vssd1 vssd1 vccd1 vccd1 _17685_/S sky130_fd_sc_hd__clkbuf_2
X_14639_ _14639_/A vssd1 vssd1 vccd1 vccd1 _18883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17358_ _17358_/A vssd1 vssd1 vccd1 vccd1 _17358_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16309_ _16321_/D _16308_/Y _16303_/X vssd1 vssd1 vccd1 vccd1 _16309_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_174_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17289_ _15764_/Y _19868_/Q _17291_/S vssd1 vssd1 vccd1 vccd1 _17290_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19028_ _19478_/CLK _19028_/D vssd1 vssd1 vccd1 vccd1 _19028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14821__S _14823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16287__A0 _19529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09939__S1 _09929_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14122__A _14133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09614_ _09614_/A vssd1 vssd1 vccd1 vccd1 _09615_/A sky130_fd_sc_hd__buf_4
XANTENNA__16975__C _19748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09545_ _11190_/A vssd1 vssd1 vccd1 vccd1 _11482_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14268__S _14268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09476_ _09476_/A vssd1 vssd1 vccd1 vccd1 _10314_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16211__A0 _19516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10097__A _10812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13900__S _13900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09875__S0 _09872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15099__S _15105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10485__S1 _10397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10320_ _10311_/X _10315_/X _10317_/X _10319_/X _09605_/A vssd1 vssd1 vccd1 vccd1
+ _10320_/X sky130_fd_sc_hd__a221o_1
XFILLER_4_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_162_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10251_ _10147_/A _10248_/X _10250_/X _09580_/A vssd1 vssd1 vccd1 vccd1 _10251_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14731__S _14735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10182_ _09712_/A _10172_/Y _10177_/X _10181_/Y _09741_/X vssd1 vssd1 vccd1 vccd1
+ _10182_/X sky130_fd_sc_hd__o311a_1
XANTENNA__13855__B _18297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14990_ _15046_/A vssd1 vssd1 vccd1 vccd1 _15059_/S sky130_fd_sc_hd__buf_6
X_13941_ _13998_/S vssd1 vssd1 vccd1 vccd1 _13950_/S sky130_fd_sc_hd__buf_2
XFILLER_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16660_ _16661_/A _16661_/C _16659_/Y vssd1 vssd1 vccd1 vccd1 _19661_/D sky130_fd_sc_hd__o21a_1
XFILLER_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13872_ _13771_/X _18577_/Q _13878_/S vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15611_ _14605_/X _19299_/Q _15611_/S vssd1 vssd1 vccd1 vccd1 _15612_/A sky130_fd_sc_hd__mux2_1
X_12823_ _17322_/A vssd1 vssd1 vccd1 vccd1 _12824_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16591_ _16629_/A _16591_/B _16597_/C vssd1 vssd1 vccd1 vccd1 _19637_/D sky130_fd_sc_hd__nor3_1
XANTENNA__13264__B1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18330_ _13136_/B _18323_/X _18328_/X _18329_/X vssd1 vssd1 vccd1 vccd1 _20011_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_87_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15542_ _19268_/Q _15231_/X _15550_/S vssd1 vssd1 vccd1 vccd1 _15543_/A sky130_fd_sc_hd__mux2_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _19659_/Q _12752_/X _12753_/X _19791_/Q vssd1 vssd1 vccd1 vccd1 _13316_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11853_/S vssd1 vssd1 vccd1 vccd1 _12937_/C sky130_fd_sc_hd__clkbuf_4
X_18261_ _18261_/A vssd1 vssd1 vccd1 vccd1 _19984_/D sky130_fd_sc_hd__clkbuf_1
X_15473_ _15473_/A vssd1 vssd1 vccd1 vccd1 _19237_/D sky130_fd_sc_hd__clkbuf_1
X_12685_ _12791_/B vssd1 vssd1 vccd1 vccd1 _17245_/S sky130_fd_sc_hd__buf_2
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13810__S _13813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17212_ _17229_/A vssd1 vssd1 vccd1 vccd1 _17212_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14424_ _14628_/A vssd1 vssd1 vccd1 vccd1 _14424_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11636_ _11636_/A _17392_/B _11636_/C _17395_/B vssd1 vssd1 vccd1 vccd1 _11651_/B
+ sky130_fd_sc_hd__or4_1
X_18192_ _16361_/A _19986_/Q _18192_/S vssd1 vssd1 vccd1 vccd1 _18193_/A sky130_fd_sc_hd__mux2_1
X_17143_ _19815_/Q _17140_/X _17141_/X _17142_/X vssd1 vssd1 vccd1 vccd1 _19815_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14355_ _18788_/Q _13718_/X _14363_/S vssd1 vssd1 vccd1 vccd1 _14356_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11567_ _11567_/A vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__inv_2
XFILLER_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13319__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ _10523_/A _10515_/X _10517_/X _10307_/A vssd1 vssd1 vccd1 vccd1 _10519_/C
+ sky130_fd_sc_hd__o211a_1
X_13306_ _13354_/A vssd1 vssd1 vccd1 vccd1 _13306_/X sky130_fd_sc_hd__clkbuf_2
X_14286_ _13838_/X _18758_/Q _14290_/S vssd1 vssd1 vccd1 vccd1 _14287_/A sky130_fd_sc_hd__mux2_1
X_17074_ _17074_/A vssd1 vssd1 vccd1 vccd1 _17079_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11498_ _19128_/Q _18894_/Q _19576_/Q _19224_/Q _10119_/X _10054_/A vssd1 vssd1 vccd1
+ vccd1 _11499_/B sky130_fd_sc_hd__mux4_1
XFILLER_109_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16025_ _16047_/A vssd1 vssd1 vccd1 vccd1 _16034_/S sky130_fd_sc_hd__buf_2
X_13237_ input4/X _13172_/X _13175_/X vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__a21o_1
XFILLER_171_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10228__S1 _09874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10449_ _19502_/Q _18914_/Q _18951_/Q _18525_/Q _10325_/X _10497_/A vssd1 vssd1 vccd1
+ vccd1 _10449_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16269__A0 _12874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13168_ _19933_/Q _13170_/B vssd1 vssd1 vccd1 vccd1 _13214_/C sky130_fd_sc_hd__and2_1
XFILLER_151_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10553__A1 _09749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _12119_/A _12119_/B vssd1 vssd1 vccd1 vccd1 _12178_/C sky130_fd_sc_hd__and2_1
XANTENNA__10470__A _11428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13099_ _13099_/A vssd1 vssd1 vccd1 vccd1 _13099_/X sky130_fd_sc_hd__buf_2
X_17976_ _17976_/A _17976_/B vssd1 vssd1 vccd1 vccd1 _17978_/C sky130_fd_sc_hd__nor2_1
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19715_ _19718_/CLK _19715_/D vssd1 vssd1 vccd1 vccd1 _19715_/Q sky130_fd_sc_hd__dfxtp_1
X_16927_ _16946_/A _16959_/B vssd1 vssd1 vccd1 vccd1 _16927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17769__A0 _17772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18349__A _18349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15472__S _15478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19646_ _19783_/CLK _19646_/D vssd1 vssd1 vccd1 vccd1 _19646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16858_ _16946_/A _16870_/D vssd1 vssd1 vccd1 vccd1 _16858_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15809_ _15807_/X _19349_/Q _15835_/S vssd1 vssd1 vccd1 vccd1 _15810_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19577_ _19577_/CLK _19577_/D vssd1 vssd1 vccd1 vccd1 _19577_/Q sky130_fd_sc_hd__dfxtp_1
X_16789_ _19700_/Q _16790_/C _19701_/Q vssd1 vssd1 vccd1 vccd1 _16791_/B sky130_fd_sc_hd__a21oi_1
XFILLER_80_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09330_ _11785_/A _11787_/A _11682_/B vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__nand3b_4
X_18528_ _19504_/CLK _18528_/D vssd1 vssd1 vccd1 vccd1 _18528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09261_ _11730_/A _11789_/A _11663_/B vssd1 vssd1 vccd1 vccd1 _09420_/A sky130_fd_sc_hd__a21o_2
X_18459_ _19985_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_166_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13720__S _13736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09192_ _20034_/Q vssd1 vssd1 vccd1 vccd1 _09264_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12781__A2 _12677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15647__S _15655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14551__S _14557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17147__B _17346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15382__S _15384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_109_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13246__B1 _13205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _11259_/S vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__buf_4
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10155__S0 _10244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _15662_/B _11952_/D vssd1 vssd1 vccd1 vccd1 _14477_/A sky130_fd_sc_hd__or2b_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17610__B _17610_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12470_ _19842_/Q _17223_/A _12470_/C vssd1 vssd1 vccd1 vccd1 _12491_/B sky130_fd_sc_hd__and3_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11421_ _11421_/A _12661_/B vssd1 vssd1 vccd1 vccd1 _11550_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12221__A1 _12935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10555__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140_ _18695_/Q _13731_/X _14142_/S vssd1 vssd1 vccd1 vccd1 _14141_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11352_ _11352_/A _12638_/B vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__nor2_1
XFILLER_165_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10303_ _18591_/Q _18852_/Q _18751_/Q _19086_/Q _10302_/X _09817_/A vssd1 vssd1 vccd1
+ vccd1 _10304_/B sky130_fd_sc_hd__mux4_1
XANTENNA__15557__S _15561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14071_ _14071_/A vssd1 vssd1 vccd1 vccd1 _18665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11283_ _11283_/A _11283_/B vssd1 vssd1 vccd1 vccd1 _11283_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17338__A _17338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13022_ _19643_/Q vssd1 vssd1 vccd1 vccd1 _16609_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10234_ _19474_/Q _19312_/Q _18721_/Q _18491_/Q _10175_/S _09858_/X vssd1 vssd1 vccd1
+ vccd1 _10234_/X sky130_fd_sc_hd__mux4_1
XANTENNA_input51_A io_ibus_inst[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17830_ _17832_/A _17832_/B _18077_/S vssd1 vssd1 vccd1 vccd1 _17830_/X sky130_fd_sc_hd__mux2_1
X_10165_ _18594_/Q _18855_/Q _18754_/Q _19089_/Q _09508_/A _10148_/X vssd1 vssd1 vccd1
+ vccd1 _10166_/B sky130_fd_sc_hd__mux4_2
XFILLER_117_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17761_ _17759_/X _17760_/X _17930_/S vssd1 vssd1 vccd1 vccd1 _17761_/X sky130_fd_sc_hd__mux2_1
X_10096_ _10630_/A _10096_/B vssd1 vssd1 vccd1 vccd1 _10096_/X sky130_fd_sc_hd__or2_1
X_14973_ _14973_/A vssd1 vssd1 vccd1 vccd1 _19026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19500_ _19500_/CLK _19500_/D vssd1 vssd1 vccd1 vccd1 _19500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16712_ _16731_/A _16717_/C vssd1 vssd1 vccd1 vccd1 _16712_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17073__A _17073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13924_ _13847_/X _18601_/Q _13926_/S vssd1 vssd1 vccd1 vccd1 _13925_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17692_ _17922_/S vssd1 vssd1 vccd1 vccd1 _17702_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19431_ _19431_/CLK _19431_/D vssd1 vssd1 vccd1 vccd1 _19431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16643_ _16645_/A _16645_/C _16624_/X vssd1 vssd1 vccd1 vccd1 _16643_/Y sky130_fd_sc_hd__a21oi_1
X_13855_ _15061_/A _18297_/A _14844_/C _14844_/D vssd1 vssd1 vccd1 vccd1 _14502_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ _19816_/Q _17140_/C _12804_/Y _19741_/Q _12805_/Y vssd1 vssd1 vccd1 vccd1
+ _12806_/X sky130_fd_sc_hd__a221o_1
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19362_ _19552_/CLK _19362_/D vssd1 vssd1 vccd1 vccd1 _19362_/Q sky130_fd_sc_hd__dfxtp_1
X_16574_ _19632_/Q _16574_/B vssd1 vssd1 vccd1 vccd1 _16582_/C sky130_fd_sc_hd__and2_1
XFILLER_34_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13786_ _13786_/A vssd1 vssd1 vccd1 vccd1 _18549_/D sky130_fd_sc_hd__clkbuf_1
X_10998_ _11002_/A vssd1 vssd1 vccd1 vccd1 _10999_/A sky130_fd_sc_hd__buf_4
XFILLER_62_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18313_ _18313_/A _18331_/B vssd1 vssd1 vccd1 vccd1 _18313_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15525_ _15525_/A vssd1 vssd1 vccd1 vccd1 _19260_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _15702_/A vssd1 vssd1 vccd1 vccd1 _15680_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19293_ _19293_/CLK _19293_/D vssd1 vssd1 vccd1 vccd1 _19293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16417__A _16428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18255_/A vssd1 vssd1 vccd1 vccd1 _18253_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_148_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15456_ _19230_/Q _15212_/X _15456_/S vssd1 vssd1 vccd1 vccd1 _15457_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12668_ _12669_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _12668_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09839__S0 _10160_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14407_ _14407_/A vssd1 vssd1 vccd1 vccd1 _18805_/D sky130_fd_sc_hd__clkbuf_1
X_11619_ _11619_/A _11690_/B vssd1 vssd1 vccd1 vccd1 _11910_/A sky130_fd_sc_hd__and2_2
X_18175_ _16317_/A _19978_/Q _18181_/S vssd1 vssd1 vccd1 vccd1 _18176_/A sky130_fd_sc_hd__mux2_1
X_15387_ _14592_/X _19199_/Q _15395_/S vssd1 vssd1 vccd1 vccd1 _15388_/A sky130_fd_sc_hd__mux2_1
X_12599_ _12599_/A _17391_/A _12598_/X vssd1 vssd1 vccd1 vccd1 _12609_/B sky130_fd_sc_hd__or3b_1
XANTENNA__11060__S _11114_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17126_ _16708_/B _17123_/B _17125_/Y vssd1 vssd1 vccd1 vccd1 _19805_/D sky130_fd_sc_hd__o21a_1
X_14338_ _14338_/A vssd1 vssd1 vccd1 vccd1 _18780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17151__A1 _13572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17248__A _17304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17057_ _17066_/A _17062_/C vssd1 vssd1 vccd1 vccd1 _17057_/Y sky130_fd_sc_hd__nor2_1
X_14269_ _14269_/A vssd1 vssd1 vccd1 vccd1 _18750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16008_ _13149_/X _19427_/Q _16012_/S vssd1 vssd1 vccd1 vccd1 _16009_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15991__A _16047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_191_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19745_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17959_ _17964_/B _17960_/B vssd1 vssd1 vccd1 vccd1 _17963_/B sky130_fd_sc_hd__and2b_1
XFILLER_39_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13715__S _13715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_110_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19629_ _19759_/CLK _19629_/D vssd1 vssd1 vccd1 vccd1 _19629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11235__S _11306_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13016__A _14148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09313_ _20043_/Q vssd1 vssd1 vccd1 vccd1 _12378_/A sky130_fd_sc_hd__buf_2
XANTENNA__12987__C1 _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11254__A2 _11244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14546__S _14546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12855__A _12855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15231__A _15231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09244_ _09244_/A vssd1 vssd1 vccd1 vccd1 _12595_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ _18279_/A _18276_/A _09328_/C _09328_/D vssd1 vssd1 vccd1 vccd1 _11627_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_108_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17678__C1 _17675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_144_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19727_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_35_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11714__B1 _11764_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__B _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_159_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19783_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16001__S _16001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14310__A _14367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ _11932_/A _17772_/B _11939_/B vssd1 vssd1 vccd1 vccd1 _11971_/B sky130_fd_sc_hd__a21oi_1
XFILLER_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10921_ _10051_/A _10918_/X _10920_/X vssd1 vssd1 vccd1 vccd1 _10921_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10852_ _18772_/Q _19043_/Q _19267_/Q _19011_/Q _10053_/X _10054_/X vssd1 vssd1 vccd1
+ vccd1 _10852_/X sky130_fd_sc_hd__mux4_2
XFILLER_60_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13640_ _18513_/Q _13639_/X _13652_/S vssd1 vssd1 vccd1 vccd1 _13641_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14839__A1_N _18319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10778_/X _10780_/Y _10043_/X _10782_/Y vssd1 vssd1 vccd1 vccd1 _10783_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12549__A2_N _12668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13571_ _15737_/A _18437_/Q vssd1 vssd1 vccd1 vccd1 _13571_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12442__A1 _19538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12765__A _18454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _19165_/Q _15209_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _15311_/A sky130_fd_sc_hd__mux2_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12506_/X _12503_/X _12521_/D _12483_/Y _12504_/A vssd1 vssd1 vccd1 vccd1
+ _12534_/B sky130_fd_sc_hd__a221oi_1
XANTENNA__12993__A2 _12992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16290_ _19941_/Q _16290_/B vssd1 vssd1 vccd1 vccd1 _16291_/B sky130_fd_sc_hd__nand2_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15241_ _15241_/A vssd1 vssd1 vccd1 vccd1 _15241_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12453_ _18058_/A _12453_/B vssd1 vssd1 vccd1 vccd1 _12457_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13299__C _13299_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11402__C1 _10063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ _09998_/X _11393_/X _11402_/X _10065_/X _11403_/Y vssd1 vssd1 vccd1 vccd1
+ _12649_/A sky130_fd_sc_hd__o32a_4
X_15172_ _15172_/A vssd1 vssd1 vccd1 vccd1 _19117_/D sky130_fd_sc_hd__clkbuf_1
X_12384_ _19979_/Q _10240_/A _17464_/S vssd1 vssd1 vccd1 vccd1 _12385_/A sky130_fd_sc_hd__mux2_4
XANTENNA__15795__B _17220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14123_ _18687_/Q _13697_/X _14131_/S vssd1 vssd1 vccd1 vccd1 _14124_/A sky130_fd_sc_hd__mux2_1
X_11335_ _11183_/A _11332_/X _11334_/X vssd1 vssd1 vccd1 vccd1 _11335_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13596__A _15806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19980_ _19981_/CLK _19980_/D vssd1 vssd1 vccd1 vccd1 _19980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18931_ _19930_/CLK _18931_/D vssd1 vssd1 vccd1 vccd1 _18931_/Q sky130_fd_sc_hd__dfxtp_1
X_14054_ _14054_/A vssd1 vssd1 vccd1 vccd1 _18657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11266_ _11271_/A _11263_/X _11265_/X _18968_/Q vssd1 vssd1 vccd1 vccd1 _11266_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10732__B _10732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10217_ _10217_/A vssd1 vssd1 vccd1 vccd1 _10217_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13005_ _18930_/Q vssd1 vssd1 vccd1 vccd1 _13305_/A sky130_fd_sc_hd__inv_2
XFILLER_97_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18862_ _19299_/CLK _18862_/D vssd1 vssd1 vccd1 vccd1 _18862_/Q sky130_fd_sc_hd__dfxtp_1
X_11197_ _11274_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11197_/X sky130_fd_sc_hd__or2_1
XFILLER_95_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17813_ _17813_/A vssd1 vssd1 vccd1 vccd1 _17998_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10148_ _10148_/A vssd1 vssd1 vccd1 vccd1 _10148_/X sky130_fd_sc_hd__buf_2
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18793_ _19514_/CLK _18793_/D vssd1 vssd1 vccd1 vccd1 _18793_/Q sky130_fd_sc_hd__dfxtp_1
X_17744_ _17702_/A _17661_/X _17694_/X vssd1 vssd1 vccd1 vccd1 _17744_/Y sky130_fd_sc_hd__o21ai_2
X_14956_ _14956_/A vssd1 vssd1 vccd1 vccd1 _19018_/D sky130_fd_sc_hd__clkbuf_1
X_10079_ _10606_/A vssd1 vssd1 vccd1 vccd1 _10746_/A sky130_fd_sc_hd__buf_2
XFILLER_82_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12659__B _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ _13822_/X _18593_/Q _13911_/S vssd1 vssd1 vccd1 vccd1 _13908_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17675_ _17673_/X _17674_/X _17675_/S vssd1 vssd1 vccd1 vccd1 _17676_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14887_ _14634_/X _18988_/Q _14889_/S vssd1 vssd1 vccd1 vccd1 _14888_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19414_ _19510_/CLK _19414_/D vssd1 vssd1 vccd1 vccd1 _19414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16626_ _16627_/A _16627_/C _16625_/Y vssd1 vssd1 vccd1 vccd1 _19649_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17531__A _17542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13838_ _14663_/A vssd1 vssd1 vccd1 vccd1 _13838_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19345_ _19844_/CLK _19345_/D vssd1 vssd1 vccd1 vccd1 _19345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16557_ _17101_/A vssd1 vssd1 vccd1 vccd1 _16593_/A sky130_fd_sc_hd__clkbuf_2
X_13769_ _13767_/X _18544_/Q _13781_/S vssd1 vssd1 vccd1 vccd1 _13770_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16147__A _16204_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15508_ _15508_/A vssd1 vssd1 vccd1 vccd1 _19253_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19276_ _19406_/CLK _19276_/D vssd1 vssd1 vccd1 vccd1 _19276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17372__A1 _09188_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16488_ _19603_/Q _16487_/X _12468_/X _12471_/Y _16482_/X vssd1 vssd1 vccd1 vccd1
+ _19603_/D sky130_fd_sc_hd__o221a_1
XFILLER_50_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18227_ _19969_/Q _12119_/A _18231_/S vssd1 vssd1 vccd1 vccd1 _18228_/A sky130_fd_sc_hd__mux2_1
X_15439_ _14669_/X _19223_/Q _15439_/S vssd1 vssd1 vccd1 vccd1 _15440_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_61_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19480_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09984__A _10812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18158_ _18158_/A vssd1 vssd1 vccd1 vccd1 _19938_/D sky130_fd_sc_hd__clkbuf_1
X_17109_ _19798_/Q _17106_/B _17108_/Y vssd1 vssd1 vccd1 vccd1 _19798_/D sky130_fd_sc_hd__o21a_1
XFILLER_144_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18089_ _18087_/Y _18088_/X _18089_/S vssd1 vssd1 vccd1 vccd1 _18089_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_76_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19063_/CLK sky130_fd_sc_hd__clkbuf_16
X_09931_ _18787_/Q _19058_/Q _19282_/Q _19026_/Q _10270_/S _09929_/A vssd1 vssd1 vccd1
+ vccd1 _09931_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15925__S _15929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20051_ _20052_/CLK _20051_/D vssd1 vssd1 vccd1 vccd1 _20051_/Q sky130_fd_sc_hd__dfxtp_1
X_09862_ _18692_/Q _19187_/Q _10216_/S vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09793_ _09800_/A _09790_/X _09792_/X vssd1 vssd1 vccd1 vccd1 _09793_/Y sky130_fd_sc_hd__o21ai_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19971_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17363__A1 _09202_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17363__B2 _19888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19500_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09227_ _20048_/Q _20047_/Q _20046_/Q vssd1 vssd1 vccd1 vccd1 _09238_/A sky130_fd_sc_hd__or3_4
XFILLER_10_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09894__A _19918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13137__C1 _12805_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11120_ _18575_/Q _18836_/Q _18735_/Q _19070_/Q _10999_/A _11065_/A vssd1 vssd1 vccd1
+ vccd1 _11121_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11648__B _17331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11051_ _09746_/A _11040_/X _11049_/X _09753_/A _11050_/Y vssd1 vssd1 vccd1 vccd1
+ _12638_/B sky130_fd_sc_hd__o32a_4
XFILLER_89_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18434__A1_N _18349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10002_ _10792_/A vssd1 vssd1 vccd1 vccd1 _11395_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14810_ _14810_/A vssd1 vssd1 vccd1 vccd1 _14819_/S sky130_fd_sc_hd__buf_4
XANTENNA__11664__A _17338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15790_ _18459_/Q _12853_/X _15789_/X vssd1 vssd1 vccd1 vccd1 _17217_/A sky130_fd_sc_hd__a21oi_2
XFILLER_76_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18379__B1 _18374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14741_ _14741_/A vssd1 vssd1 vccd1 vccd1 _18922_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input14_A io_dbus_rdata[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10123__C1 _09738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11953_ _19822_/Q _13597_/A vssd1 vssd1 vccd1 vccd1 _11953_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17460_ _17832_/B _12385_/A _17460_/S vssd1 vssd1 vccd1 vccd1 _17460_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10904_ _19106_/Q _18872_/Q _19554_/Q _19202_/Q _11493_/S _09660_/A vssd1 vssd1 vccd1
+ vccd1 _10905_/B sky130_fd_sc_hd__mux4_1
XFILLER_33_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14672_ _14672_/A vssd1 vssd1 vccd1 vccd1 _14672_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ _17162_/A _13592_/A vssd1 vssd1 vccd1 vccd1 _11885_/B sky130_fd_sc_hd__or2_1
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16411_ _13321_/X _19563_/Q _16415_/S vssd1 vssd1 vccd1 vccd1 _16412_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13623_ _18509_/Q _13622_/X _13631_/S vssd1 vssd1 vccd1 vccd1 _13624_/A sky130_fd_sc_hd__mux2_1
X_10835_ _19365_/Q _18979_/Q _19429_/Q _18548_/Q _10735_/S _09970_/X vssd1 vssd1 vccd1
+ vccd1 _10836_/B sky130_fd_sc_hd__mux4_1
X_17391_ _17391_/A _17391_/B _17391_/C _17391_/D vssd1 vssd1 vccd1 vccd1 _17392_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13090__S _13090_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19130_ _19258_/CLK _19130_/D vssd1 vssd1 vccd1 vccd1 _19130_/Q sky130_fd_sc_hd__dfxtp_1
X_16342_ _16342_/A vssd1 vssd1 vccd1 vccd1 _19539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13554_ _13543_/Y _13553_/X _13554_/S vssd1 vssd1 vccd1 vccd1 _13554_/X sky130_fd_sc_hd__mux2_1
X_10766_ _11399_/A _10765_/X _10056_/X vssd1 vssd1 vccd1 vccd1 _10766_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10727__B _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12505_ _12520_/A vssd1 vssd1 vccd1 vccd1 _12505_/Y sky130_fd_sc_hd__inv_2
X_19061_ _19285_/CLK _19061_/D vssd1 vssd1 vccd1 vccd1 _19061_/Q sky130_fd_sc_hd__dfxtp_1
X_16273_ _19938_/Q _16273_/B vssd1 vssd1 vccd1 vccd1 _16274_/B sky130_fd_sc_hd__nand2_1
X_10697_ _10632_/A _10696_/X _10621_/X vssd1 vssd1 vccd1 vccd1 _10697_/X sky130_fd_sc_hd__o21a_1
XFILLER_139_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13485_ _13054_/A _13476_/Y _13484_/X _13324_/A vssd1 vssd1 vccd1 vccd1 _13485_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_145_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18012_ _18012_/A _18012_/B vssd1 vssd1 vccd1 vccd1 _18012_/Y sky130_fd_sc_hd__nor2_1
X_15224_ _15224_/A vssd1 vssd1 vccd1 vccd1 _19137_/D sky130_fd_sc_hd__clkbuf_1
X_12436_ _12459_/A _12436_/B vssd1 vssd1 vccd1 vccd1 _12436_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_154_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15155_ _19109_/Q vssd1 vssd1 vccd1 vccd1 _15156_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_126_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10743__A _11440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ _12538_/A _12362_/Y _11871_/X vssd1 vssd1 vccd1 vccd1 _12367_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12426__A2_N _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ _14106_/A vssd1 vssd1 vccd1 vccd1 _18679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output82_A _11740_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11318_ _19356_/Q _18970_/Q _19420_/Q _18539_/Q _11262_/X _11113_/A vssd1 vssd1 vccd1
+ vccd1 _11319_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09309__A _20042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15086_ _14608_/X _19076_/Q _15094_/S vssd1 vssd1 vccd1 vccd1 _15087_/A sky130_fd_sc_hd__mux2_1
X_12298_ _18321_/A _17334_/B _12190_/X vssd1 vssd1 vccd1 vccd1 _12298_/Y sky130_fd_sc_hd__a21oi_1
X_19963_ _19963_/CLK _19963_/D vssd1 vssd1 vccd1 vccd1 _19963_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09347__A1 _19890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18914_ _19439_/CLK _18914_/D vssd1 vssd1 vccd1 vccd1 _18914_/Q sky130_fd_sc_hd__dfxtp_1
X_14037_ _14059_/A vssd1 vssd1 vccd1 vccd1 _14046_/S sky130_fd_sc_hd__clkbuf_4
X_11249_ _19455_/Q _19293_/Q _18702_/Q _18472_/Q _11057_/S _11115_/A vssd1 vssd1 vccd1
+ vccd1 _11250_/B sky130_fd_sc_hd__mux4_1
XFILLER_79_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19894_ _19963_/CLK _19894_/D vssd1 vssd1 vccd1 vccd1 _19894_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18845_ _18845_/CLK _18845_/D vssd1 vssd1 vccd1 vccd1 _18845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15046__A _15046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18776_ _19559_/CLK _18776_/D vssd1 vssd1 vccd1 vccd1 _18776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15988_ _19419_/Q _15298_/X _15988_/S vssd1 vssd1 vccd1 vccd1 _15989_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15840__A1 _15839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17727_ _11625_/B _17729_/B _17865_/S _17726_/X vssd1 vssd1 vccd1 vccd1 _17727_/X
+ sky130_fd_sc_hd__o211a_1
X_14939_ _19011_/Q _14401_/X _14939_/S vssd1 vssd1 vccd1 vccd1 _14940_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17042__B1 _17021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17658_ _17477_/X _17497_/X _17686_/S vssd1 vssd1 vccd1 vccd1 _17658_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16609_ _16609_/A _16609_/B _19644_/Q vssd1 vssd1 vccd1 vccd1 _16611_/B sky130_fd_sc_hd__and3_1
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17589_ _17499_/X _17506_/X _17590_/S vssd1 vssd1 vccd1 vccd1 _17589_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14096__S _14098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19328_ _19881_/CLK _19328_/D vssd1 vssd1 vccd1 vccd1 _19328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19259_ _19389_/CLK _19259_/D vssd1 vssd1 vccd1 vccd1 _19259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10653__A _10700_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10815__S1 _10609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__A1 _10000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09219__A _19888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15655__S _15655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09914_ _19508_/Q _18920_/Q _18957_/Q _18531_/Q _10197_/S _09899_/X vssd1 vssd1 vccd1
+ vccd1 _09915_/B sky130_fd_sc_hd__mux4_1
XFILLER_99_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20034_ _20049_/CLK _20034_/D vssd1 vssd1 vccd1 vccd1 _20034_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input6_A io_dbus_rdata[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _10207_/A _09839_/X _09844_/X _09826_/X vssd1 vssd1 vccd1 vccd1 _09845_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11240__S1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _18663_/Q _19254_/Q _19416_/Q _18631_/Q _09542_/S _09526_/X vssd1 vssd1 vccd1
+ vccd1 _09777_/B sky130_fd_sc_hd__mux4_1
XFILLER_58_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13903__S _13911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ _11443_/A _10620_/B vssd1 vssd1 vccd1 vccd1 _10620_/X sky130_fd_sc_hd__or2_1
XANTENNA__12948__A2 _12946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10551_ _10544_/Y _10546_/Y _10548_/Y _10550_/Y _09718_/A vssd1 vssd1 vccd1 vccd1
+ _10551_/X sky130_fd_sc_hd__o221a_1
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10482_ _10478_/A _10479_/X _10481_/X _10307_/X vssd1 vssd1 vccd1 vccd1 _10482_/X
+ sky130_fd_sc_hd__o211a_1
X_13270_ _19907_/Q _13269_/X _13553_/S vssd1 vssd1 vccd1 vccd1 _13270_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12221_ _12935_/A _17334_/B _12190_/X vssd1 vssd1 vccd1 vccd1 _12221_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10806__S1 _10691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ _12152_/A _12178_/C vssd1 vssd1 vccd1 vccd1 _12153_/D sky130_fd_sc_hd__nand2_1
XFILLER_151_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11103_ _11153_/A _11103_/B vssd1 vssd1 vccd1 vccd1 _11103_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16960_ _19746_/Q _16971_/C _16833_/X vssd1 vssd1 vccd1 vccd1 _16961_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__17346__A _17346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12083_ _12083_/A _12083_/B vssd1 vssd1 vccd1 vccd1 _12084_/A sky130_fd_sc_hd__xnor2_4
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15911_ _15911_/A vssd1 vssd1 vccd1 vccd1 _19384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11034_ _18577_/Q _18838_/Q _18737_/Q _19072_/Q _10914_/X _11225_/A vssd1 vssd1 vccd1
+ vccd1 _11034_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16891_ _16923_/C _19727_/Q _19726_/Q _16891_/D vssd1 vssd1 vccd1 vccd1 _16900_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__17272__A0 _15724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18630_ _19511_/CLK _18630_/D vssd1 vssd1 vccd1 vccd1 _18630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15842_ _15842_/A vssd1 vssd1 vccd1 vccd1 _19354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15822__A1 _15818_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10990__S0 _10018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18561_ _19476_/CLK _18561_/D vssd1 vssd1 vccd1 vccd1 _18561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _15773_/A vssd1 vssd1 vccd1 vccd1 _19343_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output120_A _12632_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14909__S _14911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16396__S _16404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12985_ _19890_/Q vssd1 vssd1 vccd1 vccd1 _13173_/A sky130_fd_sc_hd__inv_2
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_4_clock_A _19998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13813__S _13813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17512_ _17493_/Y _17782_/A _17688_/A vssd1 vssd1 vccd1 vccd1 _17513_/A sky130_fd_sc_hd__mux2_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10647__B1 _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14724_ _18915_/Q _14433_/X _14724_/S vssd1 vssd1 vccd1 vccd1 _14725_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_157_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ _19569_/CLK _18492_/D vssd1 vssd1 vccd1 vccd1 _18492_/Q sky130_fd_sc_hd__dfxtp_1
X_11936_ _11936_/A _11936_/B vssd1 vssd1 vccd1 vccd1 _11938_/B sky130_fd_sc_hd__or2_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10742__S0 _10608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _17428_/X _17439_/X _17802_/B vssd1 vssd1 vccd1 vccd1 _17443_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14655_ _14655_/A vssd1 vssd1 vccd1 vccd1 _18888_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _11867_/A vssd1 vssd1 vccd1 vccd1 _12366_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12350__A2_N _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13606_ _13606_/A vssd1 vssd1 vccd1 vccd1 _18506_/D sky130_fd_sc_hd__clkbuf_1
X_10818_ _10613_/A _10815_/X _10817_/X _09976_/A vssd1 vssd1 vccd1 vccd1 _10818_/X
+ sky130_fd_sc_hd__o211a_1
X_17374_ _17374_/A vssd1 vssd1 vccd1 vccd1 _19891_/D sky130_fd_sc_hd__clkbuf_1
X_14586_ _14586_/A vssd1 vssd1 vccd1 vccd1 _14586_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11798_ _19580_/Q _12247_/A vssd1 vssd1 vccd1 vccd1 _11798_/X sky130_fd_sc_hd__and2_1
X_19113_ _19561_/CLK _19113_/D vssd1 vssd1 vccd1 vccd1 _19113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16325_ _19536_/Q _16324_/X _16325_/S vssd1 vssd1 vccd1 vccd1 _16326_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13537_ _13066_/X _13543_/B _13536_/X _13324_/A vssd1 vssd1 vccd1 vccd1 _13537_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10749_ _09614_/A _10739_/X _10748_/X _09621_/A _19904_/Q vssd1 vssd1 vccd1 vccd1
+ _11359_/A sky130_fd_sc_hd__a32o_2
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19044_ _19366_/CLK _19044_/D vssd1 vssd1 vccd1 vccd1 _19044_/Q sky130_fd_sc_hd__dfxtp_1
X_16256_ _16265_/C _16256_/B vssd1 vssd1 vccd1 vccd1 _16256_/Y sky130_fd_sc_hd__nand2_1
X_13468_ _19919_/Q _13467_/X _13468_/S vssd1 vssd1 vccd1 vccd1 _13468_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15207_ _19132_/Q _15206_/X _15213_/S vssd1 vssd1 vccd1 vccd1 _15208_/A sky130_fd_sc_hd__mux2_1
X_12419_ _19840_/Q _19839_/Q _12419_/C vssd1 vssd1 vccd1 vccd1 _12470_/C sky130_fd_sc_hd__and3_1
X_16187_ _19507_/Q _14650_/A _16189_/S vssd1 vssd1 vccd1 vccd1 _16188_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13399_ _19664_/Q vssd1 vssd1 vccd1 vccd1 _16670_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15138_ _15138_/A vssd1 vssd1 vccd1 vccd1 _19100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13784__A _13851_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15069_ _15069_/A vssd1 vssd1 vccd1 vccd1 _19068_/D sky130_fd_sc_hd__clkbuf_1
X_19946_ _19981_/CLK _19946_/D vssd1 vssd1 vccd1 vccd1 _19946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12875__A1 _16315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19877_ _19877_/CLK _19877_/D vssd1 vssd1 vccd1 vccd1 _19877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09630_ _10116_/A vssd1 vssd1 vccd1 vccd1 _10794_/A sky130_fd_sc_hd__buf_2
XFILLER_110_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18828_ _19666_/CLK _18828_/D vssd1 vssd1 vccd1 vccd1 _18828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15813__A1 _18463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09561_ _10426_/A vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12627__A1 _19848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18759_ _19511_/CLK _18759_/D vssd1 vssd1 vccd1 vccd1 _18759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14819__S _14819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09492_ _10243_/A vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09502__A _11428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10648__A _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_4_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12863__A _13343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12563__B1 _14477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18294__A2 _18291_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11461__S1 _10754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17166__A _17166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11118__A1 _11001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11669__A2 _11749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11213__S1 _10024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12866__B2 _19526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17254__A0 _13591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20017_ _20020_/CLK _20017_/D vssd1 vssd1 vccd1 vccd1 _20017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09828_ _10205_/A _09828_/B _09828_/C vssd1 vssd1 vccd1 vccd1 _09828_/X sky130_fd_sc_hd__or3_2
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15804__A1 _18462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09759_ _09720_/X _09742_/X _09750_/X _09757_/X _09758_/Y vssd1 vssd1 vccd1 vccd1
+ _12670_/B sky130_fd_sc_hd__o32ai_4
XANTENNA__14729__S _14735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10629__B1 _09979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12903_/A vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _12475_/A _18336_/A vssd1 vssd1 vccd1 vccd1 _11724_/B sky130_fd_sc_hd__or2_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11841__A2 _11950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14644_/A vssd1 vssd1 vccd1 vccd1 _14440_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11854_/B _11621_/Y _11628_/X _11651_/X vssd1 vssd1 vccd1 vccd1 _11652_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_70_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13043__B2 _19516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ _18809_/Q _19144_/Q _10811_/S vssd1 vssd1 vccd1 vccd1 _10604_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13869__A _13926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14371_ _15301_/A _15373_/C _15918_/B vssd1 vssd1 vccd1 vccd1 _14453_/A sky130_fd_sc_hd__nor3_4
XFILLER_70_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11583_ _11302_/A _12632_/B _11324_/X _12631_/B _11348_/Y vssd1 vssd1 vccd1 vccd1
+ _11586_/C sky130_fd_sc_hd__a221o_1
XFILLER_168_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16110_ _16110_/A vssd1 vssd1 vccd1 vccd1 _19472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13322_ _18486_/Q _13321_/X _13358_/S vssd1 vssd1 vccd1 vccd1 _13323_/A sky130_fd_sc_hd__mux2_1
X_10534_ _10534_/A _10534_/B vssd1 vssd1 vccd1 vccd1 _10534_/Y sky130_fd_sc_hd__nand2_1
X_17090_ _17090_/A vssd1 vssd1 vccd1 vccd1 _17095_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13588__B _13588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16041_ _13412_/X _19442_/Q _16045_/S vssd1 vssd1 vccd1 vccd1 _16042_/A sky130_fd_sc_hd__mux2_1
X_10465_ _18812_/Q _19147_/Q _10465_/S vssd1 vssd1 vccd1 vccd1 _10465_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13253_ _16265_/B _13254_/C _19938_/Q vssd1 vssd1 vccd1 vccd1 _13255_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12204_ _12204_/A vssd1 vssd1 vccd1 vccd1 _12204_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10396_ _10396_/A vssd1 vssd1 vccd1 vccd1 _10592_/A sky130_fd_sc_hd__clkbuf_2
X_13184_ _19333_/Q _12802_/A _12704_/A _19523_/Q _13183_/X vssd1 vssd1 vccd1 vccd1
+ _13184_/X sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_83_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19800_ _19803_/CLK _19800_/D vssd1 vssd1 vccd1 vccd1 _19800_/Q sky130_fd_sc_hd__dfxtp_1
X_12135_ _12188_/A _12649_/A _12134_/Y vssd1 vssd1 vccd1 vccd1 _12136_/A sky130_fd_sc_hd__a21o_1
XFILLER_97_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17992_ _17619_/X _17877_/X _17991_/X vssd1 vssd1 vccd1 vccd1 _17992_/X sky130_fd_sc_hd__a21o_1
XFILLER_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19731_ _19734_/CLK _19731_/D vssd1 vssd1 vccd1 vccd1 _19731_/Q sky130_fd_sc_hd__dfxtp_1
X_16943_ _17052_/A _16945_/B vssd1 vssd1 vccd1 vccd1 _16943_/X sky130_fd_sc_hd__or2_1
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12066_ _12086_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12066_/X sky130_fd_sc_hd__or2_1
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13109__A _15215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _18641_/Q _19232_/Q _19394_/Q _18609_/Q _10872_/S _09955_/A vssd1 vssd1 vccd1
+ vccd1 _11017_/X sky130_fd_sc_hd__mux4_1
X_16874_ _16874_/A _16874_/B _16883_/D vssd1 vssd1 vccd1 vccd1 _19722_/D sky130_fd_sc_hd__nor3_1
X_19662_ _19794_/CLK _19662_/D vssd1 vssd1 vccd1 vccd1 _19662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18613_ _19268_/CLK _18613_/D vssd1 vssd1 vccd1 vccd1 _18613_/Q sky130_fd_sc_hd__dfxtp_1
X_15825_ _15825_/A vssd1 vssd1 vccd1 vccd1 _19351_/D sky130_fd_sc_hd__clkbuf_1
X_19593_ _19608_/CLK _19593_/D vssd1 vssd1 vccd1 vccd1 _19593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _15756_/A vssd1 vssd1 vccd1 vccd1 _19339_/D sky130_fd_sc_hd__clkbuf_1
X_18544_ _19553_/CLK _18544_/D vssd1 vssd1 vccd1 vccd1 _18544_/Q sky130_fd_sc_hd__dfxtp_1
X_12968_ _18456_/Q _12966_/X _11415_/A _12962_/X vssd1 vssd1 vccd1 vccd1 _18456_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12667__B _12667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ _18907_/Q _14408_/X _14713_/S vssd1 vssd1 vccd1 vccd1 _14708_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11293__B1 _10988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _19822_/Q _11919_/B vssd1 vssd1 vccd1 vccd1 _11919_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18475_ _19895_/CLK _18475_/D vssd1 vssd1 vccd1 vccd1 _18475_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ _15737_/A _18442_/Q vssd1 vssd1 vccd1 vccd1 _15687_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12899_ _16923_/B _12719_/X _12723_/X _19697_/Q _12898_/X vssd1 vssd1 vccd1 vccd1
+ _12899_/X sky130_fd_sc_hd__a221o_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16220__A1 _16219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17426_ _17581_/S vssd1 vssd1 vccd1 vccd1 _17677_/S sky130_fd_sc_hd__clkbuf_2
X_14638_ _14637_/X _18883_/Q _14638_/S vssd1 vssd1 vccd1 vccd1 _14639_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14231__A0 _13758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17357_ _17376_/A vssd1 vssd1 vccd1 vccd1 _17373_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14569_ _14569_/A vssd1 vssd1 vccd1 vccd1 _18861_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14374__S _14386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11140__S0 _11035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16308_ _19944_/Q _16308_/B vssd1 vssd1 vccd1 vccd1 _16308_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17288_ _17288_/A vssd1 vssd1 vccd1 vccd1 _19867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19027_ _19027_/CLK _19027_/D vssd1 vssd1 vccd1 vccd1 _19027_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11299__A _19894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17338__C_N _18343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16239_ _19932_/Q _16239_/B vssd1 vssd1 vccd1 vccd1 _16240_/B sky130_fd_sc_hd__nand2_1
XFILLER_127_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18370__A input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11_0_clock_A clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19929_ _19930_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _19929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13019__A _13558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10954__S0 _09530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09613_ _09613_/A vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__buf_4
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14549__S _14557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__A _14476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _10082_/A vssd1 vssd1 vccd1 vccd1 _11190_/A sky130_fd_sc_hd__inv_2
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09475_ _09475_/A vssd1 vssd1 vccd1 vccd1 _09476_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13689__A _14634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14284__S _14290_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12593__A _12593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11131__S0 _11003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__S1 _09874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_105_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10250_ _10373_/A _10250_/B vssd1 vssd1 vccd1 vccd1 _10250_/X sky130_fd_sc_hd__or2_1
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17608__B _17610_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10181_ _10188_/A _10178_/X _10180_/X vssd1 vssd1 vccd1 vccd1 _10181_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_106_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13855__C _14844_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13940_ _13940_/A vssd1 vssd1 vccd1 vccd1 _18607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13871_ _13871_/A vssd1 vssd1 vccd1 vccd1 _18576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15610_ _15610_/A vssd1 vssd1 vccd1 vccd1 _19298_/D sky130_fd_sc_hd__clkbuf_1
X_12822_ _19810_/Q _12819_/X _14752_/B vssd1 vssd1 vccd1 vccd1 _12822_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16590_ _19637_/Q _19636_/Q _16590_/C vssd1 vssd1 vccd1 vccd1 _16597_/C sky130_fd_sc_hd__and3_1
XFILLER_46_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_3_0_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_15541_ _15587_/S vssd1 vssd1 vccd1 vccd1 _15550_/S sky130_fd_sc_hd__buf_2
XANTENNA__10078__B2 _10805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12753_ _13117_/A vssd1 vssd1 vccd1 vccd1 _12753_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11704_/A _11704_/B _12670_/A vssd1 vssd1 vccd1 vccd1 _11704_/X sky130_fd_sc_hd__or3_2
X_18260_ _19984_/Q _19605_/Q _18264_/S vssd1 vssd1 vccd1 vccd1 _18261_/A sky130_fd_sc_hd__mux2_1
X_15472_ _19237_/Q _15235_/X _15478_/S vssd1 vssd1 vccd1 vccd1 _15473_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12684_ _17322_/A _12684_/B _12684_/C vssd1 vssd1 vccd1 vccd1 _12791_/B sky130_fd_sc_hd__and3_1
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17950__A1 _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17211_ _17209_/Y _17197_/X _17210_/X _17201_/X vssd1 vssd1 vccd1 vccd1 _19837_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14423_/A vssd1 vssd1 vccd1 vccd1 _18810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18191_ _18191_/A vssd1 vssd1 vccd1 vccd1 _19953_/D sky130_fd_sc_hd__clkbuf_1
X_11635_ _12594_/B _11634_/X _11682_/A _11680_/C vssd1 vssd1 vccd1 vccd1 _17395_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14194__S _14196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17142_ _17185_/A vssd1 vssd1 vccd1 vccd1 _17142_/X sky130_fd_sc_hd__clkbuf_2
X_14354_ _14354_/A vssd1 vssd1 vccd1 vccd1 _14363_/S sky130_fd_sc_hd__clkbuf_4
X_11566_ _10674_/Y _11569_/B _10673_/A vssd1 vssd1 vccd1 vccd1 _11566_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13305_ _13305_/A _13436_/A vssd1 vssd1 vccd1 vccd1 _13354_/A sky130_fd_sc_hd__or2_1
XFILLER_156_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10517_ _10574_/A _10517_/B vssd1 vssd1 vccd1 vccd1 _10517_/X sky130_fd_sc_hd__or2_1
XFILLER_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17073_ _17073_/A vssd1 vssd1 vccd1 vccd1 _17108_/A sky130_fd_sc_hd__buf_2
X_14285_ _14285_/A vssd1 vssd1 vccd1 vccd1 _18757_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14922__S _14928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ _10665_/A _11494_/Y _11496_/Y _10116_/A vssd1 vssd1 vccd1 vccd1 _11497_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16024_ _16024_/A vssd1 vssd1 vccd1 vccd1 _19434_/D sky130_fd_sc_hd__clkbuf_1
X_13236_ _13233_/X _13235_/X _13299_/C vssd1 vssd1 vccd1 vccd1 _13236_/X sky130_fd_sc_hd__mux2_1
X_10448_ _10448_/A _10448_/B vssd1 vssd1 vccd1 vccd1 _10448_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17518__B _17542_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13167_ _13316_/A _15709_/B _15709_/C _13164_/X _13418_/A vssd1 vssd1 vccd1 vccd1
+ _13167_/X sky130_fd_sc_hd__o311a_1
X_10379_ _19375_/Q _18989_/Q _19439_/Q _18558_/Q _09505_/A _10312_/X vssd1 vssd1 vccd1
+ vccd1 _10380_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10553__A2 _10542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11750__A1 _11745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12118_ _12119_/A _12119_/B vssd1 vssd1 vccd1 vccd1 _12118_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13098_ _19743_/Q vssd1 vssd1 vccd1 vccd1 _16958_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17975_ _18078_/S _17976_/B _17974_/X _17723_/A vssd1 vssd1 vccd1 vccd1 _17978_/B
+ sky130_fd_sc_hd__o211a_1
X_19714_ _19718_/CLK _19714_/D vssd1 vssd1 vccd1 vccd1 _19714_/Q sky130_fd_sc_hd__dfxtp_1
X_16926_ _19738_/Q _19737_/Q _16926_/C vssd1 vssd1 vccd1 vccd1 _16959_/B sky130_fd_sc_hd__and3_1
X_12049_ _12049_/A _17462_/A vssd1 vssd1 vccd1 vccd1 _12050_/B sky130_fd_sc_hd__or2_1
XANTENNA__17769__A1 _17772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11502__A1 _10039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19645_ _19805_/CLK _19645_/D vssd1 vssd1 vccd1 vccd1 _19645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16857_ _19718_/Q _19717_/Q _19716_/Q _16857_/D vssd1 vssd1 vccd1 vccd1 _16870_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_1_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15808_ _15808_/A vssd1 vssd1 vccd1 vccd1 _15835_/S sky130_fd_sc_hd__clkbuf_2
X_16788_ _19700_/Q _16790_/C _16787_/Y vssd1 vssd1 vccd1 vccd1 _19700_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19576_ _19576_/CLK _19576_/D vssd1 vssd1 vccd1 vccd1 _19576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18527_ _19503_/CLK _18527_/D vssd1 vssd1 vccd1 vccd1 _18527_/Q sky130_fd_sc_hd__dfxtp_1
X_15739_ hold15/X _15738_/X _15757_/S vssd1 vssd1 vccd1 vccd1 _15739_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18365__A _18365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11361__S0 _10614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ _09426_/A _12601_/B vssd1 vssd1 vccd1 vccd1 _11663_/B sky130_fd_sc_hd__or2_1
X_18458_ _19985_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09191_ _20027_/Q _09191_/B _09271_/B vssd1 vssd1 vccd1 vccd1 _09269_/C sky130_fd_sc_hd__or3b_1
X_17409_ _17966_/B vssd1 vssd1 vccd1 vccd1 _17554_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_147_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18389_ _20032_/Q _18373_/X _18374_/X _18388_/Y vssd1 vssd1 vccd1 vccd1 _18390_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_14_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16613__A _16631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09926__S _09926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14133__A _14133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__buf_2
XFILLER_29_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14279__S _14279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12588__A _17240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09527_ _18965_/Q vssd1 vssd1 vccd1 vccd1 _11259_/S sky130_fd_sc_hd__clkbuf_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13911__S _13911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10155__S1 _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09465__A3 _17342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09458_ _09336_/Y _12678_/A _09412_/X _09403_/X vssd1 vssd1 vccd1 vccd1 _15662_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10836__A _10840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ _09389_/A _12688_/A _12688_/B vssd1 vssd1 vccd1 vccd1 _09391_/B sky130_fd_sc_hd__or3_2
XANTENNA__11104__S0 _11224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11420_ _11556_/A _11558_/A _11556_/C _10364_/A _11419_/Y vssd1 vssd1 vccd1 vccd1
+ _11552_/C sky130_fd_sc_hd__a311o_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10555__B _12653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11351_ _11581_/A _11349_/X _11582_/B vssd1 vssd1 vccd1 vccd1 _11351_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14742__S _14746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10302_ _10559_/S vssd1 vssd1 vccd1 vccd1 _10302_/X sky130_fd_sc_hd__clkbuf_4
X_14070_ _18665_/Q _13739_/X _14072_/S vssd1 vssd1 vccd1 vccd1 _14071_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11282_ _18796_/Q _19131_/Q _11327_/S vssd1 vssd1 vccd1 vccd1 _11283_/B sky130_fd_sc_hd__mux2_1
XANTENNA__17338__B _17338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17448__A0 _17937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13358__S _13358_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ _13021_/A vssd1 vssd1 vccd1 vccd1 _18469_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11667__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ _10233_/A _10233_/B vssd1 vssd1 vccd1 vccd1 _10233_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10164_ _10207_/A _10159_/X _10161_/X _10163_/X vssd1 vssd1 vccd1 vccd1 _10164_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input44_A io_ibus_inst[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10095_ _19511_/Q _18923_/Q _18960_/Q _18534_/Q _10081_/X _10691_/A vssd1 vssd1 vccd1
+ vccd1 _10096_/B sky130_fd_sc_hd__mux4_1
X_14972_ _19026_/Q _14449_/X _14972_/S vssd1 vssd1 vccd1 vccd1 _14973_/A sky130_fd_sc_hd__mux2_1
X_17760_ _17652_/X _17657_/X _17760_/S vssd1 vssd1 vccd1 vccd1 _17760_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13485__A1 _13054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__S0 _10914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13923_ _13923_/A vssd1 vssd1 vccd1 vccd1 _18600_/D sky130_fd_sc_hd__clkbuf_1
X_16711_ _16719_/D vssd1 vssd1 vccd1 vccd1 _16717_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17691_ _17681_/Y _17689_/X _17931_/S vssd1 vssd1 vccd1 vccd1 _17691_/X sky130_fd_sc_hd__mux2_1
X_19430_ _19430_/CLK _19430_/D vssd1 vssd1 vccd1 vccd1 _19430_/Q sky130_fd_sc_hd__dfxtp_1
X_16642_ _19654_/Q _16638_/B _16641_/Y vssd1 vssd1 vccd1 vccd1 _19654_/D sky130_fd_sc_hd__o21a_1
X_13854_ _16062_/A vssd1 vssd1 vccd1 vccd1 _16134_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__13237__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12805_ _12837_/A _12810_/B vssd1 vssd1 vccd1 vccd1 _12805_/Y sky130_fd_sc_hd__nor2_4
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16573_ _16573_/A _16573_/B _16574_/B vssd1 vssd1 vccd1 vccd1 _19631_/D sky130_fd_sc_hd__nor3_1
XFILLER_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19361_ _19553_/CLK _19361_/D vssd1 vssd1 vccd1 vccd1 _19361_/Q sky130_fd_sc_hd__dfxtp_1
X_13785_ _13783_/X _18549_/Q _13797_/S vssd1 vssd1 vccd1 vccd1 _13786_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10997_ _09746_/A _10983_/X _10995_/X _09753_/A _10996_/Y vssd1 vssd1 vccd1 vccd1
+ _12639_/B sky130_fd_sc_hd__o32a_4
XANTENNA__11343__S0 _11030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11799__A1 _11771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18312_ _20004_/Q _18310_/X _18311_/X _18303_/X vssd1 vssd1 vccd1 vccd1 _20004_/D
+ sky130_fd_sc_hd__o211a_1
X_15524_ _19260_/Q _15206_/X _15528_/S vssd1 vssd1 vccd1 vccd1 _15525_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15602__A _15659_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ _19292_/CLK _19292_/D vssd1 vssd1 vccd1 vccd1 _19292_/Q sky130_fd_sc_hd__dfxtp_1
X_12736_ _13578_/A vssd1 vssd1 vccd1 vccd1 _15702_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _18243_/A vssd1 vssd1 vccd1 vccd1 _19976_/D sky130_fd_sc_hd__clkbuf_1
X_15455_ _15455_/A vssd1 vssd1 vccd1 vccd1 _19229_/D sky130_fd_sc_hd__clkbuf_1
X_12667_ _12669_/A _12667_/B vssd1 vssd1 vccd1 vccd1 _12667_/Y sky130_fd_sc_hd__nor2_8
XFILLER_169_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10746__A _10746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09839__S1 _09809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14406_ _18805_/Q _14404_/X _14418_/S vssd1 vssd1 vccd1 vccd1 _14407_/A sky130_fd_sc_hd__mux2_1
X_11618_ _12378_/B vssd1 vssd1 vccd1 vccd1 _12475_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_18174_ _18174_/A vssd1 vssd1 vccd1 vccd1 _19945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15386_ _15443_/S vssd1 vssd1 vccd1 vccd1 _15395_/S sky130_fd_sc_hd__buf_2
XFILLER_156_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12598_ _12598_/A _12598_/B _12598_/C _12598_/D vssd1 vssd1 vccd1 vccd1 _12598_/X
+ sky130_fd_sc_hd__and4_1
X_17125_ _16708_/B _17123_/B _17101_/X vssd1 vssd1 vccd1 vccd1 _17125_/Y sky130_fd_sc_hd__a21oi_1
X_14337_ _18780_/Q _13685_/X _14341_/S vssd1 vssd1 vccd1 vccd1 _14338_/A sky130_fd_sc_hd__mux2_1
X_11549_ _11552_/A _11554_/A _11552_/C _10241_/A vssd1 vssd1 vccd1 vccd1 _11549_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17056_ _17056_/A vssd1 vssd1 vccd1 vccd1 _17062_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14268_ _13812_/X _18750_/Q _14268_/S vssd1 vssd1 vccd1 vccd1 _14269_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12592__B1_N _12319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16007_ _16007_/A vssd1 vssd1 vccd1 vccd1 _19426_/D sky130_fd_sc_hd__clkbuf_1
X_13219_ _15231_/A vssd1 vssd1 vccd1 vccd1 _13219_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11988__A2_N _12643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14199_ _13815_/X _18719_/Q _14207_/S vssd1 vssd1 vccd1 vccd1 _14200_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15483__S _15489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _17958_/A vssd1 vssd1 vccd1 vccd1 _18078_/S sky130_fd_sc_hd__buf_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16909_ _16925_/C _19733_/Q _16924_/B _16909_/D vssd1 vssd1 vccd1 vccd1 _16918_/D
+ sky130_fd_sc_hd__and4_1
X_17889_ _17729_/A _17695_/Y _17888_/Y vssd1 vssd1 vccd1 vccd1 _17983_/B sky130_fd_sc_hd__a21oi_2
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19628_ _19759_/CLK _19628_/D vssd1 vssd1 vccd1 vccd1 _19628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13228__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13016__B _14501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19559_ _19559_/CLK _19559_/D vssd1 vssd1 vccd1 vccd1 _19559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09312_ _20041_/Q _14501_/B vssd1 vssd1 vccd1 vccd1 _09320_/A sky130_fd_sc_hd__xor2_1
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11254__A3 _11253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09243_ _09243_/A vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09174_ _20021_/Q vssd1 vssd1 vccd1 vccd1 _09328_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14562__S _14568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16343__A _16347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11637__D _18288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10920_ _10920_/A vssd1 vssd1 vccd1 vccd1 _10920_/X sky130_fd_sc_hd__buf_2
XANTENNA__17902__A _17976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ _10665_/X _10848_/Y _10850_/Y _10794_/A vssd1 vssd1 vccd1 vccd1 _10851_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11325__S0 _11030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12978__B1 _10139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11950__A _19823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ _15837_/A vssd1 vssd1 vccd1 vccd1 _15737_/A sky130_fd_sc_hd__clkbuf_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10794_/A _10782_/B vssd1 vssd1 vccd1 vccd1 _10782_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17905__A1 _17705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12765__B _13316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12521_/A _12521_/B _12521_/C _12521_/D vssd1 vssd1 vccd1 vccd1 _12534_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09420__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15240_/A vssd1 vssd1 vccd1 vccd1 _19142_/D sky130_fd_sc_hd__clkbuf_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _18046_/A _12429_/B _17525_/A vssd1 vssd1 vccd1 vccd1 _12453_/B sky130_fd_sc_hd__o21ai_1
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12073__A2_N _12647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11403_ hold15/A vssd1 vssd1 vccd1 vccd1 _11403_/Y sky130_fd_sc_hd__clkinv_2
X_15171_ _19117_/Q vssd1 vssd1 vccd1 vccd1 _15172_/A sky130_fd_sc_hd__clkbuf_1
X_12383_ _12428_/A _12383_/B vssd1 vssd1 vccd1 vccd1 _12387_/A sky130_fd_sc_hd__nor2_1
XANTENNA__14472__S _14472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ _14133_/A vssd1 vssd1 vccd1 vccd1 _14131_/S sky130_fd_sc_hd__buf_2
X_11334_ _11291_/A _11333_/X _10980_/A vssd1 vssd1 vccd1 vccd1 _11334_/X sky130_fd_sc_hd__o21a_1
XANTENNA__16341__A0 _19539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14053_ _18657_/Q _13706_/X _14057_/S vssd1 vssd1 vccd1 vccd1 _14054_/A sky130_fd_sc_hd__mux2_1
X_18930_ _19895_/CLK _18930_/D vssd1 vssd1 vccd1 vccd1 _18930_/Q sky130_fd_sc_hd__dfxtp_1
X_11265_ _18967_/Q _11265_/B vssd1 vssd1 vccd1 vccd1 _11265_/X sky130_fd_sc_hd__or2_1
XFILLER_107_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13004_ _19925_/Q _13001_/X _13554_/S vssd1 vssd1 vccd1 vccd1 _13004_/X sky130_fd_sc_hd__mux2_1
X_10216_ _18689_/Q _19184_/Q _10216_/S vssd1 vssd1 vccd1 vccd1 _10217_/A sky130_fd_sc_hd__mux2_1
X_18861_ _19575_/CLK _18861_/D vssd1 vssd1 vccd1 vccd1 _18861_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output150_A _12269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11196_ _18573_/Q _18834_/Q _18733_/Q _19068_/Q _11259_/S _10880_/A vssd1 vssd1 vccd1
+ vccd1 _11197_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17812_ _17666_/S _17804_/X _17719_/X vssd1 vssd1 vccd1 vccd1 _17812_/X sky130_fd_sc_hd__o21ba_1
X_10147_ _10147_/A vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18792_ _19417_/CLK _18792_/D vssd1 vssd1 vccd1 vccd1 _18792_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14501__A _18293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11469__B1 _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14955_ _19018_/Q _14424_/X _14961_/S vssd1 vssd1 vccd1 vccd1 _14956_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17743_ _17738_/X _17742_/Y _17805_/S vssd1 vssd1 vccd1 vccd1 _17743_/X sky130_fd_sc_hd__mux2_2
X_10078_ _10070_/X _10072_/X _10075_/X _10805_/A _09979_/A vssd1 vssd1 vccd1 vccd1
+ _10090_/B sky130_fd_sc_hd__o221a_1
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_0_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13906_ _13906_/A vssd1 vssd1 vccd1 vccd1 _18592_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09314__B _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14886_ _14886_/A vssd1 vssd1 vccd1 vccd1 _18987_/D sky130_fd_sc_hd__clkbuf_1
X_17674_ _17590_/X _17579_/X _17674_/S vssd1 vssd1 vccd1 vccd1 _17674_/X sky130_fd_sc_hd__mux2_1
X_19413_ _19443_/CLK _19413_/D vssd1 vssd1 vccd1 vccd1 _19413_/Q sky130_fd_sc_hd__dfxtp_1
X_13837_ _13837_/A vssd1 vssd1 vccd1 vccd1 _18565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16625_ _16627_/A _16627_/C _16624_/X vssd1 vssd1 vccd1 vccd1 _16625_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_62_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16428__A _16428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__S0 _11003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16556_ _16573_/A _16556_/B _16558_/B vssd1 vssd1 vccd1 vccd1 _19625_/D sky130_fd_sc_hd__nor3_1
X_19344_ _19844_/CLK _19344_/D vssd1 vssd1 vccd1 vccd1 _19344_/Q sky130_fd_sc_hd__dfxtp_1
X_13768_ _13851_/S vssd1 vssd1 vccd1 vccd1 _13781_/S sky130_fd_sc_hd__buf_2
XFILLER_31_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15507_ _19253_/Q _15286_/X _15511_/S vssd1 vssd1 vccd1 vccd1 _15508_/A sky130_fd_sc_hd__mux2_1
X_12719_ _13341_/A vssd1 vssd1 vccd1 vccd1 _12719_/X sky130_fd_sc_hd__clkbuf_2
X_19275_ _19406_/CLK _19275_/D vssd1 vssd1 vccd1 vccd1 _19275_/Q sky130_fd_sc_hd__dfxtp_1
X_16487_ _16487_/A vssd1 vssd1 vccd1 vccd1 _16487_/X sky130_fd_sc_hd__clkbuf_2
X_13699_ _18527_/Q _13697_/X _13715_/S vssd1 vssd1 vccd1 vccd1 _13700_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15438_ _15438_/A vssd1 vssd1 vccd1 vccd1 _19222_/D sky130_fd_sc_hd__clkbuf_1
X_18226_ _18226_/A vssd1 vssd1 vccd1 vccd1 _19968_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15478__S _15478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _19192_/Q _15295_/X _15371_/S vssd1 vssd1 vccd1 vccd1 _15370_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18157_ _19938_/Q _19970_/Q _18159_/S vssd1 vssd1 vccd1 vccd1 _18158_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11944__A1 _19323_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17108_ _17108_/A _17112_/C vssd1 vssd1 vccd1 vccd1 _17108_/Y sky130_fd_sc_hd__nor2_1
X_18088_ _18090_/A _18090_/B _18088_/S vssd1 vssd1 vccd1 vccd1 _18088_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13146__A0 _19900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09930_ _18595_/Q _18856_/Q _18755_/Q _19090_/Q _10218_/S _09929_/X vssd1 vssd1 vccd1
+ vccd1 _09930_/X sky130_fd_sc_hd__mux4_1
X_17039_ _17039_/A _17039_/B vssd1 vssd1 vccd1 vccd1 _19769_/D sky130_fd_sc_hd__nor2_1
XANTENNA__18085__A0 _19920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10055__S0 _10053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20050_ _20052_/CLK _20050_/D vssd1 vssd1 vccd1 vccd1 _20050_/Q sky130_fd_sc_hd__dfxtp_2
X_09861_ _09924_/S vssd1 vssd1 vccd1 vccd1 _10216_/S sky130_fd_sc_hd__buf_4
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09770__C1 _09580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16102__S _16106_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09792_ _10188_/A _09791_/X _09712_/A vssd1 vssd1 vccd1 vccd1 _09792_/X sky130_fd_sc_hd__o21a_1
XFILLER_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14411__A _14615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09505__A _09505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12121__A1 _11745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10132__B1 _09706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14557__S _14557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16338__A _19950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11770__A _16487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17363__A2 _18301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09226_ _20050_/Q _20049_/Q _20051_/Q vssd1 vssd1 vccd1 vccd1 _09248_/B sky130_fd_sc_hd__or3b_1
XANTENNA__13697__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09589__C1 _10205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17169__A _17242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14292__S _14294_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16323__B1 _12444_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11148__C1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11010__A _11202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11050_ _19899_/Q vssd1 vssd1 vccd1 vccd1 _11050_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10001_ _10116_/A vssd1 vssd1 vccd1 vccd1 _10792_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13636__S _13652_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14321__A _14367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11664__B _18328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15851__S _15857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18379__B2 _18378_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14740_ _18922_/Q _14456_/X _14746_/S vssd1 vssd1 vccd1 vccd1 _14741_/A sky130_fd_sc_hd__mux2_1
X_11952_ _12693_/A _11952_/B _11952_/C _11952_/D vssd1 vssd1 vccd1 vccd1 _13597_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _10903_/A vssd1 vssd1 vccd1 vccd1 _11493_/S sky130_fd_sc_hd__clkbuf_4
X_14671_ _14671_/A vssd1 vssd1 vccd1 vccd1 _18893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11883_ _17162_/A _13592_/A vssd1 vssd1 vccd1 vccd1 _11917_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12776__A _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16410_ _16410_/A vssd1 vssd1 vccd1 vccd1 _19562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13622_ _14583_/A vssd1 vssd1 vccd1 vccd1 _13622_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10834_ _10834_/A _10834_/B _10834_/C vssd1 vssd1 vccd1 vccd1 _10834_/X sky130_fd_sc_hd__or3_1
X_17390_ _11627_/C _12594_/C _11692_/C _11901_/A vssd1 vssd1 vccd1 vccd1 _17391_/D
+ sky130_fd_sc_hd__a211o_1
X_16341_ _19539_/Q _16340_/X _16365_/S vssd1 vssd1 vccd1 vccd1 _16342_/A sky130_fd_sc_hd__mux2_1
X_13553_ _19924_/Q _13600_/B _13553_/S vssd1 vssd1 vccd1 vccd1 _13553_/X sky130_fd_sc_hd__mux2_1
X_10765_ _19495_/Q _18907_/Q _18944_/Q _18518_/Q _11451_/S _10037_/X vssd1 vssd1 vccd1
+ vccd1 _10765_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10296__A _10296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14991__A _15059_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19060_ _19478_/CLK _19060_/D vssd1 vssd1 vccd1 vccd1 _19060_/Q sky130_fd_sc_hd__dfxtp_1
X_12504_ _12504_/A _12503_/X vssd1 vssd1 vccd1 vccd1 _12520_/B sky130_fd_sc_hd__or2b_1
XFILLER_41_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_190_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19857_/CLK sky130_fd_sc_hd__clkbuf_16
X_16272_ _19938_/Q _16273_/B vssd1 vssd1 vccd1 vccd1 _16282_/C sky130_fd_sc_hd__or2_2
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ _13534_/S _10134_/Y _13147_/S _13483_/Y vssd1 vssd1 vccd1 vccd1 _13484_/X
+ sky130_fd_sc_hd__o211a_1
X_10696_ _18647_/Q _19238_/Q _19400_/Q _18615_/Q _10625_/X _10691_/X vssd1 vssd1 vccd1
+ vccd1 _10696_/X sky130_fd_sc_hd__mux4_1
X_18011_ _18008_/Y _18010_/X _18110_/S vssd1 vssd1 vccd1 vccd1 _18011_/X sky130_fd_sc_hd__mux2_1
X_15223_ _19137_/Q _15222_/X _15229_/S vssd1 vssd1 vccd1 vccd1 _15224_/A sky130_fd_sc_hd__mux2_1
X_12435_ _12521_/A _12521_/B vssd1 vssd1 vccd1 vccd1 _12436_/B sky130_fd_sc_hd__nand2_2
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15154_ _15154_/A vssd1 vssd1 vccd1 vccd1 _19108_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_0_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12366_ _12366_/A _12366_/B _12393_/B vssd1 vssd1 vccd1 vccd1 _12366_/X sky130_fd_sc_hd__or3_1
XANTENNA__16314__B1 _12127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_153_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14105_ _18679_/Q _13664_/X _14109_/S vssd1 vssd1 vccd1 vccd1 _14106_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11317_ _11317_/A _11317_/B vssd1 vssd1 vccd1 vccd1 _11317_/Y sky130_fd_sc_hd__nor2_1
X_15085_ _15131_/S vssd1 vssd1 vccd1 vccd1 _15094_/S sky130_fd_sc_hd__buf_4
XANTENNA__09309__B _14148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19962_ _19963_/CLK _19962_/D vssd1 vssd1 vccd1 vccd1 _19962_/Q sky130_fd_sc_hd__dfxtp_2
X_12297_ _12339_/B _12115_/X _12292_/X _12296_/X vssd1 vssd1 vccd1 vccd1 _12297_/X
+ sky130_fd_sc_hd__o22a_4
XANTENNA_output75_A _12148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14036_ _14036_/A vssd1 vssd1 vccd1 vccd1 _18649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18913_ _19501_/CLK _18913_/D vssd1 vssd1 vccd1 vccd1 _18913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09347__A2 _13173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11248_ _11117_/X _11247_/X _10875_/A vssd1 vssd1 vccd1 vccd1 _11248_/X sky130_fd_sc_hd__o21a_1
X_19893_ _19997_/CLK _19893_/D vssd1 vssd1 vccd1 vccd1 _19893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18844_ _19302_/CLK _18844_/D vssd1 vssd1 vccd1 vccd1 _18844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ _11179_/A vssd1 vssd1 vccd1 vccd1 _11179_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09325__A _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18775_ _18777_/CLK _18775_/D vssd1 vssd1 vccd1 vccd1 _18775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15987_ _15987_/A vssd1 vssd1 vccd1 vccd1 _19418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17542__A _17542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17726_ _17849_/A _17888_/A vssd1 vssd1 vccd1 vccd1 _17726_/X sky130_fd_sc_hd__or2_1
X_14938_ _14938_/A vssd1 vssd1 vccd1 vccd1 _19010_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_143_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19734_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17657_ _17481_/X _17490_/X _17660_/S vssd1 vssd1 vccd1 vccd1 _17657_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14377__S _14386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16158__A _16204_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14869_ _14915_/S vssd1 vssd1 vccd1 vccd1 _14878_/S sky130_fd_sc_hd__buf_6
XANTENNA__12686__A _17245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15062__A _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16608_ _16609_/A _16609_/B _16607_/Y vssd1 vssd1 vccd1 vccd1 _19643_/D sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_78_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17588_ _17586_/X _17587_/Y _17601_/S vssd1 vssd1 vccd1 vccd1 _17628_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19327_ _19762_/CLK _19327_/D vssd1 vssd1 vccd1 vccd1 _19327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16539_ _16573_/A _16539_/B _16539_/C vssd1 vssd1 vccd1 vccd1 _19619_/D sky130_fd_sc_hd__nor3_1
XANTENNA__18373__A _18413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_158_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19877_/CLK sky130_fd_sc_hd__clkbuf_16
X_19258_ _19258_/CLK _19258_/D vssd1 vssd1 vccd1 vccd1 _19258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18209_ _19961_/Q _19582_/Q _18209_/S vssd1 vssd1 vccd1 vccd1 _18210_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19189_ _19510_/CLK _19189_/D vssd1 vssd1 vccd1 vccd1 _19189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11749__B _11749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16621__A _16631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ _10254_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09913_/X sky130_fd_sc_hd__or2_1
XANTENNA__12342__A1 _11745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20033_ _20049_/CLK _20033_/D vssd1 vssd1 vccd1 vccd1 _20033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09844_ _10147_/A _09844_/B vssd1 vssd1 vccd1 vccd1 _09844_/X sky130_fd_sc_hd__or2_1
XFILLER_112_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09235__A _09238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ _09777_/A _09774_/X _09479_/X vssd1 vssd1 vccd1 vccd1 _09775_/X sky130_fd_sc_hd__o21a_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09316__B_N _14074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11853__A0 _18333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15700__A _15700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11081__A1 _10875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ _10588_/A _10549_/X _10323_/A vssd1 vssd1 vccd1 vccd1 _10550_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ _09209_/A vssd1 vssd1 vccd1 vccd1 _09209_/Y sky130_fd_sc_hd__inv_6
XFILLER_139_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10481_ _10521_/A _10481_/B vssd1 vssd1 vccd1 vccd1 _10481_/X sky130_fd_sc_hd__or2_1
XFILLER_120_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13220__A _13558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ _12338_/A _12115_/X _12213_/X _12219_/Y vssd1 vssd1 vccd1 vccd1 _12220_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11659__B _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12151_ _12152_/A _12178_/C vssd1 vssd1 vccd1 vccd1 _12153_/C sky130_fd_sc_hd__or2_1
XFILLER_163_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14750__S _14750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11102_ _19457_/Q _19295_/Q _18704_/Q _18474_/Q _11035_/X _11168_/A vssd1 vssd1 vccd1
+ vccd1 _11103_/B sky130_fd_sc_hd__mux4_1
XFILLER_150_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17346__B _17346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13125__A3 _15693_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ _12055_/A _12055_/B _12050_/A vssd1 vssd1 vccd1 vccd1 _12083_/B sky130_fd_sc_hd__a21bo_1
X_15910_ _13506_/X _19384_/Q _15912_/S vssd1 vssd1 vccd1 vccd1 _15911_/A sky130_fd_sc_hd__mux2_1
X_11033_ _11032_/A _11027_/Y _11032_/Y _11221_/A vssd1 vssd1 vccd1 vccd1 _11033_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16890_ _16923_/C _16896_/D vssd1 vssd1 vccd1 vccd1 _16892_/B sky130_fd_sc_hd__nor2_1
XFILLER_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15841_ _15840_/X _19354_/Q _15844_/S vssd1 vssd1 vccd1 vccd1 _15842_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15581__S _15583_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19512_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15822__A2 _18464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10990__S1 _11225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18560_ _19570_/CLK _18560_/D vssd1 vssd1 vccd1 vccd1 _18560_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _15771_/X _19343_/Q _15772_/S vssd1 vssd1 vccd1 vccd1 _15773_/A sky130_fd_sc_hd__mux2_1
X_12984_ _18468_/Q _12980_/X _12593_/Y _12947_/A vssd1 vssd1 vccd1 vccd1 _18468_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17511_ _17799_/S _17502_/X _17510_/X vssd1 vssd1 vccd1 vccd1 _17782_/A sky130_fd_sc_hd__o21ai_2
X_14723_ _14723_/A vssd1 vssd1 vccd1 vccd1 _18914_/D sky130_fd_sc_hd__clkbuf_1
X_11935_ _11905_/A _17421_/A _11934_/X vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__o21a_1
XFILLER_91_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ _19476_/CLK _18491_/D vssd1 vssd1 vccd1 vccd1 _18491_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output113_A _12649_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__S1 _10609_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12937__C _12937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14654_ _14653_/X _18888_/Q _14654_/S vssd1 vssd1 vccd1 vccd1 _14655_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _17602_/S vssd1 vssd1 vccd1 vccd1 _17802_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _19582_/Q _12218_/A vssd1 vssd1 vccd1 vccd1 _11892_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_75_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19575_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13605_ _13604_/X _18506_/Q _13605_/S vssd1 vssd1 vccd1 vccd1 _13606_/A sky130_fd_sc_hd__mux2_1
X_10817_ _10817_/A _10817_/B vssd1 vssd1 vccd1 vccd1 _10817_/X sky130_fd_sc_hd__or2_1
X_14585_ _14585_/A vssd1 vssd1 vccd1 vccd1 _18866_/D sky130_fd_sc_hd__clkbuf_1
X_17373_ _17373_/A _17373_/B vssd1 vssd1 vccd1 vccd1 _17374_/A sky130_fd_sc_hd__and2_1
X_11797_ _11797_/A vssd1 vssd1 vccd1 vccd1 _12247_/A sky130_fd_sc_hd__clkbuf_2
X_19112_ _19302_/CLK _19112_/D vssd1 vssd1 vccd1 vccd1 _19112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16324_ _16324_/A _16324_/B vssd1 vssd1 vccd1 vccd1 _16324_/X sky130_fd_sc_hd__or2_1
X_13536_ _19955_/Q _13536_/B vssd1 vssd1 vccd1 vccd1 _13536_/X sky130_fd_sc_hd__or2_1
XFILLER_174_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10748_ _09476_/A _10741_/X _10743_/X _10747_/X _09603_/A vssd1 vssd1 vccd1 vccd1
+ _10748_/X sky130_fd_sc_hd__a311o_2
XFILLER_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16255_ _19935_/Q _16255_/B vssd1 vssd1 vccd1 vccd1 _16256_/B sky130_fd_sc_hd__nand2_1
X_19043_ _19204_/CLK _19043_/D vssd1 vssd1 vccd1 vccd1 _19043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13467_ _19668_/Q _12832_/X _12833_/X _19800_/Q _13466_/X vssd1 vssd1 vccd1 vccd1
+ _13467_/X sky130_fd_sc_hd__a221o_4
XANTENNA__10754__A _10754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10679_ _18679_/Q _19174_/Q _11429_/S vssd1 vssd1 vccd1 vccd1 _10679_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14226__A _14294_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _15206_/A vssd1 vssd1 vccd1 vccd1 _15206_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12418_ _19537_/Q _12206_/X _12262_/X _12417_/X _12212_/X vssd1 vssd1 vccd1 vccd1
+ _12418_/X sky130_fd_sc_hd__o221a_1
X_16186_ _16186_/A vssd1 vssd1 vccd1 vccd1 _19506_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11569__B _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13398_ _13418_/A _13398_/B _13417_/B vssd1 vssd1 vccd1 vccd1 _13398_/X sky130_fd_sc_hd__or3_1
XFILLER_126_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10032__C1 _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15137_ _19100_/Q vssd1 vssd1 vccd1 vccd1 _15138_/A sky130_fd_sc_hd__clkbuf_1
X_12349_ _20042_/Q _12378_/B vssd1 vssd1 vccd1 vccd1 _12349_/X sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_13_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19966_/CLK sky130_fd_sc_hd__clkbuf_16
X_15068_ _14583_/X _19068_/Q _15072_/S vssd1 vssd1 vccd1 vccd1 _15069_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19945_ _19981_/CLK _19945_/D vssd1 vssd1 vccd1 vccd1 _19945_/Q sky130_fd_sc_hd__dfxtp_1
X_14019_ _14019_/A vssd1 vssd1 vccd1 vccd1 _18641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19876_ _19876_/CLK _19876_/D vssd1 vssd1 vccd1 vccd1 _19876_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold15_A hold15/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18827_ _19671_/CLK _18827_/D vssd1 vssd1 vccd1 vccd1 _18827_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_28_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19049_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15274__A0 _19153_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ _10523_/A vssd1 vssd1 vccd1 vccd1 _10426_/A sky130_fd_sc_hd__clkbuf_2
X_18758_ _19317_/CLK _18758_/D vssd1 vssd1 vccd1 vccd1 _18758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12627__A2 _17240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18212__A0 _19962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17709_ _11816_/A _17554_/B _18019_/A vssd1 vssd1 vccd1 vccd1 _17709_/Y sky130_fd_sc_hd__o21ai_1
X_09491_ _10373_/A vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18689_ _19411_/CLK _18689_/D vssd1 vssd1 vccd1 vccd1 _18689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11063__A1 _11001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10664__A _11460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12563__A1 _19543_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14570__S _14572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10603__S _10811_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11669__A3 _12562_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09827_ _09833_/A _09823_/X _09825_/X _09826_/X vssd1 vssd1 vccd1 vccd1 _09828_/C
+ sky130_fd_sc_hd__o211a_1
X_20016_ _20020_/CLK _20016_/D vssd1 vssd1 vccd1 vccd1 _20016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13914__S _13922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17182__A _17197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15804__A2 _13449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09758_ _19924_/Q vssd1 vssd1 vccd1 vccd1 _09758_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_101_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18203__A0 _19958_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10629__A1 _10296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _19515_/Q _18927_/Q _18964_/Q _18538_/Q _09726_/S _09788_/A vssd1 vssd1 vccd1
+ vccd1 _09689_/X sky130_fd_sc_hd__mux4_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _20046_/Q vssd1 vssd1 vccd1 vccd1 _18336_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09590__S1 _09526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11673_/C _11651_/B _11651_/C _11651_/D vssd1 vssd1 vccd1 vccd1 _11651_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_30_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15430__A _15430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ _10813_/A vssd1 vssd1 vccd1 vccd1 _10604_/A sky130_fd_sc_hd__clkbuf_4
X_14370_ _16371_/B vssd1 vssd1 vccd1 vccd1 _15373_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_23_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11582_ _11582_/A _11582_/B _11582_/C _11582_/D vssd1 vssd1 vccd1 vccd1 _11582_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13321_ _15254_/A vssd1 vssd1 vccd1 vccd1 _13321_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10533_ _18811_/Q _19146_/Q _10533_/S vssd1 vssd1 vccd1 vccd1 _10534_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10574__A _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16040_ _16040_/A vssd1 vssd1 vccd1 vccd1 _19441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13252_ hold15/A _15736_/B _13468_/S vssd1 vssd1 vccd1 vccd1 _13252_/X sky130_fd_sc_hd__mux2_1
X_10464_ _10476_/A _10464_/B vssd1 vssd1 vccd1 vccd1 _10464_/X sky130_fd_sc_hd__or2_1
XFILLER_129_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12203_ _12203_/A _12203_/B vssd1 vssd1 vccd1 vccd1 _12204_/A sky130_fd_sc_hd__xnor2_1
XFILLER_142_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13183_ _19859_/Q _12842_/A _13343_/A _19826_/Q vssd1 vssd1 vccd1 vccd1 _13183_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10395_ _18782_/Q _19053_/Q _19277_/Q _19021_/Q _10268_/S _10335_/A vssd1 vssd1 vccd1
+ vccd1 _10395_/X sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_26_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12134_ _12600_/A _12189_/A _12190_/A vssd1 vssd1 vccd1 vccd1 _12134_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17991_ _17560_/A _17983_/Y _17990_/X _17966_/Y vssd1 vssd1 vccd1 vccd1 _17991_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13503__A0 _19921_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19730_ _19734_/CLK _19730_/D vssd1 vssd1 vccd1 vccd1 _19730_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_96_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16942_ _16958_/B _16965_/C _16964_/A vssd1 vssd1 vccd1 vccd1 _16945_/B sky130_fd_sc_hd__and3_1
X_12065_ _17180_/A _12092_/C _12064_/Y vssd1 vssd1 vccd1 vccd1 _12065_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17245__A1 _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11016_ _11016_/A _11016_/B vssd1 vssd1 vccd1 vccd1 _11016_/X sky130_fd_sc_hd__or2_1
X_19661_ _19792_/CLK _19661_/D vssd1 vssd1 vccd1 vccd1 _19661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16873_ _16921_/C _19721_/Q _19720_/Q _16873_/D vssd1 vssd1 vccd1 vccd1 _16883_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_38_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18612_ _19204_/CLK _18612_/D vssd1 vssd1 vccd1 vccd1 _18612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15824_ _15823_/X _19351_/Q _15835_/S vssd1 vssd1 vccd1 vccd1 _15825_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16200__S _16200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19592_ _19592_/CLK _19592_/D vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfxtp_2
XFILLER_161_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09603__A _09603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18543_ _19794_/CLK _18543_/D vssd1 vssd1 vccd1 vccd1 _18543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ _18455_/Q _12966_/X _10459_/A _12962_/X vssd1 vssd1 vccd1 vccd1 _18455_/D
+ sky130_fd_sc_hd__a22o_1
X_15755_ _15753_/X _19339_/Q _15772_/S vssd1 vssd1 vccd1 vccd1 _15756_/A sky130_fd_sc_hd__mux2_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _14706_/A vssd1 vssd1 vccd1 vccd1 _18906_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11293__A1 _11170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11918_ _11885_/B _11917_/Y _11958_/B vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__a21boi_1
X_18474_ _19551_/CLK _18474_/D vssd1 vssd1 vccd1 vccd1 _18474_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ _19633_/Q _12891_/X _12897_/X vssd1 vssd1 vccd1 vccd1 _12898_/X sky130_fd_sc_hd__o21a_1
X_15686_ _18442_/Q _15686_/B vssd1 vssd1 vccd1 vccd1 _15686_/X sky130_fd_sc_hd__or2_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _17420_/X _17422_/X _17582_/S vssd1 vssd1 vccd1 vccd1 _17425_/X sky130_fd_sc_hd__mux2_1
X_14637_ _14637_/A vssd1 vssd1 vccd1 vccd1 _14637_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11849_ _17467_/A _11849_/B _11849_/C _11849_/D vssd1 vssd1 vccd1 vccd1 _11990_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_33_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _13844_/X _18861_/Q _14568_/S vssd1 vssd1 vccd1 vccd1 _14569_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10479__S0 _10417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17356_ _17356_/A vssd1 vssd1 vccd1 vccd1 _19886_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12242__B1 _12026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11140__S1 _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16307_ _19944_/Q _16308_/B vssd1 vssd1 vccd1 vccd1 _16321_/D sky130_fd_sc_hd__or2_2
X_13519_ _19671_/Q _12832_/X _12833_/X _19803_/Q _13518_/X vssd1 vssd1 vccd1 vccd1
+ _13519_/X sky130_fd_sc_hd__a221o_4
X_17287_ _12772_/B _19867_/Q _17291_/S vssd1 vssd1 vccd1 vccd1 _17288_/A sky130_fd_sc_hd__mux2_1
X_14499_ _18333_/A _14485_/X _14486_/X _14498_/Y vssd1 vssd1 vccd1 vccd1 _18412_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_173_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19026_ _19058_/CLK _19026_/D vssd1 vssd1 vccd1 vccd1 _19026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16238_ _19932_/Q _16239_/B vssd1 vssd1 vccd1 vccd1 _16248_/C sky130_fd_sc_hd__or2_2
XFILLER_155_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14390__S _14402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16169_ _16191_/A vssd1 vssd1 vccd1 vccd1 _16178_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_114_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17484__A1 _17937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19928_ _19930_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _19928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19859_ _19859_/CLK _19859_/D vssd1 vssd1 vccd1 vccd1 _19859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18098__A _18118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09612_ _09612_/A vssd1 vssd1 vccd1 vccd1 _09613_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10954__S1 _11236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12858__B _16268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ _18966_/Q vssd1 vssd1 vccd1 vccd1 _10082_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11762__B _17429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11808__B1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11284__A1 _11179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ _09979_/A vssd1 vssd1 vccd1 vccd1 _09475_/A sky130_fd_sc_hd__buf_2
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13025__A2 _13546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11131__S1 _11059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10890__S0 _09967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13909__S _13911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10180_ _09860_/A _10179_/X _09891_/X vssd1 vssd1 vccd1 vccd1 _10180_/X sky130_fd_sc_hd__o21a_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11429__S _11429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12114__A _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13644__S _13652_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15789__A1 _18459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870_ _13767_/X _18576_/Q _13878_/S vssd1 vssd1 vccd1 vccd1 _13871_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12768__B _18454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ _12855_/B vssd1 vssd1 vccd1 vccd1 _14752_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11275__A1 _10941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ _13116_/A vssd1 vssd1 vccd1 vccd1 _12752_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15540_ _15540_/A vssd1 vssd1 vccd1 vccd1 _19267_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11703_ _11894_/A vssd1 vssd1 vccd1 vccd1 _11856_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__10483__C1 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15471_ _15471_/A vssd1 vssd1 vccd1 vccd1 _19236_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _17146_/A _13560_/B vssd1 vssd1 vccd1 vccd1 _12684_/C sky130_fd_sc_hd__and2b_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _18810_/Q _14420_/X _14434_/S vssd1 vssd1 vccd1 vccd1 _14423_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17210_ _17210_/A _17210_/B vssd1 vssd1 vccd1 vccd1 _17210_/X sky130_fd_sc_hd__or2_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12379__A2_N _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ _09425_/B _11634_/B vssd1 vssd1 vccd1 vccd1 _11634_/X sky130_fd_sc_hd__and2b_1
X_18190_ _19953_/Q _19985_/Q _18192_/S vssd1 vssd1 vccd1 vccd1 _18191_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14353_ _14353_/A vssd1 vssd1 vccd1 vccd1 _18787_/D sky130_fd_sc_hd__clkbuf_1
X_17141_ _17141_/A _17140_/X vssd1 vssd1 vccd1 vccd1 _17141_/X sky130_fd_sc_hd__or2b_1
X_11565_ _11565_/A _11568_/A _11565_/C vssd1 vssd1 vccd1 vccd1 _11565_/Y sky130_fd_sc_hd__nand3_1
XFILLER_155_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _13173_/A _13173_/B _09349_/A input7/X _13174_/B vssd1 vssd1 vccd1 vccd1
+ _13436_/A sky130_fd_sc_hd__a41o_1
X_10516_ _18587_/Q _18848_/Q _18747_/Q _19082_/Q _10509_/S _10461_/A vssd1 vssd1 vccd1
+ vccd1 _10517_/B sky130_fd_sc_hd__mux4_1
XFILLER_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17072_ _17089_/A _17072_/B _17072_/C vssd1 vssd1 vccd1 vccd1 _19785_/D sky130_fd_sc_hd__nor3_1
X_14284_ _13835_/X _18757_/Q _14290_/S vssd1 vssd1 vccd1 vccd1 _14285_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15713__A1 _19901_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11496_ _11496_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11496_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16023_ _13277_/X _19434_/Q _16023_/S vssd1 vssd1 vccd1 vccd1 _16024_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13235_ _16265_/B _13254_/C vssd1 vssd1 vccd1 vccd1 _13235_/X sky130_fd_sc_hd__xor2_1
X_10447_ _19374_/Q _18988_/Q _19438_/Q _18557_/Q _10337_/X _10326_/X vssd1 vssd1 vccd1
+ vccd1 _10448_/B sky130_fd_sc_hd__mux4_1
XFILLER_143_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14504__A _14572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10633__S0 _10678_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ _13255_/A vssd1 vssd1 vccd1 vccd1 _13418_/A sky130_fd_sc_hd__buf_2
X_10378_ _10378_/A _10378_/B vssd1 vssd1 vccd1 vccd1 _10378_/X sky130_fd_sc_hd__or2_1
XFILLER_124_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11750__A2 _11740_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12117_ _12538_/A _12117_/B vssd1 vssd1 vccd1 vccd1 _12117_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17974_ _18033_/A _17977_/B _17539_/A _17973_/Y vssd1 vssd1 vccd1 vccd1 _17974_/X
+ sky130_fd_sc_hd__a211o_1
X_13097_ _19615_/Q vssd1 vssd1 vccd1 vccd1 _16527_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19713_ _19718_/CLK _19713_/D vssd1 vssd1 vccd1 vccd1 _19713_/Q sky130_fd_sc_hd__dfxtp_1
X_16925_ _19736_/Q _16925_/B _16925_/C _16925_/D vssd1 vssd1 vccd1 vccd1 _16926_/C
+ sky130_fd_sc_hd__and4_2
X_12048_ _12049_/A _17462_/A vssd1 vssd1 vccd1 vccd1 _12050_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17534__B _17534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12959__A _17861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13554__S _13554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19644_ _19805_/CLK _19644_/D vssd1 vssd1 vccd1 vccd1 _19644_/Q sky130_fd_sc_hd__dfxtp_1
X_16856_ _16874_/A _16856_/B _16856_/C vssd1 vssd1 vccd1 vccd1 _19717_/D sky130_fd_sc_hd__nor3_1
XFILLER_92_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15807_ _19918_/Q _12127_/A _16340_/A vssd1 vssd1 vccd1 vccd1 _15807_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19575_ _19575_/CLK _19575_/D vssd1 vssd1 vccd1 vccd1 _19575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16787_ _19700_/Q _16790_/C _16768_/X vssd1 vssd1 vccd1 vccd1 _16787_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13999_ _13999_/A vssd1 vssd1 vccd1 vccd1 _18634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18526_ _19503_/CLK _18526_/D vssd1 vssd1 vccd1 vccd1 _18526_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ _13587_/X _15736_/X _15737_/Y _12770_/X _18450_/Q vssd1 vssd1 vccd1 vccd1
+ _15738_/X sky130_fd_sc_hd__a32o_4
XFILLER_61_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10474__C1 _10519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11361__S1 _11371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18457_ _19985_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15669_ _09345_/X _15668_/X _13583_/Y vssd1 vssd1 vccd1 vccd1 _15669_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17408_ _17596_/B vssd1 vssd1 vccd1 vccd1 _17966_/B sky130_fd_sc_hd__buf_2
X_09190_ _09196_/A vssd1 vssd1 vccd1 vccd1 _09275_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18388_ input36/X vssd1 vssd1 vccd1 vccd1 _18388_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17339_ _17339_/A _18324_/A _17339_/C _18328_/A vssd1 vssd1 vccd1 vccd1 _17339_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12518__A1 _12421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19009_ _19491_/CLK _19009_/D vssd1 vssd1 vccd1 vccd1 _19009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10529__B1 _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09508__A _09508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_57_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16968__B1 _16833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ _09526_/A vssd1 vssd1 vccd1 vccd1 _09526_/X sky130_fd_sc_hd__buf_2
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09457_ _16816_/C _17346_/A vssd1 vssd1 vccd1 vccd1 _14479_/C sky130_fd_sc_hd__nand2_2
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09388_ _20015_/Q vssd1 vssd1 vccd1 vccd1 _18338_/A sky130_fd_sc_hd__inv_2
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11104__S1 _10917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ _11135_/X _12636_/B _11254_/Y _12634_/B vssd1 vssd1 vccd1 vccd1 _11582_/B
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10863__S0 _10702_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _10476_/A vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11281_ _11281_/A vssd1 vssd1 vccd1 vccd1 _11281_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16015__S _16023_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17448__A1 _17949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13020_ _18469_/Q _13009_/X _13090_/S vssd1 vssd1 vccd1 vccd1 _13021_/A sky130_fd_sc_hd__mux2_1
X_10232_ _18657_/Q _19248_/Q _19410_/Q _18625_/Q _09872_/X _09874_/X vssd1 vssd1 vccd1
+ vccd1 _10233_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09418__A _18138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10163_ _09569_/A _10162_/X _09833_/A vssd1 vssd1 vccd1 vccd1 _10163_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17635__A _17675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input37_A io_ibus_inst[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ _11443_/A _10094_/B vssd1 vssd1 vccd1 vccd1 _10094_/X sky130_fd_sc_hd__or2_1
X_14971_ _14971_/A vssd1 vssd1 vccd1 vccd1 _19025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16710_ _19675_/Q _19674_/Q _19805_/Q _16710_/D vssd1 vssd1 vccd1 vccd1 _16719_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__10918__S1 _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13922_ _13844_/X _18600_/Q _13922_/S vssd1 vssd1 vccd1 vccd1 _13923_/A sky130_fd_sc_hd__mux2_1
X_17690_ _17690_/A vssd1 vssd1 vccd1 vccd1 _17931_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16641_ _16674_/A _16645_/C vssd1 vssd1 vccd1 vccd1 _16641_/Y sky130_fd_sc_hd__nor2_1
X_13853_ _14148_/A _14501_/B vssd1 vssd1 vccd1 vccd1 _16062_/A sky130_fd_sc_hd__or2_1
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ _12804_/A _12810_/B vssd1 vssd1 vccd1 vccd1 _12804_/Y sky130_fd_sc_hd__nor2_2
X_19360_ _19455_/CLK _19360_/D vssd1 vssd1 vccd1 vccd1 _19360_/Q sky130_fd_sc_hd__dfxtp_1
X_16572_ hold14/X _19630_/Q _16572_/C vssd1 vssd1 vccd1 vccd1 _16574_/B sky130_fd_sc_hd__and3_1
XANTENNA__12445__B1 _12444_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13784_ _13851_/S vssd1 vssd1 vccd1 vccd1 _13797_/S sky130_fd_sc_hd__clkbuf_8
X_10996_ _19900_/Q vssd1 vssd1 vccd1 vccd1 _10996_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11343__S1 _09658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18311_ _18311_/A _18311_/B vssd1 vssd1 vccd1 vccd1 _18311_/X sky130_fd_sc_hd__or2_1
XFILLER_163_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15523_ _15523_/A vssd1 vssd1 vccd1 vccd1 _19259_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16187__A1 _14650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19291_ _19727_/CLK _19291_/D vssd1 vssd1 vccd1 vccd1 _19291_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12735_ _13580_/A vssd1 vssd1 vccd1 vccd1 _12735_/X sky130_fd_sc_hd__buf_2
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _19976_/Q _12339_/C _18242_/S vssd1 vssd1 vccd1 vccd1 _18243_/A sky130_fd_sc_hd__mux2_1
X_12666_ _12669_/A _12666_/B vssd1 vssd1 vccd1 vccd1 _12666_/Y sky130_fd_sc_hd__nor2_8
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15454_ _19229_/Q _15209_/X _15456_/S vssd1 vssd1 vccd1 vccd1 _15455_/A sky130_fd_sc_hd__mux2_1
X_14405_ _14472_/S vssd1 vssd1 vccd1 vccd1 _14418_/S sky130_fd_sc_hd__buf_2
X_11617_ _12320_/B vssd1 vssd1 vccd1 vccd1 _12378_/B sky130_fd_sc_hd__buf_2
X_18173_ _16313_/A _19977_/Q _18181_/S vssd1 vssd1 vccd1 vccd1 _18174_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15385_ _15385_/A vssd1 vssd1 vccd1 vccd1 _19198_/D sky130_fd_sc_hd__clkbuf_1
X_12597_ _17325_/A _12595_/B _11729_/A _17378_/A vssd1 vssd1 vccd1 vccd1 _12598_/C
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14933__S _14939_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17124_ _19804_/Q _17122_/B _17123_/Y vssd1 vssd1 vccd1 vccd1 _19804_/D sky130_fd_sc_hd__o21a_1
X_14336_ _14336_/A vssd1 vssd1 vccd1 vccd1 _18779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11548_ _11548_/A _11550_/A _11548_/C vssd1 vssd1 vccd1 vccd1 _11548_/Y sky130_fd_sc_hd__nand3_1
XFILLER_129_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14267_ _14267_/A vssd1 vssd1 vccd1 vccd1 _18749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17055_ _17089_/A _17055_/B _17055_/C vssd1 vssd1 vccd1 vccd1 _19779_/D sky130_fd_sc_hd__nor3_1
X_11479_ _11473_/A _11476_/X _11478_/X _09976_/A vssd1 vssd1 vccd1 vccd1 _11479_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13218_ _11656_/X _13216_/X _13217_/X vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__o21a_4
X_16006_ _13128_/X _19426_/Q _16012_/S vssd1 vssd1 vccd1 vccd1 _16007_/A sky130_fd_sc_hd__mux2_1
X_14198_ _14209_/A vssd1 vssd1 vccd1 vccd1 _14207_/S sky130_fd_sc_hd__buf_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12920__A1 _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13149_ _15222_/A vssd1 vssd1 vccd1 vccd1 _13149_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _17971_/A _17957_/B vssd1 vssd1 vccd1 vccd1 _17957_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16908_ _16925_/C _16915_/D vssd1 vssd1 vccd1 vccd1 _16910_/B sky130_fd_sc_hd__nor2_1
XFILLER_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17888_ _17888_/A _17888_/B vssd1 vssd1 vccd1 vccd1 _17888_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19627_ _19759_/CLK _19627_/D vssd1 vssd1 vccd1 vccd1 _19627_/Q sky130_fd_sc_hd__dfxtp_2
X_16839_ _19713_/Q _19712_/Q vssd1 vssd1 vccd1 vccd1 _16848_/D sky130_fd_sc_hd__and2_1
XFILLER_66_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09998__A _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19558_ _19560_/CLK _19558_/D vssd1 vssd1 vccd1 vccd1 _19558_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_148_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09311_ _19996_/Q vssd1 vssd1 vccd1 vccd1 _14501_/B sky130_fd_sc_hd__buf_4
XFILLER_62_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18509_ _19486_/CLK _18509_/D vssd1 vssd1 vccd1 vccd1 _18509_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16178__A1 _14637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19489_ _19489_/CLK _19489_/D vssd1 vssd1 vccd1 vccd1 _19489_/Q sky130_fd_sc_hd__dfxtp_1
X_09242_ _17379_/B _11650_/A _17379_/C vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__or3_2
XFILLER_22_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09173_ _20022_/Q vssd1 vssd1 vccd1 vccd1 _09328_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__11098__S0 _11035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10845__S0 _10702_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15689__A0 _19898_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10672__A _10672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09238__A _09238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17850__A1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13922__S _13922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10850_ _11387_/A _10850_/B vssd1 vssd1 vccd1 vccd1 _10850_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12978__A1 _18463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__S1 _09658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09509_ _18966_/Q vssd1 vssd1 vccd1 vccd1 _10880_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11950__B _11950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781_ _19108_/Q _18874_/Q _19556_/Q _19204_/Q _10849_/S _11496_/A vssd1 vssd1 vccd1
+ vccd1 _10782_/B sky130_fd_sc_hd__mux4_2
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18436__D input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12520_/A _12520_/B vssd1 vssd1 vccd1 vccd1 _12521_/D sky130_fd_sc_hd__nor2_1
XFILLER_13_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12451_/A vssd1 vssd1 vccd1 vccd1 _18058_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15849__S _15857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17118__B1 _17101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11402_ _11395_/Y _11397_/Y _11399_/Y _11401_/Y _10063_/X vssd1 vssd1 vccd1 vccd1
+ _11402_/X sky130_fd_sc_hd__o221a_2
X_15170_ _15170_/A vssd1 vssd1 vccd1 vccd1 _19116_/D sky130_fd_sc_hd__clkbuf_1
X_12382_ _18023_/A _12382_/B vssd1 vssd1 vccd1 vccd1 _12383_/B sky130_fd_sc_hd__and2_1
XFILLER_138_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14121_ _14121_/A vssd1 vssd1 vccd1 vccd1 _18686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11333_ _18571_/Q _18832_/Q _18731_/Q _19066_/Q _11035_/A _10006_/A vssd1 vssd1 vccd1
+ vccd1 _11333_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13155__A1 _12837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ _14052_/A vssd1 vssd1 vccd1 vccd1 _18656_/D sky130_fd_sc_hd__clkbuf_1
X_11264_ _18572_/Q _18833_/Q _18732_/Q _19067_/Q _11002_/A _10880_/A vssd1 vssd1 vccd1
+ vccd1 _11265_/B sky130_fd_sc_hd__mux4_1
XFILLER_4_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13003_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13554_/S sky130_fd_sc_hd__buf_2
X_10215_ _09616_/X _10205_/X _10214_/X _09623_/X _19915_/Q vssd1 vssd1 vccd1 vccd1
+ _10240_/A sky130_fd_sc_hd__a32o_2
XFILLER_106_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18860_ _19574_/CLK _18860_/D vssd1 vssd1 vccd1 vccd1 _18860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11195_ _18765_/Q _19036_/Q _19260_/Q _19004_/Q _09981_/A _09511_/A vssd1 vssd1 vccd1
+ vccd1 _11195_/X sky130_fd_sc_hd__mux4_1
X_17811_ _17783_/X _17810_/X _17931_/S vssd1 vssd1 vccd1 vccd1 _17811_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10146_ _10146_/A _11548_/A vssd1 vssd1 vccd1 vccd1 _11540_/A sky130_fd_sc_hd__or2b_1
X_18791_ _19512_/CLK _18791_/D vssd1 vssd1 vccd1 vccd1 _18791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output143_A _16465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14501__B _14501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11469__A1 _09748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11013__S0 _10893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17742_ _17742_/A vssd1 vssd1 vccd1 vccd1 _17742_/Y sky130_fd_sc_hd__clkinv_2
X_14954_ _14954_/A vssd1 vssd1 vccd1 vccd1 _19017_/D sky130_fd_sc_hd__clkbuf_1
X_10077_ _10817_/A vssd1 vssd1 vccd1 vccd1 _10805_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13905_ _13819_/X _18592_/Q _13911_/S vssd1 vssd1 vccd1 vccd1 _13906_/A sky130_fd_sc_hd__mux2_1
X_17673_ _17580_/X _17583_/X _17674_/S vssd1 vssd1 vccd1 vccd1 _17673_/X sky130_fd_sc_hd__mux2_1
X_14885_ _14631_/X _18987_/Q _14889_/S vssd1 vssd1 vccd1 vccd1 _14886_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14928__S _14928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19412_ _19412_/CLK _19412_/D vssd1 vssd1 vccd1 vccd1 _19412_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15613__A _15659_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16624_ _16860_/A vssd1 vssd1 vccd1 vccd1 _16624_/X sky130_fd_sc_hd__buf_2
X_13836_ _13835_/X _18565_/Q _13845_/S vssd1 vssd1 vccd1 vccd1 _13837_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11316__S1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _19873_/CLK _19343_/D vssd1 vssd1 vccd1 vccd1 _19343_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11860__B _17418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16555_ _19625_/Q _19624_/Q _16555_/C vssd1 vssd1 vccd1 vccd1 _16558_/B sky130_fd_sc_hd__and3_1
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10757__A _10757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13767_ _14592_/A vssd1 vssd1 vccd1 vccd1 _13767_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10979_ _18770_/Q _19041_/Q _19265_/Q _19009_/Q _11224_/S _11330_/A vssd1 vssd1 vccd1
+ vccd1 _10979_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15506_ _15506_/A vssd1 vssd1 vccd1 vccd1 _19252_/D sky130_fd_sc_hd__clkbuf_1
X_19274_ _19405_/CLK _19274_/D vssd1 vssd1 vccd1 vccd1 _19274_/Q sky130_fd_sc_hd__dfxtp_1
X_12718_ _12989_/A vssd1 vssd1 vccd1 vccd1 _13341_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16486_ _19602_/Q _16449_/X _12447_/X _16480_/X vssd1 vssd1 vccd1 vccd1 _19602_/D
+ sky130_fd_sc_hd__o211a_1
X_13698_ _13719_/A vssd1 vssd1 vccd1 vccd1 _13715_/S sky130_fd_sc_hd__clkbuf_4
X_18225_ _19968_/Q _19589_/Q _18231_/S vssd1 vssd1 vccd1 vccd1 _18226_/A sky130_fd_sc_hd__mux2_1
X_15437_ _14666_/X _19222_/Q _15439_/S vssd1 vssd1 vccd1 vccd1 _15438_/A sky130_fd_sc_hd__mux2_1
X_12649_ _12649_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _12649_/Y sky130_fd_sc_hd__nor2_2
XFILLER_30_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16444__A _18341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18156_ _18156_/A vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__clkbuf_1
X_15368_ _15368_/A vssd1 vssd1 vccd1 vccd1 _19191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17107_ _17107_/A vssd1 vssd1 vccd1 vccd1 _17112_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11944__A2 _11665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14319_ _18772_/Q _13651_/X _14319_/S vssd1 vssd1 vccd1 vccd1 _14320_/A sky130_fd_sc_hd__mux2_1
X_18087_ _18090_/A _18090_/B vssd1 vssd1 vccd1 vccd1 _18087_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15299_ _19161_/Q _15298_/X _15299_/S vssd1 vssd1 vccd1 vccd1 _15300_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17038_ _19769_/Q hold20/A _17034_/C _16635_/A vssd1 vssd1 vccd1 vccd1 _17039_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_74_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09860_ _09860_/A _09860_/B vssd1 vssd1 vccd1 vccd1 _09860_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10055__S1 _10054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _18791_/Q _19062_/Q _19286_/Q _19030_/Q _09787_/S _09688_/A vssd1 vssd1 vccd1
+ vccd1 _09791_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18989_ _19311_/CLK _18989_/D vssd1 vssd1 vccd1 vccd1 _18989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15843__B1 _13604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12212__A _13591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10668__C1 _09717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16619__A _16629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09521__A _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09225_ _11627_/B _09467_/B _09243_/A vssd1 vssd1 vccd1 vccd1 _11704_/B sky130_fd_sc_hd__and3_2
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12882__A _18273_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11935__A2 _17421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14602__A _14602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10000_ _10655_/A vssd1 vssd1 vccd1 vccd1 _10000_/X sky130_fd_sc_hd__buf_2
XFILLER_104_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09989_ _09989_/A _09989_/B vssd1 vssd1 vccd1 vccd1 _09989_/X sky130_fd_sc_hd__or2_1
XANTENNA__15834__A0 _19922_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10123__A1 _09706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _11951_/A _11951_/B vssd1 vssd1 vccd1 vccd1 _11956_/A sky130_fd_sc_hd__or2_1
XANTENNA__14748__S _14750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13652__S _13652_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ _11147_/A vssd1 vssd1 vccd1 vccd1 _10903_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14670_ _14669_/X _18893_/Q _14670_/S vssd1 vssd1 vccd1 vccd1 _14671_/A sky130_fd_sc_hd__mux2_1
X_11882_ _11878_/X _11879_/Y _11881_/X vssd1 vssd1 vccd1 vccd1 _13592_/A sky130_fd_sc_hd__a21oi_1
XFILLER_33_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09431__A _20041_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10833_ _09989_/A _10830_/X _10832_/X _10621_/A vssd1 vssd1 vccd1 vccd1 _10834_/C
+ sky130_fd_sc_hd__o211a_1
X_13621_ _15206_/A vssd1 vssd1 vccd1 vccd1 _14583_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16340_ _16340_/A _16340_/B vssd1 vssd1 vccd1 vccd1 _16340_/X sky130_fd_sc_hd__or2_1
X_10764_ _10764_/A _10764_/B vssd1 vssd1 vccd1 vccd1 _10764_/Y sky130_fd_sc_hd__nor2_1
X_13552_ _16507_/B _12727_/X _12729_/X _16708_/B _13551_/X vssd1 vssd1 vccd1 vccd1
+ _13600_/B sky130_fd_sc_hd__a221o_2
XFILLER_160_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12503_ _12503_/A _18079_/B vssd1 vssd1 vccd1 vccd1 _12503_/X sky130_fd_sc_hd__or2_1
XANTENNA__15579__S _15583_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16271_ _16271_/A vssd1 vssd1 vccd1 vccd1 _19526_/D sky130_fd_sc_hd__clkbuf_1
X_13483_ _13483_/A _13483_/B vssd1 vssd1 vccd1 vccd1 _13483_/Y sky130_fd_sc_hd__nand2_1
X_10695_ _11438_/A _10695_/B vssd1 vssd1 vccd1 vccd1 _10695_/X sky130_fd_sc_hd__or2_1
XFILLER_157_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18010_ _18012_/A _18012_/B _18088_/S vssd1 vssd1 vccd1 vccd1 _18010_/X sky130_fd_sc_hd__mux2_1
X_12434_ _12390_/A _12391_/A _12390_/B _12411_/B _12388_/A vssd1 vssd1 vccd1 vccd1
+ _12521_/B sky130_fd_sc_hd__a311o_2
XFILLER_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15222_ _15222_/A vssd1 vssd1 vccd1 vccd1 _15222_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10809__S0 _10073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15153_ _19108_/Q vssd1 vssd1 vccd1 vccd1 _15154_/A sky130_fd_sc_hd__clkbuf_1
X_12365_ _19597_/Q _19598_/Q _19599_/Q _12365_/D vssd1 vssd1 vccd1 vccd1 _12393_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_154_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14104_ _14104_/A vssd1 vssd1 vccd1 vccd1 _18678_/D sky130_fd_sc_hd__clkbuf_1
X_11316_ _19452_/Q _19290_/Q _18699_/Q _18469_/Q _11003_/A _11065_/A vssd1 vssd1 vccd1
+ vccd1 _11317_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19961_ _19997_/CLK _19961_/D vssd1 vssd1 vccd1 vccd1 _19961_/Q sky130_fd_sc_hd__dfxtp_2
X_15084_ _15084_/A vssd1 vssd1 vccd1 vccd1 _19075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12296_ _12127_/X _12294_/X _12295_/Y _12131_/X vssd1 vssd1 vccd1 vccd1 _12296_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11925__A2_N _12638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14035_ _18649_/Q _13672_/X _14035_/S vssd1 vssd1 vccd1 vccd1 _14036_/A sky130_fd_sc_hd__mux2_1
X_18912_ _19500_/CLK _18912_/D vssd1 vssd1 vccd1 vccd1 _18912_/Q sky130_fd_sc_hd__dfxtp_1
X_11247_ _19487_/Q _18899_/Q _18936_/Q _18510_/Q _11057_/S _10943_/X vssd1 vssd1 vccd1
+ vccd1 _11247_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11234__S0 _11129_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19892_ _19892_/CLK _19892_/D vssd1 vssd1 vccd1 vccd1 _19892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18843_ _19301_/CLK _18843_/D vssd1 vssd1 vccd1 vccd1 _18843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11178_ _11178_/A _11178_/B vssd1 vssd1 vccd1 vccd1 _11178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10129_ _19479_/Q _19317_/Q _18726_/Q _18496_/Q _10702_/S _09662_/A vssd1 vssd1 vccd1
+ vccd1 _10130_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13128__A _15219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18774_ _19369_/CLK _18774_/D vssd1 vssd1 vccd1 vccd1 _18774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15986_ _19418_/Q _15295_/X _15988_/S vssd1 vssd1 vccd1 vccd1 _15987_/A sky130_fd_sc_hd__mux2_1
X_17725_ _17725_/A vssd1 vssd1 vccd1 vccd1 _17865_/S sky130_fd_sc_hd__clkbuf_2
X_14937_ _19010_/Q _14398_/X _14939_/S vssd1 vssd1 vccd1 vccd1 _14938_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14658__S _14670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17656_ _17651_/Y _17655_/Y _17845_/A vssd1 vssd1 vccd1 vccd1 _17656_/X sky130_fd_sc_hd__mux2_1
X_14868_ _14868_/A vssd1 vssd1 vccd1 vccd1 _18979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16607_ _16609_/A _16609_/B _16577_/X vssd1 vssd1 vccd1 vccd1 _16607_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13819_ _14644_/A vssd1 vssd1 vccd1 vccd1 _13819_/X sky130_fd_sc_hd__clkbuf_1
X_17587_ _17721_/A _17486_/S _17802_/C vssd1 vssd1 vccd1 vccd1 _17587_/Y sky130_fd_sc_hd__a21boi_1
X_14799_ _14810_/A vssd1 vssd1 vccd1 vccd1 _14808_/S sky130_fd_sc_hd__clkbuf_4
X_19326_ _19756_/CLK _19326_/D vssd1 vssd1 vccd1 vccd1 _19326_/Q sky130_fd_sc_hd__dfxtp_1
X_16538_ _19619_/Q _16538_/B _16538_/C vssd1 vssd1 vccd1 vccd1 _16539_/C sky130_fd_sc_hd__and3_1
XFILLER_149_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15489__S _15489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19257_ _19952_/CLK _19257_/D vssd1 vssd1 vccd1 vccd1 _19257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16469_ _12119_/A _16449_/X _12125_/Y _12132_/X _16468_/X vssd1 vssd1 vccd1 vccd1
+ _19590_/D sky130_fd_sc_hd__o221a_1
XANTENNA__14393__S _14402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18208_ _18208_/A vssd1 vssd1 vccd1 vccd1 _19960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19188_ _19510_/CLK _19188_/D vssd1 vssd1 vccd1 vccd1 _19188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18139_ _18183_/A vssd1 vssd1 vccd1 vccd1 _18148_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__16305__A1 _12127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12207__A _17338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13119__B2 _19823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09912_ _19380_/Q _18994_/Q _19444_/Q _18563_/Q _10197_/S _09899_/X vssd1 vssd1 vccd1
+ vccd1 _09913_/B sky130_fd_sc_hd__mux4_1
XANTENNA__15518__A _15574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16113__S _16117_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09516__A _09813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20032_ _20032_/CLK _20032_/D vssd1 vssd1 vccd1 vccd1 _20032_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12342__A2 _12336_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09843_ _18660_/Q _19251_/Q _19413_/Q _18628_/Q _09904_/S _10151_/A vssd1 vssd1 vccd1
+ vccd1 _09844_/B sky130_fd_sc_hd__mux4_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _19512_/Q _18924_/Q _18961_/Q _18535_/Q _09542_/S _09526_/X vssd1 vssd1 vccd1
+ vccd1 _09774_/X sky130_fd_sc_hd__mux4_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14568__S _14568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13472__S _13524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11853__A1 _18321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16241__A0 _17127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13055__B1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09208_ _12610_/A _12610_/B _11638_/A vssd1 vssd1 vccd1 vccd1 _09209_/A sky130_fd_sc_hd__or3_2
X_10480_ _19469_/Q _19307_/Q _18716_/Q _18486_/Q _10559_/S _10510_/A vssd1 vssd1 vccd1
+ vccd1 _10481_/B sky130_fd_sc_hd__mux4_1
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12150_ _12152_/A _12150_/B vssd1 vssd1 vccd1 vccd1 _12160_/A sky130_fd_sc_hd__or2_1
XFILLER_118_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11101_ _10976_/X _11100_/X _10988_/X vssd1 vssd1 vccd1 vccd1 _11101_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_162_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12081_ _12081_/A _12081_/B vssd1 vssd1 vccd1 vccd1 _12083_/A sky130_fd_sc_hd__nor2_2
XANTENNA__16023__S _16023_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14332__A _14354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _11032_/A _11032_/B vssd1 vssd1 vccd1 vccd1 _11032_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10071__S _10675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15840_ _19923_/Q _15839_/X _15840_/S vssd1 vssd1 vccd1 vccd1 _15840_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_clock _19998_/CLK vssd1 vssd1 vccd1 vccd1 _19997_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _19912_/Q _15770_/X _15800_/S vssd1 vssd1 vccd1 vccd1 _15771_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15822__A3 _15819_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12787__A _18455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ _18467_/Q _12980_/X _11520_/A _12947_/A vssd1 vssd1 vccd1 vccd1 _18467_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _17649_/A _17510_/B vssd1 vssd1 vccd1 vccd1 _17510_/X sky130_fd_sc_hd__or2_1
XFILLER_45_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _18914_/Q _14430_/X _14724_/S vssd1 vssd1 vccd1 vccd1 _14723_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18490_ _19570_/CLK _18490_/D vssd1 vssd1 vccd1 vccd1 _18490_/Q sky130_fd_sc_hd__dfxtp_1
X_11934_ _11860_/A _17418_/A _11905_/A _17421_/A vssd1 vssd1 vccd1 vccd1 _11934_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17441_ _17649_/A vssd1 vssd1 vccd1 vccd1 _17602_/S sky130_fd_sc_hd__clkbuf_2
X_14653_ _14653_/A vssd1 vssd1 vccd1 vccd1 _14653_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _12066_/B vssd1 vssd1 vccd1 vccd1 _12218_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output106_A _17379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13604_ _13604_/A _13604_/B vssd1 vssd1 vccd1 vccd1 _13604_/X sky130_fd_sc_hd__or2_1
XANTENNA__10100__A _10817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10816_ _18581_/Q _18842_/Q _18741_/Q _19076_/Q _11483_/S _10074_/A vssd1 vssd1 vccd1
+ vccd1 _10817_/B sky130_fd_sc_hd__mux4_1
X_17372_ _09188_/Y _12824_/A _17358_/X _19891_/Q vssd1 vssd1 vccd1 vccd1 _17373_/B
+ sky130_fd_sc_hd__a22o_1
X_14584_ _14583_/X _18866_/Q _14590_/S vssd1 vssd1 vccd1 vccd1 _14585_/A sky130_fd_sc_hd__mux2_1
X_11796_ _11779_/X _11780_/Y _11784_/X _11795_/X vssd1 vssd1 vccd1 vccd1 _11796_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_158_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19111_ _19559_/CLK _19111_/D vssd1 vssd1 vccd1 vccd1 _19111_/Q sky130_fd_sc_hd__dfxtp_1
X_16323_ _16332_/C _16322_/Y _12444_/X vssd1 vssd1 vccd1 vccd1 _16324_/B sky130_fd_sc_hd__a21oi_2
XFILLER_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13535_ _19955_/Q _13536_/B vssd1 vssd1 vccd1 vccd1 _13543_/B sky130_fd_sc_hd__nand2_1
X_10747_ _11362_/A _10744_/X _10746_/X _10621_/X vssd1 vssd1 vccd1 vccd1 _10747_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19042_ _19042_/CLK _19042_/D vssd1 vssd1 vccd1 vccd1 _19042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16254_ _19935_/Q _16255_/B vssd1 vssd1 vccd1 vccd1 _16265_/C sky130_fd_sc_hd__or2_1
X_10678_ _18807_/Q _19142_/Q _10678_/S vssd1 vssd1 vccd1 vccd1 _10678_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13466_ _19732_/Q _13202_/X _13203_/X _19700_/Q _13465_/X vssd1 vssd1 vccd1 vccd1
+ _13466_/X sky130_fd_sc_hd__a221o_1
X_15205_ _15205_/A vssd1 vssd1 vccd1 vccd1 _19131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12417_ _12414_/Y _12416_/X _12562_/S vssd1 vssd1 vccd1 vccd1 _12417_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10258__S1 _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16185_ _19506_/Q _14647_/A _16189_/S vssd1 vssd1 vccd1 vccd1 _16186_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11455__S0 _10053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13397_ _19946_/Q _19947_/Q _13397_/C vssd1 vssd1 vccd1 vccd1 _13417_/B sky130_fd_sc_hd__and3_1
XFILLER_154_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15136_ _15136_/A vssd1 vssd1 vccd1 vccd1 _19099_/D sky130_fd_sc_hd__clkbuf_1
X_12348_ _12340_/A _11771_/X _12347_/X vssd1 vssd1 vccd1 vccd1 _12348_/X sky130_fd_sc_hd__o21a_4
XFILLER_153_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11780__B1 _19819_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15067_ _15067_/A vssd1 vssd1 vccd1 vccd1 _19067_/D sky130_fd_sc_hd__clkbuf_1
X_19944_ _19981_/CLK _19944_/D vssd1 vssd1 vccd1 vccd1 _19944_/Q sky130_fd_sc_hd__dfxtp_1
X_12279_ _12279_/A _12279_/B vssd1 vssd1 vccd1 vccd1 _12283_/A sky130_fd_sc_hd__and2_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14018_ _18641_/Q _13639_/X _14024_/S vssd1 vssd1 vccd1 vccd1 _14019_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19875_ _19879_/CLK _19875_/D vssd1 vssd1 vccd1 vccd1 _19875_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12875__A3 _12874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18826_ _19952_/CLK _18826_/D vssd1 vssd1 vccd1 vccd1 _18826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10430__S1 _10312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18757_ _19092_/CLK _18757_/D vssd1 vssd1 vccd1 vccd1 _18757_/Q sky130_fd_sc_hd__dfxtp_1
X_15969_ _19410_/Q _15270_/X _15973_/S vssd1 vssd1 vccd1 vccd1 _15970_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16169__A _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17708_ _17560_/X _17691_/X _17707_/X _17598_/X vssd1 vssd1 vccd1 vccd1 _17708_/X
+ sky130_fd_sc_hd__o211a_1
X_09490_ _10428_/A vssd1 vssd1 vccd1 vccd1 _10373_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18688_ _19409_/CLK _18688_/D vssd1 vssd1 vccd1 vccd1 _18688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16223__A0 _19518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ _18118_/A _17803_/S _17958_/A _17638_/X vssd1 vssd1 vccd1 vccd1 _17639_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18384__A _18396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19309_ _19564_/CLK _19309_/D vssd1 vssd1 vccd1 vccd1 _19309_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14417__A _14621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13321__A _15254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15947__S _15951_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__S1 _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15248__A hold10/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20015_ _20020_/CLK _20015_/D vssd1 vssd1 vccd1 vccd1 _20015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09826_ _09826_/A vssd1 vssd1 vccd1 vccd1 _09826_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10421__S1 _10312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09757_ _09757_/A vssd1 vssd1 vccd1 vccd1 _09757_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09688_/A vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10185__S0 _09881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16807__A _17247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11650_/A _17379_/C _17336_/A _11650_/D vssd1 vssd1 vccd1 vccd1 _11651_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10601_ _11411_/A _12651_/A vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__or2_1
X_11581_ _11581_/A vssd1 vssd1 vccd1 vccd1 _11582_/C sky130_fd_sc_hd__clkinv_2
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10532_ _10589_/S vssd1 vssd1 vccd1 vccd1 _10533_/S sky130_fd_sc_hd__buf_2
XFILLER_7_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13320_ _13060_/X _13315_/Y _13317_/X _13319_/X vssd1 vssd1 vccd1 vccd1 _15254_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_128_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17190__A1 _15738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15857__S _15857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__S0 _10625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10463_ _19115_/Q _18881_/Q _19563_/Q _19211_/Q _10382_/X _10462_/X vssd1 vssd1 vccd1
+ vccd1 _10464_/B sky130_fd_sc_hd__mux4_1
XFILLER_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13251_ _16645_/A _13116_/X _13117_/X _17079_/A _13250_/X vssd1 vssd1 vccd1 vccd1
+ _15736_/B sky130_fd_sc_hd__a221o_2
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12202_ _12174_/A _12174_/B _12170_/A vssd1 vssd1 vccd1 vccd1 _12203_/B sky130_fd_sc_hd__a21bo_1
X_13182_ _13255_/A vssd1 vssd1 vccd1 vccd1 _13337_/A sky130_fd_sc_hd__clkbuf_2
X_10394_ _10393_/A _10391_/Y _10393_/Y _10436_/A vssd1 vssd1 vccd1 vccd1 _10394_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_input67_A io_irq_motor_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_142_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19389_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12133_ _12119_/A _12115_/X _12125_/Y _12132_/X vssd1 vssd1 vccd1 vccd1 _12133_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _18002_/A _17990_/B _17990_/C _17990_/D vssd1 vssd1 vccd1 vccd1 _17990_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13503__A1 _13502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16941_ _16958_/B vssd1 vssd1 vccd1 vccd1 _16941_/Y sky130_fd_sc_hd__inv_2
X_12064_ _17180_/A _12092_/C _11778_/A vssd1 vssd1 vccd1 vccd1 _12064_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__15592__S _15600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11015_ _19490_/Q _18902_/Q _18939_/Q _18513_/Q _10893_/X _09955_/A vssd1 vssd1 vccd1
+ vccd1 _11016_/B sky130_fd_sc_hd__mux4_1
X_19660_ _19792_/CLK _19660_/D vssd1 vssd1 vccd1 vccd1 _19660_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_157_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19682_/CLK sky130_fd_sc_hd__clkbuf_16
X_16872_ _16921_/C _16880_/D vssd1 vssd1 vccd1 vccd1 _16874_/B sky130_fd_sc_hd__nor2_1
X_18611_ _19493_/CLK _18611_/D vssd1 vssd1 vccd1 vccd1 _18611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15823_ _19920_/Q _15822_/X _15840_/S vssd1 vssd1 vccd1 vccd1 _15823_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19591_ _19594_/CLK _19591_/D vssd1 vssd1 vccd1 vccd1 _19591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18542_ _18973_/CLK _18542_/D vssd1 vssd1 vccd1 vccd1 _18542_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15808_/A vssd1 vssd1 vccd1 vccd1 _15772_/S sky130_fd_sc_hd__clkbuf_2
X_12966_ _17861_/A vssd1 vssd1 vccd1 vccd1 _12966_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _18906_/Q _14404_/X _14713_/S vssd1 vssd1 vccd1 vccd1 _14706_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _11917_/A _11917_/B vssd1 vssd1 vccd1 vccd1 _11917_/Y sky130_fd_sc_hd__nand2_1
X_18473_ _19794_/CLK _18473_/D vssd1 vssd1 vccd1 vccd1 _18473_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17820__B _17820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _15685_/A vssd1 vssd1 vccd1 vccd1 _19328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _19761_/Q _12892_/X _12895_/X _12896_/X vssd1 vssd1 vccd1 vccd1 _12897_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ _17508_/S vssd1 vssd1 vccd1 vccd1 _17582_/S sky130_fd_sc_hd__clkbuf_2
X_14636_ _14636_/A vssd1 vssd1 vccd1 vccd1 _18882_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11848_ _19581_/Q _12150_/B _11829_/X _11847_/X vssd1 vssd1 vccd1 vccd1 _16453_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17355_/A _17355_/B vssd1 vssd1 vccd1 vccd1 _17356_/A sky130_fd_sc_hd__and2_1
XANTENNA__12242__A1 _19530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14567_ _14567_/A vssd1 vssd1 vccd1 vccd1 _18860_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10479__S1 _09841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11779_ _19819_/Q _11773_/X _11957_/A _12492_/A vssd1 vssd1 vccd1 vccd1 _11779_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__14237__A _14294_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16306_ _19532_/Q _16300_/X _16304_/Y _16305_/Y vssd1 vssd1 vccd1 vccd1 _19532_/D
+ sky130_fd_sc_hd__o22a_1
X_13518_ _19735_/Q _13202_/X _13203_/X _19703_/Q _13517_/X vssd1 vssd1 vccd1 vccd1
+ _13518_/X sky130_fd_sc_hd__a221o_1
XFILLER_146_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17286_ _17286_/A vssd1 vssd1 vccd1 vccd1 _19866_/D sky130_fd_sc_hd__clkbuf_1
X_14498_ input50/X vssd1 vssd1 vccd1 vccd1 _14498_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17181__A1 _15724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19025_ _19507_/CLK _19025_/D vssd1 vssd1 vccd1 vccd1 _19025_/Q sky130_fd_sc_hd__dfxtp_1
X_16237_ _16237_/A vssd1 vssd1 vccd1 vccd1 _19520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13449_ _16680_/A _12832_/X _12833_/X _17112_/A _13448_/X vssd1 vssd1 vccd1 vccd1
+ _13449_/X sky130_fd_sc_hd__a221o_4
XFILLER_174_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12980__A _17861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16168_ _16168_/A vssd1 vssd1 vccd1 vccd1 _19498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15119_ _14656_/X _19091_/Q _15127_/S vssd1 vssd1 vccd1 vccd1 _15120_/A sky130_fd_sc_hd__mux2_1
X_16099_ _16099_/A vssd1 vssd1 vccd1 vccd1 _19467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19927_ _19930_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _19927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19858_ _19859_/CLK _19858_/D vssd1 vssd1 vccd1 vccd1 _19858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09611_ _09611_/A vssd1 vssd1 vccd1 vccd1 _09612_/A sky130_fd_sc_hd__buf_4
X_18809_ _19495_/CLK _18809_/D vssd1 vssd1 vccd1 vccd1 _18809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19789_ _19789_/CLK _19789_/D vssd1 vssd1 vccd1 vccd1 _19789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15007__S _15011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09542_ _18826_/Q _19161_/Q _09542_/S vssd1 vssd1 vccd1 vccd1 _09542_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11808__A1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11808__B2 _19896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10167__S0 _09508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09473_ _09473_/A vssd1 vssd1 vccd1 vccd1 _09979_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13430__A0 _19917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10675__A _10675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13051__A _13299_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14581__S _14590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_74_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19481_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13497__B1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18289__A _18289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09809_ _09809_/A _09809_/B vssd1 vssd1 vccd1 vccd1 _09809_/X sky130_fd_sc_hd__and2_1
XFILLER_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15789__A2 _13407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19495_/CLK sky130_fd_sc_hd__clkbuf_16
X_12820_ _17146_/A _12820_/B _16808_/D vssd1 vssd1 vccd1 vccd1 _12855_/B sky130_fd_sc_hd__or3b_2
XFILLER_75_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12130__A _17187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18188__A0 _16347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _16921_/B _12719_/X _12723_/X _19691_/Q vssd1 vssd1 vccd1 vccd1 _13316_/B
+ sky130_fd_sc_hd__a22o_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14756__S _14764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19594_/CLK sky130_fd_sc_hd__clkbuf_16
X_11702_ _11712_/C vssd1 vssd1 vccd1 vccd1 _12673_/A sky130_fd_sc_hd__clkbuf_2
X_15470_ _19236_/Q _15231_/X _15478_/S vssd1 vssd1 vccd1 vccd1 _15471_/A sky130_fd_sc_hd__mux2_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _13136_/D _12693_/C vssd1 vssd1 vccd1 vccd1 _13560_/B sky130_fd_sc_hd__and2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14421_ _14453_/A vssd1 vssd1 vccd1 vccd1 _14434_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _17394_/A _12568_/B vssd1 vssd1 vccd1 vccd1 _11636_/C sky130_fd_sc_hd__nand2_1
XFILLER_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17140_ _17149_/A _17322_/A _17140_/C vssd1 vssd1 vccd1 vccd1 _17140_/X sky130_fd_sc_hd__and3b_1
X_14352_ _18787_/Q _13714_/X _14352_/S vssd1 vssd1 vccd1 vccd1 _14353_/A sky130_fd_sc_hd__mux2_1
X_11564_ _11568_/A _11565_/C _11565_/A vssd1 vssd1 vccd1 vccd1 _11564_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_27_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19501_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15587__S _15587_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ _13353_/A vssd1 vssd1 vccd1 vccd1 _13303_/X sky130_fd_sc_hd__clkbuf_2
X_10515_ _18779_/Q _19050_/Q _19274_/Q _19018_/Q _10470_/X _10462_/A vssd1 vssd1 vccd1
+ vccd1 _10515_/X sky130_fd_sc_hd__mux4_1
X_17071_ _17070_/B _17070_/C _19785_/Q vssd1 vssd1 vccd1 vccd1 _17072_/C sky130_fd_sc_hd__a21oi_1
X_14283_ _14283_/A vssd1 vssd1 vccd1 vccd1 _18756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11495_ _18825_/Q _19160_/Q _11495_/S vssd1 vssd1 vccd1 vccd1 _11496_/B sky130_fd_sc_hd__mux2_1
XFILLER_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16022_ _16022_/A vssd1 vssd1 vccd1 vccd1 _19433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10446_ _10323_/X _10436_/Y _10441_/X _10445_/Y _09740_/A vssd1 vssd1 vccd1 vccd1
+ _10446_/X sky130_fd_sc_hd__o311a_1
X_13234_ _19937_/Q vssd1 vssd1 vccd1 vccd1 _16265_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_137_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11735__B1 _12097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10377_ _19503_/Q _18915_/Q _18952_/Q _18526_/Q _09505_/A _10312_/X vssd1 vssd1 vccd1
+ vccd1 _10378_/B sky130_fd_sc_hd__mux4_1
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13255_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__10633__S1 _09813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12116_ _12116_/A vssd1 vssd1 vccd1 vccd1 _12538_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17973_ _17985_/A _17973_/B vssd1 vssd1 vccd1 vccd1 _17973_/Y sky130_fd_sc_hd__nor2_1
X_13096_ _19679_/Q vssd1 vssd1 vccd1 vccd1 _16727_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17815__B _17820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18199__A _18255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16924_ _19733_/Q _16924_/B _16924_/C _16924_/D vssd1 vssd1 vccd1 vccd1 _16925_/D
+ sky130_fd_sc_hd__and4_1
X_19712_ _19718_/CLK _19712_/D vssd1 vssd1 vccd1 vccd1 _19712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12047_ _19967_/Q _10821_/B _12198_/S vssd1 vssd1 vccd1 vccd1 _17462_/A sky130_fd_sc_hd__mux2_2
XFILLER_111_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09614__A _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16855_ _16868_/C _16864_/A _16857_/D vssd1 vssd1 vccd1 vccd1 _16856_/C sky130_fd_sc_hd__and3_1
X_19643_ _19877_/CLK _19643_/D vssd1 vssd1 vccd1 vccd1 _19643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15806_ _15806_/A _17225_/A vssd1 vssd1 vccd1 vccd1 _16340_/A sky130_fd_sc_hd__nor2_1
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19574_ _19574_/CLK _19574_/D vssd1 vssd1 vccd1 vccd1 _19574_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09333__B _17346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16786_ _19699_/Q _16784_/B _16785_/Y vssd1 vssd1 vccd1 vccd1 _19699_/D sky130_fd_sc_hd__o21a_1
X_13998_ _18634_/Q _13743_/X _13998_/S vssd1 vssd1 vccd1 vccd1 _13999_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18525_ _19406_/CLK _18525_/D vssd1 vssd1 vccd1 vccd1 _18525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15737_ _15737_/A _18450_/Q vssd1 vssd1 vccd1 vccd1 _15737_/Y sky130_fd_sc_hd__nand2_1
X_12949_ _18443_/Q _12946_/X _11352_/A _12947_/X vssd1 vssd1 vccd1 vccd1 _18443_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17926__A0 _19907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18456_ _19985_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15668_ _16213_/A vssd1 vssd1 vccd1 vccd1 _15668_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17407_ _17668_/A _17721_/C vssd1 vssd1 vccd1 vccd1 _17596_/B sky130_fd_sc_hd__or2_1
X_14619_ _14618_/X _18877_/Q _14622_/S vssd1 vssd1 vccd1 vccd1 _14620_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18387_ _18396_/A _18387_/B vssd1 vssd1 vccd1 vccd1 _20031_/D sky130_fd_sc_hd__nor2_1
X_15599_ _15599_/A vssd1 vssd1 vccd1 vccd1 _19293_/D sky130_fd_sc_hd__clkbuf_1
X_17338_ _17338_/A _17338_/B _18343_/A vssd1 vssd1 vccd1 vccd1 _17339_/C sky130_fd_sc_hd__or3b_1
XFILLER_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17269_ _15718_/X _19859_/Q _17269_/S vssd1 vssd1 vccd1 vccd1 _17270_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19008_ _19042_/CLK _19008_/D vssd1 vssd1 vccd1 vccd1 _19008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10529__A1 _09615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10529__B2 _19909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_144_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_60_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14430__A _14634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16968__A1 _19748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15960__S _15962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ _09773_/A _09525_/B vssd1 vssd1 vccd1 vccd1 _09525_/X sky130_fd_sc_hd__or2_1
XFILLER_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16357__A _16361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_69_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ input70/X vssd1 vssd1 vccd1 vccd1 _12747_/A sky130_fd_sc_hd__inv_2
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09387_ _16809_/A _12700_/A _09392_/C vssd1 vssd1 vccd1 vccd1 _12914_/B sky130_fd_sc_hd__and3b_1
XFILLER_61_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10863__S1 _09662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14605__A _14605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10300_ _10569_/A vssd1 vssd1 vccd1 vccd1 _10476_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13167__C1 _13418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11280_ _18668_/Q _19163_/Q _11280_/S vssd1 vssd1 vccd1 vccd1 _11281_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10231_ _10233_/A _10230_/X _09696_/X vssd1 vssd1 vccd1 vccd1 _10231_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10162_ _18818_/Q _19153_/Q _10162_/S vssd1 vssd1 vccd1 vccd1 _10162_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10093_ _19383_/Q _18997_/Q _19447_/Q _18566_/Q _10081_/X _10813_/A vssd1 vssd1 vccd1
+ vccd1 _10094_/B sky130_fd_sc_hd__mux4_1
X_14970_ _19025_/Q _14446_/X _14972_/S vssd1 vssd1 vccd1 vccd1 _14971_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10379__S0 _09505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13921_ _13921_/A vssd1 vssd1 vccd1 vccd1 _18599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16640_ _16640_/A vssd1 vssd1 vccd1 vccd1 _16645_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13852_ _13852_/A vssd1 vssd1 vccd1 vccd1 _18570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ _13077_/B vssd1 vssd1 vccd1 vccd1 _13546_/B sky130_fd_sc_hd__buf_2
X_16571_ _19630_/Q _16572_/C hold14/A vssd1 vssd1 vccd1 vccd1 _16573_/B sky130_fd_sc_hd__a21oi_1
X_13783_ _14608_/A vssd1 vssd1 vccd1 vccd1 _13783_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12795__A _18413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09846__C1 _09605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10995_ _10985_/Y _10989_/Y _10991_/Y _10993_/Y _10994_/X vssd1 vssd1 vccd1 vccd1
+ _10995_/X sky130_fd_sc_hd__o221a_1
X_18310_ _18323_/A vssd1 vssd1 vccd1 vccd1 _18310_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15522_ _19259_/Q _15203_/X _15528_/S vssd1 vssd1 vccd1 vccd1 _15523_/A sky130_fd_sc_hd__mux2_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19290_ _19290_/CLK _19290_/D vssd1 vssd1 vccd1 vccd1 _19290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12734_ _15700_/A vssd1 vssd1 vccd1 vccd1 _13580_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _18241_/A vssd1 vssd1 vccd1 vccd1 _19975_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15453_/A vssd1 vssd1 vccd1 vccd1 _19228_/D sky130_fd_sc_hd__clkbuf_1
X_12665_ _12669_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _12665_/Y sky130_fd_sc_hd__nor2_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _14608_/A vssd1 vssd1 vccd1 vccd1 _14404_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11204__A _11204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11616_ _11616_/A vssd1 vssd1 vccd1 vccd1 _12320_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_18172_ _18183_/A vssd1 vssd1 vccd1 vccd1 _18181_/S sky130_fd_sc_hd__clkbuf_2
X_15384_ _14589_/X _19198_/Q _15384_/S vssd1 vssd1 vccd1 vccd1 _15385_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12596_ _12596_/A _12596_/B _12596_/C _12595_/X vssd1 vssd1 vccd1 vccd1 _12599_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_168_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17123_ _17123_/A _17123_/B vssd1 vssd1 vccd1 vccd1 _17123_/Y sky130_fd_sc_hd__nor2_1
X_14335_ _18779_/Q _13681_/X _14341_/S vssd1 vssd1 vccd1 vccd1 _14336_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _11550_/A _11548_/C _11548_/A vssd1 vssd1 vccd1 vccd1 _11547_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14515__A _14572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15110__S _15116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16895__B1 _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17054_ _17053_/B _17053_/C _19779_/Q vssd1 vssd1 vccd1 vccd1 _17055_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__09609__A _09617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output98_A _11907_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14266_ _13809_/X _18749_/Q _14268_/S vssd1 vssd1 vccd1 vccd1 _14267_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11478_ _11478_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11478_/X sky130_fd_sc_hd__or2_1
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16005_ _16005_/A vssd1 vssd1 vccd1 vccd1 _19425_/D sky130_fd_sc_hd__clkbuf_1
X_13217_ input2/X _13172_/X _13175_/X vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__a21o_1
X_10429_ _18653_/Q _19244_/Q _19406_/Q _18621_/Q _10465_/S _10291_/X vssd1 vssd1 vccd1
+ vccd1 _10429_/X sky130_fd_sc_hd__mux4_1
X_14197_ _14197_/A vssd1 vssd1 vccd1 vccd1 _18718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ input30/X _12988_/A _13147_/X _13036_/X vssd1 vssd1 vccd1 vccd1 _15222_/A
+ sky130_fd_sc_hd__a22o_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13079_ _19854_/Q _12842_/X _12863_/X _19821_/Q _13078_/X vssd1 vssd1 vccd1 vccd1
+ _13079_/X sky130_fd_sc_hd__a221o_1
X_17956_ _19909_/Q _17758_/X _17955_/X vssd1 vssd1 vccd1 vccd1 _19909_/D sky130_fd_sc_hd__o21a_1
XFILLER_97_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16907_ _16919_/A _16907_/B _16915_/D vssd1 vssd1 vccd1 vccd1 _19733_/D sky130_fd_sc_hd__nor3_1
X_17887_ _17712_/X _17715_/X _17887_/S vssd1 vssd1 vccd1 vccd1 _17888_/B sky130_fd_sc_hd__mux2_1
XFILLER_66_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19626_ _19759_/CLK _19626_/D vssd1 vssd1 vccd1 vccd1 _19626_/Q sky130_fd_sc_hd__dfxtp_1
X_16838_ _16838_/A _16838_/B vssd1 vssd1 vccd1 vccd1 _19712_/D sky130_fd_sc_hd__nor2_1
XFILLER_54_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19557_ _19557_/CLK _19557_/D vssd1 vssd1 vccd1 vccd1 _19557_/Q sky130_fd_sc_hd__dfxtp_1
X_16769_ _19694_/Q _16772_/C _16768_/X vssd1 vssd1 vccd1 vccd1 _16769_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14396__S _14402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09310_ _18331_/A _14074_/B _09309_/X vssd1 vssd1 vccd1 vccd1 _09751_/B sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_70_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18508_ _19258_/CLK _18508_/D vssd1 vssd1 vccd1 vccd1 _18508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17375__A1 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19488_ _19488_/CLK _19488_/D vssd1 vssd1 vccd1 vccd1 _19488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09241_ _12610_/B _09244_/A _09249_/A vssd1 vssd1 vccd1 vccd1 _17379_/C sky130_fd_sc_hd__nor3_1
X_18439_ _19930_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09172_ _20023_/Q vssd1 vssd1 vccd1 vccd1 _18276_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11098__S1 _11330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10845__S1 _09662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10953__A _11250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15689__A1 _15688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09519__A _09841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10672__B _12650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11270__S1 _11059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17850__A2 _17853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10781__S0 _10849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09508_ _09508_/A vssd1 vssd1 vccd1 vccd1 _09763_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10030_/A _10779_/X _10652_/A vssd1 vssd1 vccd1 vccd1 _10780_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__17366__A1 _09209_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17366__B2 _13173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10989__A1 _11216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _17339_/A _18324_/A _11723_/B _09453_/B vssd1 vssd1 vccd1 vccd1 _09439_/X
+ sky130_fd_sc_hd__or4_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _12473_/A _12663_/B _12474_/A _12449_/X vssd1 vssd1 vccd1 vccd1 _12451_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_166_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11401_ _11383_/A _11400_/X _10000_/X vssd1 vssd1 vccd1 vccd1 _11401_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16026__S _16034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12381_ _18023_/A _12382_/B vssd1 vssd1 vccd1 vccd1 _12428_/A sky130_fd_sc_hd__nor2_1
XFILLER_166_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14120_ _18686_/Q _13693_/X _14120_/S vssd1 vssd1 vccd1 vccd1 _14121_/A sky130_fd_sc_hd__mux2_1
X_11332_ _18763_/Q _19034_/Q _19258_/Q _19002_/Q _11026_/S _11179_/X vssd1 vssd1 vccd1
+ vccd1 _11332_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14051_ _18656_/Q _13702_/X _14057_/S vssd1 vssd1 vccd1 vccd1 _14052_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13155__A2 _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11263_ _18764_/Q _19035_/Q _19259_/Q _19003_/Q _11262_/X _11113_/A vssd1 vssd1 vccd1
+ vccd1 _11263_/X sky130_fd_sc_hd__mux4_2
XFILLER_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13002_ _18929_/Q vssd1 vssd1 vccd1 vccd1 _13165_/A sky130_fd_sc_hd__inv_2
X_10214_ _09479_/A _10207_/X _10209_/X _10213_/X _09605_/X vssd1 vssd1 vccd1 vccd1
+ _10214_/X sky130_fd_sc_hd__a311o_1
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11194_ _11190_/X _11192_/X _11193_/X _11319_/A _09470_/A vssd1 vssd1 vccd1 vccd1
+ _11199_/B sky130_fd_sc_hd__o221a_1
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10145_ _10145_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _11548_/A sky130_fd_sc_hd__and2_1
X_17810_ _17470_/X _17493_/A _17810_/S vssd1 vssd1 vccd1 vccd1 _17810_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18790_ _19285_/CLK _18790_/D vssd1 vssd1 vccd1 vccd1 _18790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17741_ _17740_/Y _17629_/X _17741_/S vssd1 vssd1 vccd1 vccd1 _17742_/A sky130_fd_sc_hd__mux2_2
X_14953_ _19017_/Q _14420_/X _14961_/S vssd1 vssd1 vccd1 vccd1 _14954_/A sky130_fd_sc_hd__mux2_1
X_10076_ _11014_/A vssd1 vssd1 vccd1 vccd1 _10817_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13863__A0 _13758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11013__S1 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13904_ _13904_/A vssd1 vssd1 vccd1 vccd1 _18591_/D sky130_fd_sc_hd__clkbuf_1
X_17672_ _17672_/A vssd1 vssd1 vccd1 vccd1 _19895_/D sky130_fd_sc_hd__clkbuf_1
X_14884_ _14884_/A vssd1 vssd1 vccd1 vccd1 _18986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19411_ _19411_/CLK _19411_/D vssd1 vssd1 vccd1 vccd1 _19411_/Q sky130_fd_sc_hd__dfxtp_1
X_16623_ _16820_/A vssd1 vssd1 vccd1 vccd1 _16860_/A sky130_fd_sc_hd__clkbuf_2
X_13835_ _14660_/A vssd1 vssd1 vccd1 vccd1 _13835_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12418__A1 _19537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15105__S _15105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16554_ _19624_/Q _16555_/C _19625_/Q vssd1 vssd1 vccd1 vccd1 _16556_/B sky130_fd_sc_hd__a21oi_1
X_19342_ _19859_/CLK _19342_/D vssd1 vssd1 vccd1 vccd1 _19342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13766_ _13766_/A vssd1 vssd1 vccd1 vccd1 _18543_/D sky130_fd_sc_hd__clkbuf_1
X_10978_ _10978_/A vssd1 vssd1 vccd1 vccd1 _11330_/A sky130_fd_sc_hd__buf_4
XFILLER_44_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10524__S0 _10559_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15505_ _19252_/Q _15283_/X _15511_/S vssd1 vssd1 vccd1 vccd1 _15506_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19273_ _19405_/CLK _19273_/D vssd1 vssd1 vccd1 vccd1 _19273_/Q sky130_fd_sc_hd__dfxtp_1
X_12717_ _19722_/Q vssd1 vssd1 vccd1 vccd1 _16921_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16485_ _12416_/A _16477_/X _12418_/X _12423_/Y _16482_/X vssd1 vssd1 vccd1 vccd1
+ _19601_/D sky130_fd_sc_hd__o221a_1
X_13697_ _14640_/A vssd1 vssd1 vccd1 vccd1 _13697_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18224_ _18224_/A vssd1 vssd1 vccd1 vccd1 _19967_/D sky130_fd_sc_hd__clkbuf_1
X_15436_ _15436_/A vssd1 vssd1 vccd1 vccd1 _19221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _12648_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _12648_/Y sky130_fd_sc_hd__nor2_4
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18155_ _16265_/B _19969_/Q _18159_/S vssd1 vssd1 vccd1 vccd1 _18156_/A sky130_fd_sc_hd__mux2_1
X_15367_ _19191_/Q _15292_/X _15367_/S vssd1 vssd1 vccd1 vccd1 _15368_/A sky130_fd_sc_hd__mux2_1
X_12579_ _12579_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _12579_/X sky130_fd_sc_hd__xor2_4
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17106_ _17122_/A _17106_/B _17106_/C vssd1 vssd1 vccd1 vccd1 _19797_/D sky130_fd_sc_hd__nor3_1
XANTENNA__09339__A _09339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14318_ _14318_/A vssd1 vssd1 vccd1 vccd1 _18771_/D sky130_fd_sc_hd__clkbuf_1
X_18086_ _18086_/A vssd1 vssd1 vccd1 vccd1 _19920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15298_ _15298_/A vssd1 vssd1 vccd1 vccd1 _15298_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17037_ hold20/X _17034_/C _19769_/Q vssd1 vssd1 vccd1 vccd1 _17039_/A sky130_fd_sc_hd__a21oi_1
X_14249_ _13783_/X _18741_/Q _14257_/S vssd1 vssd1 vccd1 vccd1 _14250_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13295__S _13358_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09790_ _18599_/Q _18860_/Q _18759_/Q _19094_/Q _09724_/S _09730_/X vssd1 vssd1 vccd1
+ vccd1 _09790_/X sky130_fd_sc_hd__mux4_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _19564_/CLK _18988_/D vssd1 vssd1 vccd1 vccd1 _18988_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15843__A1 _19924_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17939_ _17934_/X _17936_/Y _17938_/X vssd1 vssd1 vccd1 vccd1 _17939_/X sky130_fd_sc_hd__o21a_1
XANTENNA__18387__A _18396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10763__S0 _09647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19609_ _19988_/CLK _19609_/D vssd1 vssd1 vccd1 vccd1 _19609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10948__A _11319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10515__S0 _10470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14854__S _14856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09224_ _11634_/B _09264_/B vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__or2b_1
XFILLER_148_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09589__A1 _09479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13137__A2 _12677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11148__A1 _11083_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12345__B1 _12855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09988_ _19510_/Q _18922_/Q _18959_/Q _18533_/Q _09984_/X _09970_/X vssd1 vssd1 vccd1
+ vccd1 _09989_/B sky130_fd_sc_hd__mux4_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17913__B _17914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18297__A _18297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13933__S _13939_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ _19823_/Q _11950_/B vssd1 vssd1 vccd1 vccd1 _11951_/B sky130_fd_sc_hd__nor2_1
XFILLER_18_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10901_ _11035_/A vssd1 vssd1 vccd1 vccd1 _11147_/A sky130_fd_sc_hd__buf_4
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11881_ _19815_/Q _19811_/Q _19806_/Q _11881_/D vssd1 vssd1 vccd1 vccd1 _11881_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__10858__A _11383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13620_ _13620_/A vssd1 vssd1 vccd1 vccd1 _18508_/D sky130_fd_sc_hd__clkbuf_1
X_10832_ _11473_/A _10832_/B vssd1 vssd1 vccd1 vccd1 _10832_/X sky130_fd_sc_hd__or2_1
XFILLER_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13551_ _19737_/Q _12775_/X _12777_/X _19705_/Q _13550_/X vssd1 vssd1 vccd1 vccd1
+ _13551_/X sky130_fd_sc_hd__a221o_1
X_10763_ _19367_/Q _18981_/Q _19431_/Q _18550_/Q _09647_/A _10030_/A vssd1 vssd1 vccd1
+ vccd1 _10764_/B sky130_fd_sc_hd__mux4_2
XANTENNA__10069__S _10812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14764__S _14764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12502_ _12503_/A _18079_/B vssd1 vssd1 vccd1 vccd1 _12504_/A sky130_fd_sc_hd__and2_1
XFILLER_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16270_ _19526_/Q _16269_/X _16280_/S vssd1 vssd1 vccd1 vccd1 _16271_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13482_ _19669_/Q _13116_/X _13117_/X _19801_/Q _13481_/X vssd1 vssd1 vccd1 vccd1
+ _13483_/B sky130_fd_sc_hd__a221o_4
X_10694_ _19464_/Q _19302_/Q _18711_/Q _18481_/Q _10690_/X _11371_/A vssd1 vssd1 vccd1
+ vccd1 _10695_/B sky130_fd_sc_hd__mux4_1
XFILLER_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15221_ _15221_/A vssd1 vssd1 vccd1 vccd1 _19136_/D sky130_fd_sc_hd__clkbuf_1
X_12433_ _12460_/A _18046_/B vssd1 vssd1 vccd1 vccd1 _12459_/A sky130_fd_sc_hd__xor2_4
XFILLER_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10809__S1 _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15152_ _15152_/A vssd1 vssd1 vccd1 vccd1 _19107_/D sky130_fd_sc_hd__clkbuf_1
X_12364_ _12340_/A _12340_/B _19599_/Q vssd1 vssd1 vccd1 vccd1 _12366_/B sky130_fd_sc_hd__a21oi_1
XFILLER_153_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ _18678_/Q _13660_/X _14109_/S vssd1 vssd1 vccd1 vccd1 _14104_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11315_ _11315_/A _11315_/B vssd1 vssd1 vccd1 vccd1 _11315_/Y sky130_fd_sc_hd__nor2_1
XFILLER_154_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19960_ _19997_/CLK _19960_/D vssd1 vssd1 vccd1 vccd1 _19960_/Q sky130_fd_sc_hd__dfxtp_2
X_15083_ _14605_/X _19075_/Q _15083_/S vssd1 vssd1 vccd1 vccd1 _15084_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12295_ _17205_/A _12316_/C vssd1 vssd1 vccd1 vccd1 _12295_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18911_ _19500_/CLK _18911_/D vssd1 vssd1 vccd1 vccd1 _18911_/Q sky130_fd_sc_hd__dfxtp_1
X_14034_ _14034_/A vssd1 vssd1 vccd1 vccd1 _18648_/D sky130_fd_sc_hd__clkbuf_1
X_11246_ _11304_/A _11246_/B vssd1 vssd1 vccd1 vccd1 _11246_/X sky130_fd_sc_hd__or2_1
X_19891_ _19892_/CLK _19891_/D vssd1 vssd1 vccd1 vccd1 _19891_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11234__S1 _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18842_ _19268_/CLK _18842_/D vssd1 vssd1 vccd1 vccd1 _18842_/Q sky130_fd_sc_hd__dfxtp_1
X_11177_ _19358_/Q _18972_/Q _19422_/Q _18541_/Q _11147_/A _10007_/A vssd1 vssd1 vccd1
+ vccd1 _11178_/B sky130_fd_sc_hd__mux4_1
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10128_ _11384_/S vssd1 vssd1 vccd1 vccd1 _10702_/S sky130_fd_sc_hd__buf_4
XFILLER_94_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15985_ _15985_/A vssd1 vssd1 vccd1 vccd1 _19417_/D sky130_fd_sc_hd__clkbuf_1
X_18773_ _19559_/CLK _18773_/D vssd1 vssd1 vccd1 vccd1 _18773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14939__S _14939_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15624__A _15646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ _18661_/Q _19252_/Q _19414_/Q _18629_/Q _11451_/S _10037_/X vssd1 vssd1 vccd1
+ vccd1 _10060_/B sky130_fd_sc_hd__mux4_1
X_14936_ _14936_/A vssd1 vssd1 vccd1 vccd1 _19009_/D sky130_fd_sc_hd__clkbuf_1
X_17724_ _17805_/S _17729_/B vssd1 vssd1 vccd1 vccd1 _17724_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18000__A _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__A1 _10941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10745__S0 _10617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09622__A _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17655_ _17802_/B _17652_/X _17654_/X vssd1 vssd1 vccd1 vccd1 _17655_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_63_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14867_ _14605_/X _18979_/Q _14867_/S vssd1 vssd1 vccd1 vccd1 _14868_/A sky130_fd_sc_hd__mux2_1
X_13818_ _13818_/A vssd1 vssd1 vccd1 vccd1 _18559_/D sky130_fd_sc_hd__clkbuf_1
X_16606_ _16609_/A _17041_/B vssd1 vssd1 vccd1 vccd1 _19642_/D sky130_fd_sc_hd__nor2_1
XFILLER_63_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17586_ _17507_/X _17503_/X _17586_/S vssd1 vssd1 vccd1 vccd1 _17586_/X sky130_fd_sc_hd__mux2_1
X_14798_ _14798_/A vssd1 vssd1 vccd1 vccd1 _18952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16537_ _16538_/B _16538_/C _19619_/Q vssd1 vssd1 vccd1 vccd1 _16539_/B sky130_fd_sc_hd__a21oi_1
X_19325_ _19852_/CLK _19325_/D vssd1 vssd1 vccd1 vccd1 _19325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13749_ _18293_/A _15198_/B _14844_/D vssd1 vssd1 vccd1 vccd1 _15373_/B sky130_fd_sc_hd__or3_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16455__A _17123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19256_ _19418_/CLK _19256_/D vssd1 vssd1 vccd1 vccd1 _19256_/Q sky130_fd_sc_hd__dfxtp_1
X_16468_ _16939_/A vssd1 vssd1 vccd1 vccd1 _16468_/X sky130_fd_sc_hd__clkbuf_2
X_15419_ _15430_/A vssd1 vssd1 vccd1 vccd1 _15428_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__15761__A0 _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18207_ _19960_/Q _19581_/Q _18209_/S vssd1 vssd1 vccd1 vccd1 _18208_/A sky130_fd_sc_hd__mux2_1
X_19187_ _19287_/CLK _19187_/D vssd1 vssd1 vccd1 vccd1 _19187_/Q sky130_fd_sc_hd__dfxtp_1
X_16399_ _16399_/A vssd1 vssd1 vccd1 vccd1 _19557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18138_ _18138_/A vssd1 vssd1 vccd1 vccd1 _18183_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16305__A2 _15764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10586__C1 _09718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18069_ _17771_/X _18065_/Y _18068_/Y vssd1 vssd1 vccd1 vccd1 _18069_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10008__A _11225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09911_ _09820_/X _09906_/X _09908_/X _09910_/X _09588_/A vssd1 vssd1 vccd1 vccd1
+ _09911_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20031_ _20032_/CLK _20031_/D vssd1 vssd1 vccd1 vccd1 _20031_/Q sky130_fd_sc_hd__dfxtp_1
X_09842_ _09842_/A vssd1 vssd1 vccd1 vccd1 _10151_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10984__S0 _10018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09773_/X sky130_fd_sc_hd__or2_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13753__S _13765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_14_0_clock clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09532__A _09532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13054__A _13054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14584__S _14590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09207_ _09275_/D vssd1 vssd1 vccd1 vccd1 _11638_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11302__A _11302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12030__A2 _12024_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12117__B _12117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16812__B _16812_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11100_ _19489_/Q _18901_/Q _18938_/Q _18512_/Q _10017_/A _10007_/A vssd1 vssd1 vccd1
+ vccd1 _11100_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09707__A _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_192_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _12080_/A _12080_/B vssd1 vssd1 vccd1 vccd1 _12081_/B sky130_fd_sc_hd__and2_1
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11031_ _18801_/Q _19136_/Q _11083_/S vssd1 vssd1 vccd1 vccd1 _11032_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15807__A1 _19918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10975__S0 _10018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15770_ _13587_/X _15768_/X _15769_/Y _12770_/X _18456_/Q vssd1 vssd1 vccd1 vccd1
+ _15770_/X sky130_fd_sc_hd__a32o_2
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _18466_/Q _12980_/X _11470_/A _12976_/X vssd1 vssd1 vccd1 vccd1 _18466_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12787__B _12787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _14721_/A vssd1 vssd1 vccd1 vccd1 _18913_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input12_A io_dbus_rdata[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09442__A _20028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11933_ _11933_/A _11933_/B _11933_/C vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__and3_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17440_ _17739_/S vssd1 vssd1 vccd1 vccd1 _17649_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _14652_/A vssd1 vssd1 vccd1 vccd1 _18887_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _11864_/A vssd1 vssd1 vccd1 vccd1 _11864_/Y sky130_fd_sc_hd__inv_8
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _15760_/A _13603_/B vssd1 vssd1 vccd1 vccd1 _13604_/B sky130_fd_sc_hd__and2_2
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _18773_/Q _19044_/Q _19268_/Q _19012_/Q _10617_/X _10609_/A vssd1 vssd1 vccd1
+ vccd1 _10815_/X sky130_fd_sc_hd__mux4_1
X_17371_ _17371_/A vssd1 vssd1 vccd1 vccd1 _19890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14583_ _14583_/A vssd1 vssd1 vccd1 vccd1 _14583_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11795_ _11745_/X _11767_/Y _11794_/Y vssd1 vssd1 vccd1 vccd1 _11795_/X sky130_fd_sc_hd__a21o_1
XANTENNA__14499__A1_N _18333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__S0 _10968_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19110_ _19302_/CLK _19110_/D vssd1 vssd1 vccd1 vccd1 _19110_/Q sky130_fd_sc_hd__dfxtp_1
X_16322_ _16313_/A _16317_/A _16321_/D _19947_/Q vssd1 vssd1 vccd1 vccd1 _16322_/Y
+ sky130_fd_sc_hd__o31ai_1
X_13534_ _19923_/Q _13533_/X _13534_/S vssd1 vssd1 vccd1 vccd1 _13534_/X sky130_fd_sc_hd__mux2_1
X_10746_ _10746_/A _10746_/B vssd1 vssd1 vccd1 vccd1 _10746_/X sky130_fd_sc_hd__or2_1
XFILLER_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19041_ _19491_/CLK _19041_/D vssd1 vssd1 vccd1 vccd1 _19041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16253_ _16253_/A vssd1 vssd1 vccd1 vccd1 _19523_/D sky130_fd_sc_hd__clkbuf_1
X_13465_ _19636_/Q _12839_/X _13464_/X vssd1 vssd1 vccd1 vccd1 _13465_/X sky130_fd_sc_hd__o21a_1
XFILLER_145_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ _10732_/A _10677_/B vssd1 vssd1 vccd1 vccd1 _10677_/X sky130_fd_sc_hd__or2_1
XFILLER_139_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15204_ _19131_/Q _15203_/X _15213_/S vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__mux2_1
X_12416_ _12416_/A _12438_/C vssd1 vssd1 vccd1 vccd1 _12416_/X sky130_fd_sc_hd__xor2_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16184_ _16184_/A vssd1 vssd1 vccd1 vccd1 _19505_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11455__S1 _10054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13396_ _19946_/Q _13397_/C _19947_/Q vssd1 vssd1 vccd1 vccd1 _13398_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10032__A1 _10014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17496__A0 _12455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15135_ _19099_/Q vssd1 vssd1 vccd1 vccd1 _15136_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_5_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12347_ _12123_/X _12342_/X _12343_/X _12346_/X _12131_/X vssd1 vssd1 vccd1 vccd1
+ _12347_/X sky130_fd_sc_hd__a311o_1
XFILLER_99_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15066_ _14580_/X _19067_/Q _15072_/S vssd1 vssd1 vccd1 vccd1 _15067_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11866__B _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09617__A _09617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19943_ _19981_/CLK _19943_/D vssd1 vssd1 vccd1 vccd1 _19943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12278_ _12278_/A _17452_/A vssd1 vssd1 vccd1 vccd1 _12279_/B sky130_fd_sc_hd__or2_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14017_ _14017_/A vssd1 vssd1 vccd1 vccd1 _18640_/D sky130_fd_sc_hd__clkbuf_1
X_11229_ _11183_/A _11228_/X _10920_/A vssd1 vssd1 vccd1 vccd1 _11229_/X sky130_fd_sc_hd__o21a_1
XFILLER_136_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19874_ _19876_/CLK _19874_/D vssd1 vssd1 vccd1 vccd1 _19874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18825_ _19418_/CLK _18825_/D vssd1 vssd1 vccd1 vccd1 _18825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18756_ _19449_/CLK _18756_/D vssd1 vssd1 vccd1 vccd1 _18756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15968_ _15968_/A vssd1 vssd1 vccd1 vccd1 _19409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13285__B2 _19529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17707_ _17524_/X _17696_/Y _17706_/X _17667_/A vssd1 vssd1 vccd1 vccd1 _17707_/X
+ sky130_fd_sc_hd__a211o_1
X_14919_ _14987_/S vssd1 vssd1 vccd1 vccd1 _14928_/S sky130_fd_sc_hd__buf_2
X_15899_ _13423_/X _19379_/Q _15901_/S vssd1 vssd1 vccd1 vccd1 _15900_/A sky130_fd_sc_hd__mux2_1
X_18687_ _19409_/CLK _18687_/D vssd1 vssd1 vccd1 vccd1 _18687_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17420__A0 _17729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17638_ _17914_/A _17642_/B vssd1 vssd1 vccd1 vccd1 _17638_/X sky130_fd_sc_hd__or2_1
XFILLER_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11048__B1 _10920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17569_ _17453_/X _17446_/X _17582_/S vssd1 vssd1 vccd1 vccd1 _17569_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19308_ _19308_/CLK _19308_/D vssd1 vssd1 vccd1 vccd1 _19308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19239_ _19401_/CLK _19239_/D vssd1 vssd1 vccd1 vccd1 _19239_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10437__S _10496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12218__A _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17487__A0 _17973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16124__S _16128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14433__A _14637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09527__A _18965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20014_ _20020_/CLK _20014_/D vssd1 vssd1 vccd1 vccd1 _20014_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10957__S0 _10937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input4_A io_dbus_rdata[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _10243_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _09825_/X sky130_fd_sc_hd__or2_1
XFILLER_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12888__A _12888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15264__A hold10/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ _09756_/A vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__buf_2
XFILLER_74_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _09787_/S vssd1 vssd1 vccd1 vccd1 _09726_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_27_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10185__S1 _10219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11382__S0 _10053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17411__A0 _17772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_139_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10600_ _09749_/A _10586_/X _10598_/X _09756_/A _10599_/Y vssd1 vssd1 vccd1 vccd1
+ _12651_/A sky130_fd_sc_hd__o32a_4
XFILLER_23_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11580_ _11580_/A _11580_/B _11580_/C vssd1 vssd1 vccd1 vccd1 _11580_/Y sky130_fd_sc_hd__nand3_1
XFILLER_80_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12251__A2 _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10531_ _10531_/A vssd1 vssd1 vccd1 vccd1 _10531_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10262__B2 _19914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13250_ _16865_/A _13202_/X _13203_/X _19687_/Q _13249_/X vssd1 vssd1 vccd1 vccd1
+ _13250_/X sky130_fd_sc_hd__a221o_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10462_ _10462_/A vssd1 vssd1 vccd1 vccd1 _10462_/X sky130_fd_sc_hd__buf_2
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11437__S1 _10691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17638__B _17642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12201_ _12201_/A _12201_/B vssd1 vssd1 vccd1 vccd1 _12203_/A sky130_fd_sc_hd__and2_1
XFILLER_164_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12562__S _12562_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13181_ input32/X _13172_/A _13175_/A vssd1 vssd1 vccd1 vccd1 _13194_/A sky130_fd_sc_hd__a21o_1
XANTENNA__16034__S _16034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10393_ _10393_/A _10393_/B vssd1 vssd1 vccd1 vccd1 _10393_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14343__A _14354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10871__A _11482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09437__A _18349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ _12127_/X _12129_/X _12130_/Y _12131_/X vssd1 vssd1 vccd1 vccd1 _12132_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15873__S _15879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16940_ _16940_/A vssd1 vssd1 vccd1 vccd1 _19741_/D sky130_fd_sc_hd__clkbuf_1
X_12063_ _19827_/Q vssd1 vssd1 vccd1 vccd1 _17180_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11014_ _11014_/A _11014_/B vssd1 vssd1 vccd1 vccd1 _11014_/X sky130_fd_sc_hd__or2_1
X_16871_ _16874_/A _16871_/B _16880_/D vssd1 vssd1 vccd1 vccd1 _19721_/D sky130_fd_sc_hd__nor3_1
XANTENNA__12798__A _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18610_ _19042_/CLK _18610_/D vssd1 vssd1 vccd1 vccd1 _18610_/Q sky130_fd_sc_hd__dfxtp_1
X_15822_ _15818_/X _18464_/Q _15819_/Y _15821_/X vssd1 vssd1 vccd1 vccd1 _15822_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19590_ _19594_/CLK _19590_/D vssd1 vssd1 vccd1 vccd1 _19590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18541_ _19196_/CLK _18541_/D vssd1 vssd1 vccd1 vccd1 _18541_/Q sky130_fd_sc_hd__dfxtp_1
X_15753_ _19908_/Q _15708_/X _16285_/A vssd1 vssd1 vccd1 vccd1 _15753_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _18454_/Q _12959_/X _11562_/A _12962_/X vssd1 vssd1 vccd1 vccd1 _18454_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ _14750_/S vssd1 vssd1 vccd1 vccd1 _14713_/S sky130_fd_sc_hd__buf_2
X_11916_ _19519_/Q _12120_/A vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__or2_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10111__A _10910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15684_ _15683_/X _19328_/Q _15684_/S vssd1 vssd1 vccd1 vccd1 _15685_/A sky130_fd_sc_hd__mux2_1
X_18472_ _19455_/CLK _18472_/D vssd1 vssd1 vccd1 vccd1 _18472_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _12995_/A vssd1 vssd1 vccd1 vccd1 _12896_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14634_/X _18882_/Q _14638_/S vssd1 vssd1 vccd1 vccd1 _14636_/A sky130_fd_sc_hd__mux2_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17423_ _17586_/S vssd1 vssd1 vccd1 vccd1 _17508_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_127_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11847_ _16213_/A _11846_/X _11668_/X vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _13841_/X _18860_/Q _14568_/S vssd1 vssd1 vccd1 vccd1 _14567_/A sky130_fd_sc_hd__mux2_1
X_17354_ _18335_/A _17342_/B _17358_/A _19886_/Q vssd1 vssd1 vccd1 vccd1 _17355_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11778_/A vssd1 vssd1 vccd1 vccd1 _12492_/A sky130_fd_sc_hd__buf_2
XFILLER_158_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13517_ _19639_/Q _12839_/X _13516_/X vssd1 vssd1 vccd1 vccd1 _13517_/X sky130_fd_sc_hd__o21a_1
X_16305_ _12127_/X _15764_/A _16300_/A vssd1 vssd1 vccd1 vccd1 _16305_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_174_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10729_ _18774_/Q _19045_/Q _19269_/Q _19013_/Q _10608_/X _10609_/X vssd1 vssd1 vccd1
+ vccd1 _10730_/B sky130_fd_sc_hd__mux4_1
XANTENNA__17829__A _17832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17285_ _12741_/X _19866_/Q _17291_/S vssd1 vssd1 vccd1 vccd1 _17286_/A sky130_fd_sc_hd__mux2_1
X_14497_ _14828_/A _18411_/B vssd1 vssd1 vccd1 vccd1 _18830_/D sky130_fd_sc_hd__nor2_4
XANTENNA__12038__A _12038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19024_ _19058_/CLK _19024_/D vssd1 vssd1 vccd1 vccd1 _19024_/Q sky130_fd_sc_hd__dfxtp_1
X_16236_ _19520_/Q _16235_/X _16252_/S vssd1 vssd1 vccd1 vccd1 _16237_/A sky130_fd_sc_hd__mux2_1
X_13448_ _16924_/C _13202_/X _13203_/X _19699_/Q _13447_/X vssd1 vssd1 vccd1 vccd1
+ _13448_/X sky130_fd_sc_hd__a221o_1
XFILLER_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16167_ _19498_/Q _14621_/A _16167_/S vssd1 vssd1 vccd1 vccd1 _16168_/A sky130_fd_sc_hd__mux2_1
X_13379_ _13379_/A vssd1 vssd1 vccd1 vccd1 _18489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18130__A1 _19958_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15118_ _15118_/A vssd1 vssd1 vccd1 vccd1 _15127_/S sky130_fd_sc_hd__buf_4
XFILLER_142_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12950__B1 _10961_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16098_ _13293_/X _19467_/Q _16106_/S vssd1 vssd1 vccd1 vccd1 _16099_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15049_ _19060_/Q _14456_/X _15055_/S vssd1 vssd1 vccd1 vccd1 _15050_/A sky130_fd_sc_hd__mux2_1
X_19926_ _19930_/CLK hold5/X vssd1 vssd1 vccd1 vccd1 _19926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19857_ _19857_/CLK _19857_/D vssd1 vssd1 vccd1 vccd1 _19857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14399__S _14402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09610_ _09610_/A vssd1 vssd1 vccd1 vccd1 _09611_/A sky130_fd_sc_hd__buf_2
X_18808_ _19497_/CLK _18808_/D vssd1 vssd1 vccd1 vccd1 _18808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12501__A _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19788_ _19789_/CLK _19788_/D vssd1 vssd1 vccd1 vccd1 _19788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09541_ _09761_/S vssd1 vssd1 vccd1 vccd1 _09542_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__13316__B _13316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18739_ _19200_/CLK _18739_/D vssd1 vssd1 vccd1 vccd1 _18739_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11808__A2 _11244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10167__S1 _10148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17503__S _17507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_140_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09472_ _09472_/A vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17944__A1 _19908_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13430__A1 _12921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15958__S _15962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clock _19998_/CLK vssd1 vssd1 vccd1 vccd1 _19963_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10691__A _10691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_65_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13497__B2 _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09808_ _18820_/Q _19155_/Q _10195_/S vssd1 vssd1 vccd1 vccd1 _09809_/B sky130_fd_sc_hd__mux2_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09739_ _09739_/A vssd1 vssd1 vccd1 vccd1 _09740_/A sky130_fd_sc_hd__buf_4
XANTENNA__16818__A _16818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12750_ _19723_/Q vssd1 vssd1 vccd1 vccd1 _16921_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_83_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11849_/B vssd1 vssd1 vccd1 vccd1 _11712_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12681_ _12693_/A vssd1 vssd1 vccd1 vccd1 _17146_/A sky130_fd_sc_hd__buf_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10866__A _19902_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14624_/A vssd1 vssd1 vccd1 vccd1 _14420_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _12475_/B vssd1 vssd1 vccd1 vccd1 _12568_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__13421__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14351_ _14351_/A vssd1 vssd1 vccd1 vccd1 _18786_/D sky130_fd_sc_hd__clkbuf_1
X_11563_ _11563_/A _11563_/B vssd1 vssd1 vccd1 vccd1 _11563_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13302_ _13534_/S _19909_/Q _13418_/A _13301_/X vssd1 vssd1 vccd1 vccd1 _13302_/X
+ sky130_fd_sc_hd__o211a_1
X_10514_ _10510_/X _10512_/X _10513_/X _10569_/A _09476_/A vssd1 vssd1 vccd1 vccd1
+ _10519_/B sky130_fd_sc_hd__o221a_1
XFILLER_10_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17070_ _19785_/Q _17070_/B _17070_/C vssd1 vssd1 vccd1 vccd1 _17072_/B sky130_fd_sc_hd__and3_1
X_14282_ _13831_/X _18756_/Q _14290_/S vssd1 vssd1 vccd1 vccd1 _14283_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11494_ _11494_/A vssd1 vssd1 vccd1 vccd1 _11494_/Y sky130_fd_sc_hd__inv_2
X_16021_ _13259_/X _19433_/Q _16023_/S vssd1 vssd1 vccd1 vccd1 _16022_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09928__A1 _09874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ _19905_/Q _12872_/B _13520_/S vssd1 vssd1 vccd1 vccd1 _13233_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11697__A _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ _10448_/A _10442_/X _10444_/X vssd1 vssd1 vccd1 vccd1 _10445_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13164_ _13468_/S _19901_/Q vssd1 vssd1 vccd1 vccd1 _13164_/X sky130_fd_sc_hd__or2_1
X_10376_ _09820_/A _10371_/X _10373_/X _10375_/X _09588_/A vssd1 vssd1 vccd1 vccd1
+ _10376_/X sky130_fd_sc_hd__a221o_2
XFILLER_124_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output166_A _12629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ _12537_/A vssd1 vssd1 vccd1 vccd1 _12115_/X sky130_fd_sc_hd__buf_2
XFILLER_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13095_ _13095_/A _13132_/C vssd1 vssd1 vccd1 vccd1 _13095_/Y sky130_fd_sc_hd__nor2_1
X_17972_ _17977_/B _17973_/B vssd1 vssd1 vccd1 vccd1 _17976_/B sky130_fd_sc_hd__and2b_1
XFILLER_97_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19711_ _19718_/CLK _19711_/D vssd1 vssd1 vccd1 vccd1 _19711_/Q sky130_fd_sc_hd__dfxtp_1
X_16923_ _19730_/Q _16923_/B _16923_/C _16923_/D vssd1 vssd1 vccd1 vccd1 _16924_/D
+ sky130_fd_sc_hd__and4_1
X_12046_ _12077_/S vssd1 vssd1 vccd1 vccd1 _12198_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15108__S _15116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19642_ _19877_/CLK _19642_/D vssd1 vssd1 vccd1 vccd1 _19642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16854_ _16868_/C _16868_/D vssd1 vssd1 vccd1 vccd1 _16856_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _18462_/Q _12853_/X _15804_/X vssd1 vssd1 vccd1 vccd1 _17225_/A sky130_fd_sc_hd__a21oi_1
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19573_ _19573_/CLK _19573_/D vssd1 vssd1 vccd1 vccd1 _19573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13997_ _13997_/A vssd1 vssd1 vccd1 vccd1 _18633_/D sky130_fd_sc_hd__clkbuf_1
X_16785_ _16818_/A _16790_/C vssd1 vssd1 vccd1 vccd1 _16785_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10149__S1 _10148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13851__S _13851_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18524_ _19501_/CLK _18524_/D vssd1 vssd1 vccd1 vccd1 _18524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15736_ _18450_/Q _15736_/B vssd1 vssd1 vccd1 vccd1 _15736_/X sky130_fd_sc_hd__or2_1
X_12948_ _18442_/Q _12946_/X _11082_/X _12947_/X vssd1 vssd1 vccd1 vccd1 _18442_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16447__B _16447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18455_ _19985_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15667_ _15667_/A vssd1 vssd1 vccd1 vccd1 _19324_/D sky130_fd_sc_hd__clkbuf_1
X_12879_ _14476_/A vssd1 vssd1 vccd1 vccd1 _12880_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12467__S _12562_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14248__A _14294_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ _17549_/A _17542_/D vssd1 vssd1 vccd1 vccd1 _17721_/C sky130_fd_sc_hd__nand2_2
XFILLER_159_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14618_ _14618_/A vssd1 vssd1 vccd1 vccd1 _14618_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17139__C1 _16480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15598_ _14586_/X _19293_/Q _15600_/S vssd1 vssd1 vccd1 vccd1 _15599_/A sky130_fd_sc_hd__mux2_1
X_18386_ _20031_/Q _18373_/X _18374_/X _18385_/Y vssd1 vssd1 vccd1 vccd1 _18387_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14549_ _13815_/X _18852_/Q _14557_/S vssd1 vssd1 vccd1 vccd1 _14550_/A sky130_fd_sc_hd__mux2_1
X_17337_ _17337_/A _17337_/B vssd1 vssd1 vccd1 vccd1 _17396_/B sky130_fd_sc_hd__or2_1
XFILLER_147_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18351__B2 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17268_ _17268_/A vssd1 vssd1 vccd1 vccd1 _19858_/D sky130_fd_sc_hd__clkbuf_1
X_19007_ _19487_/CLK _19007_/D vssd1 vssd1 vccd1 vccd1 _19007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16219_ _16219_/A _16219_/B _16219_/C vssd1 vssd1 vccd1 vccd1 _16232_/C sky130_fd_sc_hd__or3_2
X_17199_ _17199_/A _17210_/B vssd1 vssd1 vccd1 vccd1 _17199_/X sky130_fd_sc_hd__or2_1
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16402__S _16404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10016__A _10977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19909_ _19914_/CLK _19909_/D vssd1 vssd1 vccd1 vccd1 _19909_/Q sky130_fd_sc_hd__dfxtp_4
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10388__S1 _10440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16638__A _16672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13100__B1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11337__S0 _11026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ _19129_/Q _18895_/Q _19577_/Q _19225_/Q _09763_/S _09526_/A vssd1 vssd1 vccd1
+ vccd1 _09525_/B sky130_fd_sc_hd__mux4_1
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_141_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19485_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09439_/X _11824_/A _11790_/A _09448_/C _11827_/A vssd1 vssd1 vccd1 vccd1
+ _17342_/B sky130_fd_sc_hd__o221a_2
XFILLER_169_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09386_ _09394_/A _13136_/B _12702_/A _11833_/A vssd1 vssd1 vccd1 vccd1 _09392_/C
+ sky130_fd_sc_hd__nor4_1
XFILLER_12_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16373__A _16441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_156_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19769_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10230_ _19506_/Q _18918_/Q _18955_/Q _18529_/Q _10175_/S _09927_/A vssd1 vssd1 vccd1
+ vccd1 _10230_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ _10161_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10161_/X sky130_fd_sc_hd__and2_1
XFILLER_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14621__A _14621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14836__A1_N _18316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09715__A _10994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10092_ _10618_/A vssd1 vssd1 vccd1 vccd1 _10813_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13920_ _13841_/X _18599_/Q _13922_/S vssd1 vssd1 vccd1 vccd1 _13921_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13851_ _13850_/X _18570_/Q _13851_/S vssd1 vssd1 vccd1 vccd1 _13852_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14767__S _14775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12802_ _12802_/A vssd1 vssd1 vccd1 vccd1 _13154_/A sky130_fd_sc_hd__buf_2
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16570_ _19630_/Q _16572_/C _16569_/Y vssd1 vssd1 vccd1 vccd1 _19630_/D sky130_fd_sc_hd__o21a_1
X_13782_ _13782_/A vssd1 vssd1 vccd1 vccd1 _18548_/D sky130_fd_sc_hd__clkbuf_1
X_10994_ _10994_/A vssd1 vssd1 vccd1 vccd1 _10994_/X sky130_fd_sc_hd__buf_2
XFILLER_76_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_109_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19285_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09450__A _20050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15521_ _15521_/A vssd1 vssd1 vccd1 vccd1 _19258_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09310__A2 _14074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12733_ _19886_/Q _15819_/B vssd1 vssd1 vccd1 vccd1 _15700_/A sky130_fd_sc_hd__and2b_2
XFILLER_163_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09941__S0 _10218_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15452_ _19228_/Q _15206_/X _15456_/S vssd1 vssd1 vccd1 vccd1 _15453_/A sky130_fd_sc_hd__mux2_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18240_ _19975_/Q _12339_/B _18242_/S vssd1 vssd1 vccd1 vccd1 _18241_/A sky130_fd_sc_hd__mux2_1
X_12664_ _12664_/A vssd1 vssd1 vccd1 vccd1 _12669_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_31_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14403_/A vssd1 vssd1 vccd1 vccd1 _18804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15598__S _15600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11615_ _11615_/A vssd1 vssd1 vccd1 vccd1 _11854_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15383_ _15383_/A vssd1 vssd1 vccd1 vccd1 _19197_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17379__A _17379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18171_ _18171_/A vssd1 vssd1 vccd1 vccd1 _19944_/D sky130_fd_sc_hd__clkbuf_1
X_12595_ _12600_/A _12595_/B _12595_/C vssd1 vssd1 vccd1 vccd1 _12595_/X sky130_fd_sc_hd__or3_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14334_ _14334_/A vssd1 vssd1 vccd1 vccd1 _18778_/D sky130_fd_sc_hd__clkbuf_1
X_17122_ _17122_/A _17122_/B _17122_/C vssd1 vssd1 vccd1 vccd1 _19803_/D sky130_fd_sc_hd__nor3_1
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11546_ _11548_/A _11550_/A _11548_/C _12662_/B _10144_/A vssd1 vssd1 vccd1 vccd1
+ _11546_/X sky130_fd_sc_hd__a32o_1
XFILLER_156_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17053_ _19779_/Q _17053_/B _17053_/C vssd1 vssd1 vccd1 vccd1 _17055_/B sky130_fd_sc_hd__and3_1
XFILLER_171_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14265_ _14265_/A vssd1 vssd1 vccd1 vccd1 _18748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11477_ _18665_/Q _19256_/Q _19418_/Q _18633_/Q _09967_/A _10074_/A vssd1 vssd1 vccd1
+ vccd1 _11478_/B sky130_fd_sc_hd__mux4_1
XFILLER_100_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14007__S _14013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09609__B _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16004_ _13109_/X _19425_/Q _16012_/S vssd1 vssd1 vccd1 vccd1 _16005_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13216_ _13363_/A _13212_/X _13215_/X vssd1 vssd1 vccd1 vccd1 _13216_/X sky130_fd_sc_hd__a21bo_1
XFILLER_171_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10428_ _10428_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10428_/X sky130_fd_sc_hd__or2_1
X_14196_ _13812_/X _18718_/Q _14196_/S vssd1 vssd1 vccd1 vccd1 _14197_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13133_/Y _13146_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13147_/X sky130_fd_sc_hd__mux2_1
X_10359_ _10349_/Y _10353_/Y _10356_/Y _10358_/Y _09719_/A vssd1 vssd1 vccd1 vccd1
+ _10359_/X sky130_fd_sc_hd__o221a_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _19328_/Q _12864_/X _12756_/A _19518_/Q _13077_/X vssd1 vssd1 vccd1 vccd1
+ _13078_/X sky130_fd_sc_hd__a221o_1
X_17955_ _12234_/B _17755_/X _17954_/X _17778_/X vssd1 vssd1 vccd1 vccd1 _17955_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_97_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16906_ _19733_/Q _19732_/Q _19731_/Q _16906_/D vssd1 vssd1 vccd1 vccd1 _16915_/D
+ sky130_fd_sc_hd__and4_1
X_12029_ _12086_/C _12153_/B _12029_/C _12029_/D vssd1 vssd1 vccd1 vccd1 _12029_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17886_ _17533_/X _17877_/X _17885_/X _18054_/A vssd1 vssd1 vccd1 vccd1 _17886_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19625_ _19759_/CLK _19625_/D vssd1 vssd1 vccd1 vccd1 _19625_/Q sky130_fd_sc_hd__dfxtp_1
X_16837_ _19712_/Q _16848_/C _16833_/X vssd1 vssd1 vccd1 vccd1 _16838_/B sky130_fd_sc_hd__o21ai_1
XFILLER_66_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12986__A _13173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16458__A _18404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__A _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19556_ _19556_/CLK _19556_/D vssd1 vssd1 vccd1 vccd1 _19556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16768_ _16860_/A vssd1 vssd1 vccd1 vccd1 _16768_/X sky130_fd_sc_hd__buf_2
XFILLER_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18507_ _19258_/CLK _18507_/D vssd1 vssd1 vccd1 vccd1 _18507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_13_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15719_ _19902_/Q _15718_/X _15719_/S vssd1 vssd1 vccd1 vccd1 _15719_/X sky130_fd_sc_hd__mux2_1
X_19487_ _19487_/CLK _19487_/D vssd1 vssd1 vccd1 vccd1 _19487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16699_ _19785_/Q _19784_/Q _19786_/Q _17065_/A vssd1 vssd1 vccd1 vccd1 _17074_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_21_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09240_ _09272_/C _09269_/B _09266_/B vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__or3_1
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18438_ _19956_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_73_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19449_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ _20024_/Q vssd1 vssd1 vccd1 vccd1 _18279_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18369_ _18380_/A _18369_/B vssd1 vssd1 vccd1 vccd1 _20026_/D sky130_fd_sc_hd__nor2_1
XFILLER_147_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13610__A _14844_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_88_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _18777_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13756__S _13765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16132__S _16132_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_clock _19998_/CLK vssd1 vssd1 vccd1 vccd1 _19592_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09535__A _10509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12124__A1 _19526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10686__A1 _11440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10230__S0 _10175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19051_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14587__S _14590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10781__S1 _11496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09507_ _10244_/S vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__clkbuf_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17366__A2 _18301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _18333_/A _11640_/A _11730_/B _11640_/C vssd1 vssd1 vccd1 vccd1 _09453_/B
+ sky130_fd_sc_hd__or4_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _20014_/Q vssd1 vssd1 vccd1 vccd1 _12688_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _19465_/Q _19303_/Q _18712_/Q _18482_/Q _10053_/X _10054_/X vssd1 vssd1 vccd1
+ vccd1 _11400_/X sky130_fd_sc_hd__mux4_2
XANTENNA__18431__A1_N _18347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12380_ _12322_/A _12324_/B _18012_/A _12429_/A vssd1 vssd1 vccd1 vccd1 _12382_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11331_ _10024_/A _11328_/Y _11330_/Y _11295_/A vssd1 vssd1 vccd1 vccd1 _11331_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10049__S0 _11451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14050_ _14050_/A vssd1 vssd1 vccd1 vccd1 _18655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _18965_/Q vssd1 vssd1 vccd1 vccd1 _11262_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13001_ _09341_/X _13569_/B _13553_/S vssd1 vssd1 vccd1 vccd1 _13001_/X sky130_fd_sc_hd__mux2_1
X_10213_ _10209_/A _10210_/X _10212_/X _09826_/X vssd1 vssd1 vccd1 vccd1 _10213_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15447__A _15515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11193_ _19100_/Q _18866_/Q _19548_/Q _19196_/Q _09981_/A _11260_/A vssd1 vssd1 vccd1
+ vccd1 _11193_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input42_A io_ibus_inst[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _10144_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _10145_/B sky130_fd_sc_hd__or2_1
XFILLER_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17740_ _17740_/A vssd1 vssd1 vccd1 vccd1 _17740_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_153_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10075_ _19125_/Q _18891_/Q _19573_/Q _19221_/Q _10073_/X _10609_/A vssd1 vssd1 vccd1
+ vccd1 _10075_/X sky130_fd_sc_hd__mux4_1
X_14952_ _14974_/A vssd1 vssd1 vccd1 vccd1 _14961_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_130_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11323__C1 _09617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13903_ _13815_/X _18591_/Q _13911_/S vssd1 vssd1 vccd1 vccd1 _13904_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10221__S0 _09653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17671_ _19895_/Q _17670_/X _17808_/S vssd1 vssd1 vccd1 vccd1 _17672_/A sky130_fd_sc_hd__mux2_1
X_14883_ _14628_/X _18986_/Q _14889_/S vssd1 vssd1 vccd1 vccd1 _14884_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output129_A _12667_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19410_ _19411_/CLK _19410_/D vssd1 vssd1 vccd1 vccd1 _19410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16622_ _19648_/Q _16619_/B _16621_/Y vssd1 vssd1 vccd1 vccd1 _19648_/D sky130_fd_sc_hd__o21a_1
X_13834_ _13834_/A vssd1 vssd1 vccd1 vccd1 _18564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19341_ _19873_/CLK _19341_/D vssd1 vssd1 vccd1 vccd1 _19341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16553_ _19624_/Q _16555_/C _16552_/Y vssd1 vssd1 vccd1 vccd1 _19624_/D sky130_fd_sc_hd__o21a_1
X_13765_ _13764_/X _18543_/Q _13765_/S vssd1 vssd1 vccd1 vccd1 _13766_/A sky130_fd_sc_hd__mux2_1
X_10977_ _10977_/A vssd1 vssd1 vccd1 vccd1 _11224_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_187_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15504_ _15504_/A vssd1 vssd1 vccd1 vccd1 _19251_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17601__S _17601_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19272_ _19272_/CLK _19272_/D vssd1 vssd1 vccd1 vccd1 _19272_/Q sky130_fd_sc_hd__dfxtp_1
X_12716_ _19626_/Q _13142_/B _12715_/X vssd1 vssd1 vccd1 vccd1 _13301_/B sky130_fd_sc_hd__o21a_2
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13696_ _15263_/A vssd1 vssd1 vccd1 vccd1 _14640_/A sky130_fd_sc_hd__buf_2
X_16484_ _19600_/Q _16477_/X _12397_/X _12400_/Y _16482_/X vssd1 vssd1 vccd1 vccd1
+ _19600_/D sky130_fd_sc_hd__o221a_1
X_18223_ _19967_/Q _12086_/A _18231_/S vssd1 vssd1 vccd1 vccd1 _18224_/A sky130_fd_sc_hd__mux2_1
X_15435_ _14663_/X _19221_/Q _15439_/S vssd1 vssd1 vccd1 vccd1 _15436_/A sky130_fd_sc_hd__mux2_1
X_12647_ _12647_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _12647_/Y sky130_fd_sc_hd__nor2_4
XFILLER_129_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14526__A _14572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15121__S _15127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15366_ _15366_/A vssd1 vssd1 vccd1 vccd1 _19190_/D sky130_fd_sc_hd__clkbuf_1
X_18154_ _18154_/A vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__clkbuf_1
X_12578_ _12532_/A _12535_/A _12555_/A _12556_/Y vssd1 vssd1 vccd1 vccd1 _12579_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17105_ _17104_/B _17104_/C _19797_/Q vssd1 vssd1 vccd1 vccd1 _17106_/C sky130_fd_sc_hd__a21oi_1
XFILLER_129_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11529_ _11524_/Y _11519_/B _11534_/B _11528_/X vssd1 vssd1 vccd1 vccd1 _11530_/C
+ sky130_fd_sc_hd__a31o_1
X_14317_ _18771_/Q _13647_/X _14319_/S vssd1 vssd1 vccd1 vccd1 _14318_/A sky130_fd_sc_hd__mux2_1
X_15297_ _15297_/A vssd1 vssd1 vccd1 vccd1 _19160_/D sky130_fd_sc_hd__clkbuf_1
X_18085_ _19920_/Q _18084_/X _18085_/S vssd1 vssd1 vccd1 vccd1 _18086_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14248_ _14294_/S vssd1 vssd1 vccd1 vccd1 _14257_/S sky130_fd_sc_hd__buf_4
X_17036_ hold20/A _17034_/C _17035_/Y vssd1 vssd1 vccd1 vccd1 _19768_/D sky130_fd_sc_hd__o21a_1
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14179_ _13787_/X _18710_/Q _14185_/S vssd1 vssd1 vccd1 vccd1 _14180_/A sky130_fd_sc_hd__mux2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _19308_/CLK _18987_/D vssd1 vssd1 vccd1 vccd1 _18987_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _18000_/A _17935_/X _17937_/X _17533_/A vssd1 vssd1 vccd1 vccd1 _17938_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17869_ _18083_/A vssd1 vssd1 vccd1 vccd1 _17869_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10763__S1 _10030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19608_ _19608_/CLK _19608_/D vssd1 vssd1 vccd1 vccd1 _19608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19539_ _19540_/CLK _19539_/D vssd1 vssd1 vccd1 vccd1 _19539_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10515__S1 _10462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ _20035_/Q vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14436__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15031__S _15033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clock clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_163_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10175__S _10175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14870__S _14878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17808__A0 _19900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15267__A _15267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10451__S0 _10337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09987_ _10732_/A _09987_/B vssd1 vssd1 vccd1 vccd1 _09987_/X sky130_fd_sc_hd__or2_1
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17482__A _17581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16492__C1 _12749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18297__B _18326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11856__A0 _11899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10900_ _18827_/Q vssd1 vssd1 vccd1 vccd1 _11035_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11880_ _19816_/Q _19849_/Q vssd1 vssd1 vccd1 vccd1 _11881_/D sky130_fd_sc_hd__nand2_1
XFILLER_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10831_ _18580_/Q _18841_/Q _18740_/Q _19075_/Q _09532_/A _09514_/A vssd1 vssd1 vccd1
+ vccd1 _10832_/B sky130_fd_sc_hd__mux4_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11035__A _11035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ _19641_/Q _12861_/X _13549_/X vssd1 vssd1 vccd1 vccd1 _13550_/X sky130_fd_sc_hd__o21a_1
X_10762_ _10655_/X _10755_/X _10757_/Y _10761_/Y _09739_/A vssd1 vssd1 vccd1 vccd1
+ _10762_/X sky130_fd_sc_hd__o311a_2
XFILLER_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12501_ _12501_/A vssd1 vssd1 vccd1 vccd1 _18079_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13481_ _19733_/Q _13341_/X _13342_/X _19701_/Q _13480_/X vssd1 vssd1 vccd1 vccd1
+ _13481_/X sky130_fd_sc_hd__a221o_1
X_10693_ _10632_/A _10692_/X _09475_/A vssd1 vssd1 vccd1 vccd1 _10693_/X sky130_fd_sc_hd__o21a_1
XANTENNA__16037__S _16045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15220_ _19136_/Q _15219_/X _15229_/S vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__mux2_1
X_12432_ _12432_/A vssd1 vssd1 vccd1 vccd1 _18046_/B sky130_fd_sc_hd__buf_2
XFILLER_32_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15770__B2 _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15151_ _19107_/Q vssd1 vssd1 vccd1 vccd1 _15152_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_148_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12363_ _12537_/A vssd1 vssd1 vccd1 vccd1 _12363_/X sky130_fd_sc_hd__buf_2
XANTENNA__14780__S _14786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _14102_/A vssd1 vssd1 vccd1 vccd1 _18677_/D sky130_fd_sc_hd__clkbuf_1
X_11314_ _18635_/Q _19226_/Q _19388_/Q _18603_/Q _10999_/A _11065_/A vssd1 vssd1 vccd1
+ vccd1 _11315_/B sky130_fd_sc_hd__mux4_2
X_15082_ _15082_/A vssd1 vssd1 vccd1 vccd1 _19074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12294_ _17205_/A _12316_/C vssd1 vssd1 vccd1 vccd1 _12294_/X sky130_fd_sc_hd__or2_1
X_18910_ _19498_/CLK _18910_/D vssd1 vssd1 vccd1 vccd1 _18910_/Q sky130_fd_sc_hd__dfxtp_1
X_14033_ _18648_/Q _13668_/X _14035_/S vssd1 vssd1 vccd1 vccd1 _14034_/A sky130_fd_sc_hd__mux2_1
X_11245_ _19359_/Q _18973_/Q _19423_/Q _18542_/Q _11129_/X _11115_/A vssd1 vssd1 vccd1
+ vccd1 _11246_/B sky130_fd_sc_hd__mux4_1
X_19890_ _20000_/CLK _19890_/D vssd1 vssd1 vccd1 vccd1 _19890_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10442__S0 _10337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10898__A1 _09612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18841_ _19203_/CLK _18841_/D vssd1 vssd1 vccd1 vccd1 _18841_/Q sky130_fd_sc_hd__dfxtp_1
X_11176_ _09703_/A _11163_/Y _11169_/X _11175_/Y _09736_/A vssd1 vssd1 vccd1 vccd1
+ _11176_/X sky130_fd_sc_hd__o311a_2
XANTENNA__10898__B2 _19901_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10127_ _09680_/A _10126_/X _09693_/A vssd1 vssd1 vccd1 vccd1 _10127_/Y sky130_fd_sc_hd__o21ai_1
X_18772_ _19556_/CLK _18772_/D vssd1 vssd1 vccd1 vccd1 _18772_/Q sky130_fd_sc_hd__dfxtp_1
X_15984_ _19417_/Q _15292_/X _15984_/S vssd1 vssd1 vccd1 vccd1 _15985_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10114__A _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09903__A _10368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17723_ _17723_/A vssd1 vssd1 vccd1 vccd1 _17723_/X sky130_fd_sc_hd__clkbuf_2
X_10058_ _10790_/A vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__clkbuf_4
X_14935_ _19009_/Q _14395_/X _14939_/S vssd1 vssd1 vccd1 vccd1 _14936_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17542__D _17542_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15116__S _15116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10745__S1 _10682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17654_ _17803_/S _17654_/B vssd1 vssd1 vccd1 vccd1 _17654_/X sky130_fd_sc_hd__or2_1
XANTENNA__14020__S _14024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14866_ _14866_/A vssd1 vssd1 vccd1 vccd1 _18978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16605_ _19642_/Q vssd1 vssd1 vccd1 vccd1 _16609_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13817_ _13815_/X _18559_/Q _13829_/S vssd1 vssd1 vccd1 vccd1 _13818_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14955__S _14961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17585_ _17581_/X _17584_/X _17759_/S vssd1 vssd1 vccd1 vccd1 _17585_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14797_ _18952_/Q _14433_/X _14797_/S vssd1 vssd1 vccd1 vccd1 _14798_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19324_ _19852_/CLK _19324_/D vssd1 vssd1 vccd1 vccd1 _19324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16536_ _16635_/A vssd1 vssd1 vccd1 vccd1 _16573_/A sky130_fd_sc_hd__buf_2
X_13748_ _19887_/Q _13748_/B vssd1 vssd1 vccd1 vccd1 _14844_/D sky130_fd_sc_hd__nand2_1
XANTENNA__12811__A2 _12888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19255_ _19417_/CLK _19255_/D vssd1 vssd1 vccd1 vccd1 _19255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16467_ _12095_/A _12095_/B _16455_/X vssd1 vssd1 vccd1 vccd1 _19589_/D sky130_fd_sc_hd__a21o_1
XFILLER_148_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13679_ _13679_/A vssd1 vssd1 vccd1 vccd1 _18522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18206_ _18206_/A vssd1 vssd1 vccd1 vccd1 _19959_/D sky130_fd_sc_hd__clkbuf_1
X_15418_ _15418_/A vssd1 vssd1 vccd1 vccd1 _19213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19186_ _19412_/CLK _19186_/D vssd1 vssd1 vccd1 vccd1 _19186_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15761__A1 _12772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11599__B _17331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16398_ _13230_/X _19557_/Q _16404_/S vssd1 vssd1 vccd1 vccd1 _16399_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18137_ _18137_/A vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15349_ _15349_/A vssd1 vssd1 vccd1 vccd1 _19182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16471__A _18352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18068_ _18068_/A _18068_/B vssd1 vssd1 vccd1 vccd1 _18068_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09910_ _09833_/A _09909_/X _09580_/A vssd1 vssd1 vccd1 vccd1 _09910_/X sky130_fd_sc_hd__o21a_1
X_17019_ _19762_/Q _17014_/C _17018_/Y vssd1 vssd1 vccd1 vccd1 _19762_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09841_ _09841_/A vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20030_ _20032_/CLK _20030_/D vssd1 vssd1 vccd1 vccd1 _20030_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10984__S1 _11225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _19384_/Q _18998_/Q _19448_/Q _18567_/Q _09568_/X _09762_/A vssd1 vssd1 vccd1
+ vccd1 _09773_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13288__C1 _13287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10024__A _10024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__A _09813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13054__B _16206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09206_ _09275_/C vssd1 vssd1 vccd1 vccd1 _12610_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_167_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11302__B _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10577__B1 _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15709__B _15709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_135_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13515__B1 _13099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11030_ _11030_/A vssd1 vssd1 vccd1 vccd1 _11083_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_1_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13944__S _13950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10975__S1 _10974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12981_ _18465_/Q _12980_/X _11537_/A _12976_/X vssd1 vssd1 vccd1 vccd1 _18465_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10869__A _10869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _18913_/Q _14427_/X _14724_/S vssd1 vssd1 vccd1 vccd1 _14721_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13245__A _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11932_ _11932_/A _11969_/A vssd1 vssd1 vccd1 vccd1 _11938_/A sky130_fd_sc_hd__xor2_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _14650_/X _18887_/Q _14654_/S vssd1 vssd1 vccd1 vccd1 _14652_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11863_ _11933_/A _11933_/B vssd1 vssd1 vccd1 vccd1 _11864_/A sky130_fd_sc_hd__xnor2_4
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14775__S _14775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _10825_/A _10811_/X _10813_/X _10613_/A vssd1 vssd1 vccd1 vccd1 _10814_/X
+ sky130_fd_sc_hd__a211o_1
X_13602_ _13580_/A _13600_/X _13601_/Y _12903_/A _18468_/Q vssd1 vssd1 vccd1 vccd1
+ _13603_/B sky130_fd_sc_hd__a32o_4
XFILLER_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _17373_/A _17370_/B vssd1 vssd1 vccd1 vccd1 _17371_/A sky130_fd_sc_hd__and2_1
X_14582_ _14582_/A vssd1 vssd1 vccd1 vccd1 _18865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11794_ _19323_/D _11665_/B _11868_/C _11792_/Y _12584_/B vssd1 vssd1 vccd1 vccd1
+ _11794_/Y sky130_fd_sc_hd__o41ai_1
XFILLER_14_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11152__S1 _10024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16321_ _19945_/Q _19946_/Q _19947_/Q _16321_/D vssd1 vssd1 vccd1 vccd1 _16332_/C
+ sky130_fd_sc_hd__or4_4
X_10745_ _18646_/Q _19237_/Q _19399_/Q _18614_/Q _10617_/X _10682_/A vssd1 vssd1 vccd1
+ vccd1 _10746_/B sky130_fd_sc_hd__mux4_1
X_13533_ _19847_/Q _12696_/X _13529_/X _13530_/X _13532_/X vssd1 vssd1 vccd1 vccd1
+ _13533_/X sky130_fd_sc_hd__a2111o_4
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19040_ _19042_/CLK _19040_/D vssd1 vssd1 vccd1 vccd1 _19040_/Q sky130_fd_sc_hd__dfxtp_1
X_13464_ _19764_/Q _12840_/X _13463_/X _12846_/X vssd1 vssd1 vccd1 vccd1 _13464_/X
+ sky130_fd_sc_hd__a211o_1
X_16252_ _19523_/Q _16251_/X _16252_/S vssd1 vssd1 vccd1 vccd1 _16253_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10676_ _19110_/Q _18876_/Q _19558_/Q _19206_/Q _10675_/X _09957_/X vssd1 vssd1 vccd1
+ vccd1 _10677_/B sky130_fd_sc_hd__mux4_1
XANTENNA__15743__A1 _18451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15203_ _15203_/A vssd1 vssd1 vccd1 vccd1 _15203_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12415_ _19601_/Q vssd1 vssd1 vccd1 vccd1 _12416_/A sky130_fd_sc_hd__clkbuf_2
X_13395_ _13395_/A vssd1 vssd1 vccd1 vccd1 _18490_/D sky130_fd_sc_hd__clkbuf_1
X_16183_ _19505_/Q _14644_/A _16189_/S vssd1 vssd1 vccd1 vccd1 _16184_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17496__A1 _11969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15134_ _15134_/A vssd1 vssd1 vccd1 vccd1 _19098_/D sky130_fd_sc_hd__clkbuf_1
X_12346_ _17210_/A _12373_/C _12345_/Y vssd1 vssd1 vccd1 vccd1 _12346_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15065_ _15065_/A vssd1 vssd1 vccd1 vccd1 _19066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19942_ _19981_/CLK _19942_/D vssd1 vssd1 vccd1 vccd1 _19942_/Q sky130_fd_sc_hd__dfxtp_1
X_12277_ _12278_/A _17452_/A vssd1 vssd1 vccd1 vccd1 _12279_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14016_ _18640_/Q _13634_/X _14024_/S vssd1 vssd1 vccd1 vccd1 _14017_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output73_A _12084_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ _18766_/Q _19037_/Q _19261_/Q _19005_/Q _11161_/X _11179_/X vssd1 vssd1 vccd1
+ vccd1 _11228_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19873_ _19873_/CLK _19873_/D vssd1 vssd1 vccd1 vccd1 _19873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15635__A _15646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18824_ _19317_/CLK _18824_/D vssd1 vssd1 vccd1 vccd1 _18824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11159_ _11082_/X _12637_/B _11135_/X _12636_/B vssd1 vssd1 vccd1 vccd1 _11582_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18755_ _19570_/CLK _18755_/D vssd1 vssd1 vccd1 vccd1 _18755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15967_ _19409_/Q _15267_/X _15973_/S vssd1 vssd1 vccd1 vccd1 _15968_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17706_ _17697_/X _17701_/X _17703_/Y _17705_/X vssd1 vssd1 vccd1 vccd1 _17706_/X
+ sky130_fd_sc_hd__o211a_1
X_14918_ _14974_/A vssd1 vssd1 vccd1 vccd1 _14987_/S sky130_fd_sc_hd__buf_6
X_18686_ _19407_/CLK _18686_/D vssd1 vssd1 vccd1 vccd1 _18686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15898_ _15898_/A vssd1 vssd1 vccd1 vccd1 _19378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17420__A1 _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17637_ _17803_/S _17642_/B vssd1 vssd1 vccd1 vccd1 _17637_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14685__S _14691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14849_ _14849_/A vssd1 vssd1 vccd1 vccd1 _18970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11048__A1 _11216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17568_ _17448_/X _17484_/X _17582_/S vssd1 vssd1 vccd1 vccd1 _17568_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19307_ _19308_/CLK _19307_/D vssd1 vssd1 vccd1 vccd1 _19307_/Q sky130_fd_sc_hd__dfxtp_1
X_16519_ _16528_/A _16519_/B _16519_/C vssd1 vssd1 vccd1 vccd1 _19613_/D sky130_fd_sc_hd__nor3_1
XFILLER_32_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17499_ _12501_/A _17729_/B _17506_/S vssd1 vssd1 vccd1 vccd1 _17499_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11403__A hold15/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19238_ _19402_/CLK _19238_/D vssd1 vssd1 vccd1 vccd1 _19238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18831__D _18831_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19169_ _19394_/CLK _19169_/D vssd1 vssd1 vccd1 vccd1 _19169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10019__A _10040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17487__A1 _17899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10406__S0 _10268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20013_ _20020_/CLK _20013_/D vssd1 vssd1 vccd1 vccd1 _20013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10957__S1 _09954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ _18596_/Q _18857_/Q _18756_/Q _19091_/Q _10245_/S _09899_/A vssd1 vssd1 vccd1
+ vccd1 _09825_/B sky130_fd_sc_hd__mux4_1
XFILLER_100_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09755_ _09755_/A vssd1 vssd1 vccd1 vccd1 _09756_/A sky130_fd_sc_hd__buf_4
XFILLER_101_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10709__S1 _10665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09686_ _10188_/A vssd1 vssd1 vccd1 vccd1 _09699_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17411__A1 _12455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11382__S1 _10054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15280__A hold10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11039__A1 _11046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_61_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13004__S _13554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10530_ _18683_/Q _19178_/Q _10589_/S vssd1 vssd1 vccd1 vccd1 _10531_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13939__S _13939_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10461_ _10461_/A vssd1 vssd1 vccd1 vccd1 _10462_/A sky130_fd_sc_hd__buf_2
XFILLER_108_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14624__A _14624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12200_ _12229_/A _17447_/A vssd1 vssd1 vccd1 vccd1 _12201_/B sky130_fd_sc_hd__or2_1
XANTENNA__09718__A _09718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ _13180_/A vssd1 vssd1 vccd1 vccd1 _18477_/D sky130_fd_sc_hd__clkbuf_1
X_10392_ _18814_/Q _19149_/Q _10392_/S vssd1 vssd1 vccd1 vccd1 _10393_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12131_ _12247_/A vssd1 vssd1 vccd1 vccd1 _12131_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09437__B _18347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16150__A1 _14596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12062_ _12057_/Y _12060_/X _12061_/X vssd1 vssd1 vccd1 vccd1 _12062_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11013_ _19362_/Q _18976_/Q _19426_/Q _18545_/Q _10893_/X _09955_/A vssd1 vssd1 vccd1
+ vccd1 _11014_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16050__S _16056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16870_ _19721_/Q _19720_/Q _19719_/Q _16870_/D vssd1 vssd1 vccd1 vccd1 _16880_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__16989__B1 _16860_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15821_ _18464_/Q _13483_/B _15820_/Y _13587_/A vssd1 vssd1 vccd1 vccd1 _15821_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10599__A _19908_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15661__A0 _09341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18540_ _19734_/CLK _18540_/D vssd1 vssd1 vccd1 vccd1 _18540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _15806_/A _17194_/A vssd1 vssd1 vccd1 vccd1 _16285_/A sky130_fd_sc_hd__nor2_1
XFILLER_46_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _18453_/Q _12959_/X _10555_/A _12962_/X vssd1 vssd1 vccd1 vccd1 _18453_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _14703_/A vssd1 vssd1 vccd1 vccd1 _18905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _19794_/CLK _18471_/D vssd1 vssd1 vccd1 vccd1 _18471_/Q sky130_fd_sc_hd__dfxtp_1
X_11915_ _11915_/A vssd1 vssd1 vccd1 vccd1 _12120_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output111_A _12647_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15683_ _19897_/Q _15668_/X _16222_/A vssd1 vssd1 vccd1 vccd1 _15683_/X sky130_fd_sc_hd__a21o_1
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _19873_/Q _12755_/A _12696_/A _19840_/Q _12894_/X vssd1 vssd1 vccd1 vccd1
+ _12895_/X sky130_fd_sc_hd__a221o_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17422_ _17749_/B _12480_/A _17450_/S vssd1 vssd1 vccd1 vccd1 _17422_/X sky130_fd_sc_hd__mux2_1
X_14634_ _14634_/A vssd1 vssd1 vccd1 vccd1 _14634_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _11958_/B _11843_/X _11844_/Y _11845_/X vssd1 vssd1 vccd1 vccd1 _11846_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _18273_/S vssd1 vssd1 vccd1 vccd1 _18335_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _14565_/A vssd1 vssd1 vccd1 vccd1 _18859_/D sky130_fd_sc_hd__clkbuf_1
X_11777_ _11958_/B vssd1 vssd1 vccd1 vccd1 _11957_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12319__A _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _16308_/B _16302_/Y _16303_/X vssd1 vssd1 vccd1 vccd1 _16304_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13516_ _19767_/Q _12692_/A _13515_/X _12714_/A vssd1 vssd1 vccd1 vccd1 _13516_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10728_ _10728_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _11570_/A sky130_fd_sc_hd__and2_1
XFILLER_158_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17284_ _17284_/A vssd1 vssd1 vccd1 vccd1 _19865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17829__B _17832_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14496_ _18331_/A _16811_/A _14481_/X _14495_/Y vssd1 vssd1 vccd1 vccd1 _18411_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_174_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19023_ _19504_/CLK _19023_/D vssd1 vssd1 vccd1 vccd1 _19023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16235_ _16235_/A _16235_/B vssd1 vssd1 vccd1 vccd1 _16235_/X sky130_fd_sc_hd__or2_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10659_ _19370_/Q _18984_/Q _19434_/Q _18553_/Q _10658_/X _10014_/X vssd1 vssd1 vccd1
+ vccd1 _10660_/B sky130_fd_sc_hd__mux4_1
XFILLER_158_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13447_ _19635_/Q _12839_/X _13446_/X vssd1 vssd1 vccd1 vccd1 _13447_/X sky130_fd_sc_hd__o21a_1
XFILLER_139_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09628__A _10899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ _18489_/Q _13376_/X _13434_/S vssd1 vssd1 vccd1 vccd1 _13379_/A sky130_fd_sc_hd__mux2_1
X_16166_ _16166_/A vssd1 vssd1 vccd1 vccd1 _19497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15117_ _15117_/A vssd1 vssd1 vccd1 vccd1 _19090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12329_ _12329_/A _18001_/B vssd1 vssd1 vccd1 vccd1 _12330_/B sky130_fd_sc_hd__nor2_1
XFILLER_170_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16097_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16106_/S sky130_fd_sc_hd__buf_2
XFILLER_141_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15048_ _15048_/A vssd1 vssd1 vccd1 vccd1 _19059_/D sky130_fd_sc_hd__clkbuf_1
X_19925_ _19930_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 _19925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12989__A _12989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11893__A _11893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19856_ _19859_/CLK _19856_/D vssd1 vssd1 vccd1 vccd1 _19856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18807_ _19495_/CLK _18807_/D vssd1 vssd1 vccd1 vccd1 _18807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19787_ _19789_/CLK _19787_/D vssd1 vssd1 vccd1 vccd1 _19787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16999_ _17005_/C _17003_/C _16860_/X vssd1 vssd1 vccd1 vccd1 _16999_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09540_ _10162_/S vssd1 vssd1 vccd1 vccd1 _09761_/S sky130_fd_sc_hd__buf_2
XFILLER_110_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18738_ _19553_/CLK _18738_/D vssd1 vssd1 vccd1 vccd1 _18738_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10302__A _10559_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11808__A3 _11253_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09471_ _10875_/A vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__buf_2
X_18669_ _19484_/CLK _18669_/D vssd1 vssd1 vccd1 vccd1 _18669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13613__A _13719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13759__S _13765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18106__C1 _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09538__A _10416_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10401__C1 _09741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17880__A1 _17884_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13497__A2 _12992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09807_ _09807_/A vssd1 vssd1 vccd1 vccd1 _09807_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09738_ _09738_/A vssd1 vssd1 vccd1 vccd1 _09739_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15722__B _15722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ _09927_/A vssd1 vssd1 vccd1 vccd1 _10176_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13523__A _15292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11894_/A _12631_/B _11696_/X _11699_/X vssd1 vssd1 vccd1 vccd1 _11849_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12680_ _17247_/D vssd1 vssd1 vccd1 vccd1 _12684_/B sky130_fd_sc_hd__clkinv_2
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _17325_/A _12595_/B vssd1 vssd1 vccd1 vccd1 _11636_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14350_ _18786_/Q _13710_/X _14352_/S vssd1 vssd1 vccd1 vccd1 _14351_/A sky130_fd_sc_hd__mux2_1
X_11562_ _11562_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _11563_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10513_ _19114_/Q _18880_/Q _19562_/Q _19210_/Q _10470_/X _10462_/A vssd1 vssd1 vccd1
+ vccd1 _10513_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13669__S _13673_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13301_ _13316_/A _13301_/B _13301_/C _13301_/D vssd1 vssd1 vccd1 vccd1 _13301_/X
+ sky130_fd_sc_hd__or4_2
X_14281_ _14281_/A vssd1 vssd1 vccd1 vccd1 _14290_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16045__S _16045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11493_ _18697_/Q _19192_/Q _11493_/S vssd1 vssd1 vccd1 vccd1 _11494_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14354__A _14354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16020_ _16020_/A vssd1 vssd1 vccd1 vccd1 _19432_/D sky130_fd_sc_hd__clkbuf_1
X_13232_ _13232_/A vssd1 vssd1 vccd1 vccd1 _18480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ _10548_/A _10443_/X _10323_/A vssd1 vssd1 vccd1 vccd1 _10444_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09448__A _17338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15884__S _15890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ _13163_/A vssd1 vssd1 vccd1 vccd1 _13468_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_10375_ _09918_/A _10374_/X _09826_/A vssd1 vssd1 vccd1 vccd1 _10375_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12114_ _12218_/A vssd1 vssd1 vccd1 vccd1 _12537_/A sky130_fd_sc_hd__buf_2
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13094_ _19929_/Q _19930_/Q _13094_/C vssd1 vssd1 vccd1 vccd1 _13132_/C sky130_fd_sc_hd__and3_1
X_17971_ _17971_/A _17971_/B vssd1 vssd1 vccd1 vccd1 _17971_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output159_A _12472_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19710_ _19718_/CLK _19710_/D vssd1 vssd1 vccd1 vccd1 _19710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16922_ _19727_/Q _16922_/B _16922_/C _16922_/D vssd1 vssd1 vccd1 vccd1 _16923_/D
+ sky130_fd_sc_hd__and4_1
X_12045_ _12045_/A _12045_/B vssd1 vssd1 vccd1 vccd1 _12049_/A sky130_fd_sc_hd__xnor2_1
XFILLER_133_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12602__A _12602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19641_ _19769_/CLK _19641_/D vssd1 vssd1 vccd1 vccd1 _19641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17623__A1 _09345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16853_ _19716_/Q _19715_/Q _16864_/C _16853_/D vssd1 vssd1 vccd1 vccd1 _16868_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15804_ _18462_/Q _13449_/X _15803_/Y _15700_/X vssd1 vssd1 vccd1 vccd1 _15804_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19572_ _19572_/CLK _19572_/D vssd1 vssd1 vccd1 vccd1 _19572_/Q sky130_fd_sc_hd__dfxtp_1
X_16784_ _19699_/Q _16784_/B vssd1 vssd1 vccd1 vccd1 _16790_/C sky130_fd_sc_hd__and2_1
XFILLER_93_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13996_ _18633_/Q _13739_/X _13998_/S vssd1 vssd1 vccd1 vccd1 _13997_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18523_ _19049_/CLK _18523_/D vssd1 vssd1 vccd1 vccd1 _18523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735_ _15735_/A vssd1 vssd1 vccd1 vccd1 _19336_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12947_ _12947_/A vssd1 vssd1 vccd1 vccd1 _12947_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13433__A _15276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18454_ _19952_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15666_ _15661_/X _19324_/Q _15684_/S vssd1 vssd1 vccd1 vccd1 _15667_/A sky130_fd_sc_hd__mux2_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _17052_/A vssd1 vssd1 vccd1 vccd1 _17122_/A sky130_fd_sc_hd__buf_4
XFILLER_61_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17419_/A vssd1 vssd1 vccd1 vccd1 _17549_/A sky130_fd_sc_hd__clkbuf_2
X_14617_ _14617_/A vssd1 vssd1 vccd1 vccd1 _18876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10268__S _10268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18385_ input35/X vssd1 vssd1 vccd1 vccd1 _18385_/Y sky130_fd_sc_hd__clkinv_2
X_11829_ _11820_/Y _11826_/X _11828_/X vssd1 vssd1 vccd1 vccd1 _11829_/X sky130_fd_sc_hd__o21a_1
X_15597_ _15597_/A vssd1 vssd1 vccd1 vccd1 _19292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17336_ _17336_/A _17336_/B vssd1 vssd1 vccd1 vccd1 _17342_/C sky130_fd_sc_hd__nor2_1
XFILLER_81_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14548_ _14559_/A vssd1 vssd1 vccd1 vccd1 _14557_/S sky130_fd_sc_hd__buf_2
XANTENNA__10857__S0 _10777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17267_ _17175_/Y _19858_/Q _17269_/S vssd1 vssd1 vccd1 vccd1 _17268_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16362__A1 _16361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14479_ _14479_/A hold12/X _14479_/C _18198_/B vssd1 vssd1 vccd1 vccd1 _14831_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_174_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19006_ _19486_/CLK _19006_/D vssd1 vssd1 vccd1 vccd1 _19006_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13176__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16218_ _16218_/A vssd1 vssd1 vccd1 vccd1 _19517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17198_ _17242_/B vssd1 vssd1 vccd1 vccd1 _17210_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12923__A1 _18461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17311__A0 _15828_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16149_ _16149_/A vssd1 vssd1 vccd1 vccd1 _19489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10934__B1 _10065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11034__S0 _10914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19908_ _19914_/CLK _19908_/D vssd1 vssd1 vccd1 vccd1 _19908_/Q sky130_fd_sc_hd__dfxtp_4
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_60_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10698__C1 _09603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10162__A1 _19153_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19839_ _19876_/CLK _19839_/D vssd1 vssd1 vccd1 vccd1 _19839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11337__S1 _11179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09523_ _09569_/A vssd1 vssd1 vccd1 vccd1 _09526_/A sky130_fd_sc_hd__buf_2
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13343__A _13343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09454_ _11824_/A _12207_/C vssd1 vssd1 vccd1 vccd1 _11827_/A sky130_fd_sc_hd__or2_2
XFILLER_169_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09385_ _20009_/Q vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14902__A _14902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10160_ _18690_/Q _19185_/Q _10160_/S vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11737__S _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _10817_/A vssd1 vssd1 vccd1 vccd1 _11443_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13850_ _14675_/A vssd1 vssd1 vccd1 vccd1 _13850_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ _19849_/Q _12798_/Y _12799_/Y _19517_/Q _12800_/X vssd1 vssd1 vccd1 vccd1
+ _12801_/X sky130_fd_sc_hd__a221o_1
XFILLER_28_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10993_ _11216_/A _10992_/X _10920_/X vssd1 vssd1 vccd1 vccd1 _10993_/Y sky130_fd_sc_hd__o21ai_1
X_13781_ _13780_/X _18548_/Q _13781_/S vssd1 vssd1 vccd1 vccd1 _13782_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18030__A1 _19915_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15520_ _19258_/Q _15197_/X _15528_/S vssd1 vssd1 vccd1 vccd1 _15521_/A sky130_fd_sc_hd__mux2_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _18453_/Q _13301_/B _13301_/C _13301_/D vssd1 vssd1 vccd1 vccd1 _12732_/X
+ sky130_fd_sc_hd__or4_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15879__S _15879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _15451_/A vssd1 vssd1 vccd1 vccd1 _19227_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12663_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _12663_/Y sky130_fd_sc_hd__nor2_4
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14402_ _18804_/Q _14401_/X _14402_/S vssd1 vssd1 vccd1 vccd1 _14403_/A sky130_fd_sc_hd__mux2_1
X_11614_ _11614_/A vssd1 vssd1 vccd1 vccd1 _18929_/D sky130_fd_sc_hd__clkbuf_1
X_18170_ _19944_/Q _19976_/Q _18170_/S vssd1 vssd1 vccd1 vccd1 _18171_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10839__S0 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15382_ _14586_/X _19197_/Q _15384_/S vssd1 vssd1 vccd1 vccd1 _15383_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12606_/A _12594_/B _12594_/C vssd1 vssd1 vccd1 vccd1 _12596_/C sky130_fd_sc_hd__and3_1
XFILLER_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ _17120_/B _17120_/C _19803_/Q vssd1 vssd1 vccd1 vccd1 _17122_/C sky130_fd_sc_hd__a21oi_1
XFILLER_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14333_ _18778_/Q _13676_/X _14341_/S vssd1 vssd1 vccd1 vccd1 _14334_/A sky130_fd_sc_hd__mux2_1
X_11545_ _11545_/A _11545_/B vssd1 vssd1 vccd1 vccd1 _11545_/X sky130_fd_sc_hd__and2_1
XANTENNA__17541__B1 _17607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13158__B2 _17176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17052_ _17052_/A vssd1 vssd1 vccd1 vccd1 _17089_/A sky130_fd_sc_hd__buf_2
X_14264_ _13806_/X _18748_/Q _14268_/S vssd1 vssd1 vccd1 vccd1 _14265_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11476_ _19482_/Q _19320_/Q _18729_/Q _18499_/Q _10675_/A _09985_/A vssd1 vssd1 vccd1
+ vccd1 _11476_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16003_ _16060_/S vssd1 vssd1 vccd1 vccd1 _16012_/S sky130_fd_sc_hd__buf_2
X_10427_ _19374_/Q _18988_/Q _19438_/Q _18557_/Q _10367_/S _10291_/X vssd1 vssd1 vccd1
+ vccd1 _10428_/B sky130_fd_sc_hd__mux4_1
X_13215_ _13255_/A _13215_/B _13225_/B vssd1 vssd1 vccd1 vccd1 _13215_/X sky130_fd_sc_hd__or3_1
X_14195_ _14195_/A vssd1 vssd1 vccd1 vccd1 _18717_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_183_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10358_ _10490_/A _10357_/X _10323_/X vssd1 vssd1 vccd1 vccd1 _10358_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13146_ _19900_/Q _15701_/B _13430_/S vssd1 vssd1 vccd1 vccd1 _13146_/X sky130_fd_sc_hd__mux2_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15119__S _15127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _18501_/Q _13077_/B vssd1 vssd1 vccd1 vccd1 _13077_/X sky130_fd_sc_hd__and2_1
X_17954_ _17928_/X _17932_/Y _17952_/X _17953_/X vssd1 vssd1 vccd1 vccd1 _17954_/X
+ sky130_fd_sc_hd__o211a_1
X_10289_ _11418_/A _12659_/B vssd1 vssd1 vccd1 vccd1 _11554_/A sky130_fd_sc_hd__or2_1
XFILLER_111_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16905_ _16924_/B _16909_/D _19733_/Q vssd1 vssd1 vccd1 vccd1 _16907_/B sky130_fd_sc_hd__a21oi_1
XFILLER_39_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12028_ _12027_/A _12027_/C hold21/A vssd1 vssd1 vccd1 vccd1 _12029_/D sky130_fd_sc_hd__a21o_1
XFILLER_78_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17885_ _18002_/A _17885_/B _17885_/C _17885_/D vssd1 vssd1 vccd1 vccd1 _17885_/X
+ sky130_fd_sc_hd__or4_1
X_19624_ _19759_/CLK _19624_/D vssd1 vssd1 vccd1 vccd1 _19624_/Q sky130_fd_sc_hd__dfxtp_1
X_16836_ _19712_/Q _16848_/C vssd1 vssd1 vccd1 vccd1 _16838_/A sky130_fd_sc_hd__and2_1
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16280__A0 _19528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16458__B _16458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19555_ _19555_/CLK _19555_/D vssd1 vssd1 vccd1 vccd1 _19555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16767_ _19693_/Q _16765_/B _16766_/Y vssd1 vssd1 vccd1 vccd1 _19693_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14259__A _14281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ _18625_/Q _13706_/X _13983_/S vssd1 vssd1 vccd1 vccd1 _13980_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18506_ _19857_/CLK _18506_/D vssd1 vssd1 vccd1 vccd1 _18506_/Q sky130_fd_sc_hd__dfxtp_1
X_15718_ _13568_/X _15716_/X _15717_/Y _12903_/X _18446_/Q vssd1 vssd1 vccd1 vccd1
+ _15718_/X sky130_fd_sc_hd__a32o_4
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19486_ _19486_/CLK _19486_/D vssd1 vssd1 vccd1 vccd1 _19486_/Q sky130_fd_sc_hd__dfxtp_1
X_16698_ _19781_/Q _19783_/Q _19782_/Q _17056_/A vssd1 vssd1 vccd1 vccd1 _17065_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18437_ _19930_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_1
X_15649_ _14660_/X _19316_/Q _15655_/S vssd1 vssd1 vccd1 vccd1 _15650_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18368_ _18283_/A _12795_/X _14831_/X _18367_/Y vssd1 vssd1 vccd1 vccd1 _18369_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_147_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17319_ _17319_/A _17319_/B vssd1 vssd1 vccd1 vccd1 _17376_/A sky130_fd_sc_hd__and2_1
XANTENNA__16335__A1 _12127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18299_ _18299_/A _18326_/B vssd1 vssd1 vccd1 vccd1 _18299_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11411__A _11411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16413__S _16415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09816__A _10312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15029__S _15033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10135__B2 _10134_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16649__A _16674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18260__A1 _19605_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10230__S1 _09927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16810__A2 _13748_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13085__A0 _19897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13073__A _16219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ _10245_/S vssd1 vssd1 vccd1 vccd1 _10244_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10843__C1 _09602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09437_ _18349_/A _18347_/A vssd1 vssd1 vccd1 vccd1 _11640_/C sky130_fd_sc_hd__or2_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16384__A _16441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09368_ _20016_/Q vssd1 vssd1 vccd1 vccd1 _09389_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09299_ _11634_/B _11678_/A vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__and2b_1
XFILLER_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11330_ _11330_/A _11330_/B vssd1 vssd1 vccd1 vccd1 _11330_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11261_ _11190_/A _11258_/X _11260_/X _10941_/X vssd1 vssd1 vccd1 vccd1 _11261_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10049__S1 _10037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10212_ _10254_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10212_/X sky130_fd_sc_hd__or2_1
XFILLER_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13000_ _13163_/A vssd1 vssd1 vccd1 vccd1 _13553_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17826__A1 _19901_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11192_ _09954_/A _11191_/X _11116_/A vssd1 vssd1 vccd1 vccd1 _11192_/X sky130_fd_sc_hd__a21o_1
XFILLER_133_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10143_ _10143_/A _09896_/Y vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__or2b_1
XFILLER_79_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14951_ _14951_/A vssd1 vssd1 vccd1 vccd1 _19016_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input35_A io_ibus_inst[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _10074_/A vssd1 vssd1 vccd1 vccd1 _10609_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14778__S _14786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__B1 _09609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13682__S _13694_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13902_ _13913_/A vssd1 vssd1 vccd1 vccd1 _13911_/S sky130_fd_sc_hd__buf_2
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11874__A1 _19518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17670_ _17624_/X _17645_/X _17667_/Y _18007_/A _11767_/Y vssd1 vssd1 vccd1 vccd1
+ _17670_/X sky130_fd_sc_hd__a32o_4
X_14882_ _14882_/A vssd1 vssd1 vccd1 vccd1 _18985_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10221__S1 _09927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16262__A0 _12854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16621_ _16631_/A _16627_/C vssd1 vssd1 vccd1 vccd1 _16621_/Y sky130_fd_sc_hd__nor2_1
X_13833_ _13831_/X _18564_/Q _13845_/S vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19340_ _19859_/CLK _19340_/D vssd1 vssd1 vccd1 vccd1 _19340_/Q sky130_fd_sc_hd__dfxtp_1
X_16552_ _19624_/Q _16555_/C _16533_/X vssd1 vssd1 vccd1 vccd1 _16552_/Y sky130_fd_sc_hd__a21oi_1
X_13764_ _14589_/A vssd1 vssd1 vccd1 vccd1 _13764_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _11091_/A vssd1 vssd1 vccd1 vccd1 _10976_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09295__A2 _14148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15503_ _19251_/Q _15279_/X _15511_/S vssd1 vssd1 vccd1 vccd1 _15504_/A sky130_fd_sc_hd__mux2_1
X_19271_ _19559_/CLK _19271_/D vssd1 vssd1 vccd1 vccd1 _19271_/Q sky130_fd_sc_hd__dfxtp_1
X_12715_ _19754_/Q _12692_/X _12710_/X _12714_/X vssd1 vssd1 vccd1 vccd1 _12715_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16483_ _19599_/Q _16477_/X _12371_/Y _12374_/Y _16482_/X vssd1 vssd1 vccd1 vccd1
+ _19599_/D sky130_fd_sc_hd__o221a_1
X_13695_ _13695_/A vssd1 vssd1 vccd1 vccd1 _18526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15402__S _15406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18222_ _18268_/S vssd1 vssd1 vccd1 vccd1 _18231_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15434_ _15434_/A vssd1 vssd1 vccd1 vccd1 _19220_/D sky130_fd_sc_hd__clkbuf_1
X_12646_ _12646_/A vssd1 vssd1 vccd1 vccd1 _12646_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18153_ _16265_/A _19968_/Q _18159_/S vssd1 vssd1 vccd1 vccd1 _18154_/A sky130_fd_sc_hd__mux2_1
X_15365_ _19190_/Q _15289_/X _15367_/S vssd1 vssd1 vccd1 vccd1 _15366_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11485__S0 _10812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12577_ _12618_/A _12577_/B vssd1 vssd1 vccd1 vccd1 _12579_/A sky130_fd_sc_hd__nand2_2
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14018__S _14024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10062__B1 _10000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17104_ _19797_/Q _17104_/B _17104_/C vssd1 vssd1 vccd1 vccd1 _17106_/B sky130_fd_sc_hd__and3_1
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _14316_/A vssd1 vssd1 vccd1 vccd1 _18770_/D sky130_fd_sc_hd__clkbuf_1
X_11528_ _11600_/A _11532_/A _09426_/B vssd1 vssd1 vccd1 vccd1 _11528_/X sky130_fd_sc_hd__o21a_1
X_18084_ _17624_/X _18082_/X _18083_/X _17754_/A _12509_/Y vssd1 vssd1 vccd1 vccd1
+ _18084_/X sky130_fd_sc_hd__a32o_1
X_15296_ _19160_/Q _15295_/X _15299_/S vssd1 vssd1 vccd1 vccd1 _15297_/A sky130_fd_sc_hd__mux2_1
X_17035_ hold20/A _17034_/C _17021_/X vssd1 vssd1 vccd1 vccd1 _17035_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14247_ _14247_/A vssd1 vssd1 vccd1 vccd1 _18740_/D sky130_fd_sc_hd__clkbuf_1
X_11459_ _19385_/Q _18999_/Q _19449_/Q _18568_/Q _10658_/X _10703_/A vssd1 vssd1 vccd1
+ vccd1 _11460_/B sky130_fd_sc_hd__mux4_1
XFILLER_125_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13551__A1 _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__C1 _10949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14178_ _14178_/A vssd1 vssd1 vccd1 vccd1 _18709_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_140_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19258_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _18475_/Q _13128_/X _13196_/S vssd1 vssd1 vccd1 vccd1 _13130_/A sky130_fd_sc_hd__mux2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18986_ _19306_/CLK _18986_/D vssd1 vssd1 vccd1 vccd1 _18986_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _17937_/A _17933_/B vssd1 vssd1 vccd1 vccd1 _17937_/X sky130_fd_sc_hd__or2b_1
XFILLER_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_155_clock clkbuf_opt_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19637_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17868_ _17697_/X _17865_/X _17867_/X vssd1 vssd1 vccd1 vccd1 _17868_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19607_ _19988_/CLK _19607_/D vssd1 vssd1 vccd1 vccd1 _19607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16819_ _19707_/Q _16814_/A _16818_/Y vssd1 vssd1 vccd1 vccd1 _19707_/D sky130_fd_sc_hd__o21a_1
XFILLER_66_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17799_ _17682_/X _17685_/X _17799_/S vssd1 vssd1 vccd1 vccd1 _17799_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11406__A _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19538_ _19542_/CLK _19538_/D vssd1 vssd1 vccd1 vccd1 _19538_/Q sky130_fd_sc_hd__dfxtp_2
X_19469_ _19563_/CLK _19469_/D vssd1 vssd1 vccd1 vccd1 _19469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15820__B _18464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13621__A _15206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09222_ _09191_/B _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09467_/B sky130_fd_sc_hd__and3b_1
XFILLER_167_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11476__S0 _10675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11141__A _11141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11228__S0 _11161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16143__S _16145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_108_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19478_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09546__A _11482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15982__S _15984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10451__S1 _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ _19382_/Q _18996_/Q _19446_/Q _18565_/Q _09984_/X _09985_/X vssd1 vssd1 vccd1
+ vccd1 _09987_/B sky130_fd_sc_hd__mux4_1
XFILLER_153_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15283__A _15283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11400__S0 _10053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10830_ _18772_/Q _19043_/Q _19267_/Q _19011_/Q _10811_/S _09970_/X vssd1 vssd1 vccd1
+ vccd1 _10830_/X sky130_fd_sc_hd__mux4_2
XANTENNA_clkbuf_leaf_131_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _10764_/A _10758_/X _10760_/X vssd1 vssd1 vccd1 vccd1 _10761_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12500_ _19984_/Q _10137_/A _12528_/S vssd1 vssd1 vccd1 vccd1 _12501_/A sky130_fd_sc_hd__mux2_4
X_10692_ _19496_/Q _18908_/Q _18945_/Q _18519_/Q _10690_/X _10691_/X vssd1 vssd1 vccd1
+ vccd1 _10692_/X sky130_fd_sc_hd__mux4_2
X_13480_ _19637_/Q _13204_/X _13479_/X vssd1 vssd1 vccd1 vccd1 _13480_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12431_ _19981_/Q _10144_/A _17464_/S vssd1 vssd1 vccd1 vccd1 _12432_/A sky130_fd_sc_hd__mux2_4
XANTENNA__12033__A1 _17176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10044__B1 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15150_ _15150_/A vssd1 vssd1 vccd1 vccd1 _19106_/D sky130_fd_sc_hd__clkbuf_1
X_12362_ _12362_/A vssd1 vssd1 vccd1 vccd1 _12362_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_154_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14101_ _18677_/Q _13655_/X _14109_/S vssd1 vssd1 vccd1 vccd1 _14102_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11313_ _10949_/X _11304_/Y _11308_/Y _11312_/Y _09599_/A vssd1 vssd1 vccd1 vccd1
+ _11313_/X sky130_fd_sc_hd__o311a_2
XANTENNA__15458__A _15515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12293_ _19835_/Q vssd1 vssd1 vccd1 vccd1 _17205_/A sky130_fd_sc_hd__clkbuf_2
X_15081_ _14602_/X _19074_/Q _15083_/S vssd1 vssd1 vccd1 vccd1 _15082_/A sky130_fd_sc_hd__mux2_1
X_14032_ _14032_/A vssd1 vssd1 vccd1 vccd1 _18647_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09456__A input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ _10875_/X _11239_/X _11241_/X _11243_/X _11012_/A vssd1 vssd1 vccd1 vccd1
+ _11244_/X sky130_fd_sc_hd__a221o_2
XFILLER_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_56_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ _11183_/A _11171_/X _11174_/X vssd1 vssd1 vccd1 vccd1 _11175_/Y sky130_fd_sc_hd__o21ai_1
X_18840_ _19074_/CLK _18840_/D vssd1 vssd1 vccd1 vccd1 _18840_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10442__S1 _10326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19571_/CLK sky130_fd_sc_hd__clkbuf_16
X_10126_ _19511_/Q _18923_/Q _18960_/Q _18534_/Q _11449_/S _10718_/A vssd1 vssd1 vccd1
+ vccd1 _10126_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18771_ _19493_/CLK _18771_/D vssd1 vssd1 vccd1 vccd1 _18771_/Q sky130_fd_sc_hd__dfxtp_1
X_15983_ _15983_/A vssd1 vssd1 vccd1 vccd1 _19416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17722_ _17722_/A vssd1 vssd1 vccd1 vccd1 _17723_/A sky130_fd_sc_hd__clkbuf_2
X_10057_ _10052_/X _10055_/X _10056_/X vssd1 vssd1 vccd1 vccd1 _10057_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14934_ _14934_/A vssd1 vssd1 vccd1 vccd1 _19008_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17653_ _17455_/X _17466_/X _17802_/D vssd1 vssd1 vccd1 vccd1 _17654_/B sky130_fd_sc_hd__mux2_1
X_14865_ _14602_/X _18978_/Q _14867_/S vssd1 vssd1 vccd1 vccd1 _14866_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_87_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19498_/CLK sky130_fd_sc_hd__clkbuf_16
X_16604_ _19641_/Q _16601_/B _16603_/Y vssd1 vssd1 vccd1 vccd1 _19641_/D sky130_fd_sc_hd__o21a_1
X_13816_ _13832_/A vssd1 vssd1 vccd1 vccd1 _13829_/S sky130_fd_sc_hd__buf_2
XANTENNA__10130__A _10846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17584_ _17582_/X _17583_/X _17686_/S vssd1 vssd1 vccd1 vccd1 _17584_/X sky130_fd_sc_hd__mux2_1
X_14796_ _14796_/A vssd1 vssd1 vccd1 vccd1 _18951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ _19594_/CLK _19323_/D vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
X_16535_ _16538_/B _16538_/C _16534_/Y vssd1 vssd1 vccd1 vccd1 _19618_/D sky130_fd_sc_hd__o21a_1
X_13747_ _14074_/A vssd1 vssd1 vccd1 vccd1 _18299_/A sky130_fd_sc_hd__inv_2
X_10959_ _11016_/A _10956_/X _10958_/X _10949_/X vssd1 vssd1 vccd1 vccd1 _10959_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14537__A _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18009__A _18009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19254_ _19416_/CLK _19254_/D vssd1 vssd1 vccd1 vccd1 _19254_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_10_clock _19998_/CLK vssd1 vssd1 vccd1 vccd1 _20000_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11480__C1 _09601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16466_ _16466_/A vssd1 vssd1 vccd1 vccd1 _19588_/D sky130_fd_sc_hd__clkbuf_1
X_13678_ _18522_/Q _13676_/X _13694_/S vssd1 vssd1 vccd1 vccd1 _13679_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_opt_3_0_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18205_ _19959_/Q _19580_/Q _18209_/S vssd1 vssd1 vccd1 vccd1 _18206_/A sky130_fd_sc_hd__mux2_1
X_15417_ _14637_/X _19213_/Q _15417_/S vssd1 vssd1 vccd1 vccd1 _15418_/A sky130_fd_sc_hd__mux2_1
X_19185_ _19411_/CLK _19185_/D vssd1 vssd1 vccd1 vccd1 _19185_/Q sky130_fd_sc_hd__dfxtp_1
X_12629_ _19609_/Q _12537_/X _12625_/Y _12628_/Y vssd1 vssd1 vccd1 vccd1 _12629_/X
+ sky130_fd_sc_hd__o22a_4
X_16397_ _16397_/A vssd1 vssd1 vccd1 vccd1 _19556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18136_ _16219_/B _19961_/Q _18136_/S vssd1 vssd1 vccd1 vccd1 _18137_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15348_ _19182_/Q _15263_/X _15356_/S vssd1 vssd1 vccd1 vccd1 _15349_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_25_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19406_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16471__B _16471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18067_ _18065_/Y _18066_/X _18089_/S vssd1 vssd1 vccd1 vccd1 _18067_/X sky130_fd_sc_hd__mux2_1
X_15279_ _15279_/A vssd1 vssd1 vccd1 vccd1 _15279_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17018_ _17066_/A _17025_/C vssd1 vssd1 vccd1 vccd1 _17018_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09840_ _09918_/A vssd1 vssd1 vccd1 vccd1 _10147_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09771_ _10205_/A _09771_/B _09771_/C vssd1 vssd1 vccd1 vccd1 _09771_/X sky130_fd_sc_hd__or3_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _19671_/CLK _18969_/D vssd1 vssd1 vccd1 vccd1 _18969_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18829__D _18829_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16927__A _16946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10040__A _10040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09205_ _12601_/A vssd1 vssd1 vccd1 vccd1 _12610_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__13212__A0 _19903_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17758__A _18019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14881__S _14889_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12015__B2 _20050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10577__A1 _09615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10577__B2 _19908_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13515__B2 _19543_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_clock clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09969_ _10074_/A vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12980_ _17861_/A vssd1 vssd1 vccd1 vccd1 _12980_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16217__A0 _19517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10869__B _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11931_ _19963_/Q _11352_/A _11966_/A vssd1 vssd1 vccd1 vccd1 _11969_/A sky130_fd_sc_hd__mux2_4
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11046__A _11046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14650_/A vssd1 vssd1 vccd1 vccd1 _14650_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _11815_/A _11815_/B _11813_/A vssd1 vssd1 vccd1 vccd1 _11933_/B sky130_fd_sc_hd__a21o_2
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _15702_/A _18468_/Q vssd1 vssd1 vccd1 vccd1 _13601_/Y sky130_fd_sc_hd__nand2_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ _10813_/A _10813_/B vssd1 vssd1 vccd1 vccd1 _10813_/X sky130_fd_sc_hd__and2_1
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _14580_/X _18865_/Q _14590_/S vssd1 vssd1 vccd1 vccd1 _14582_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16048__S _16056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _12155_/B vssd1 vssd1 vccd1 vccd1 _12584_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__10885__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16320_ _16320_/A vssd1 vssd1 vccd1 vccd1 _19535_/D sky130_fd_sc_hd__clkbuf_1
X_13532_ hold20/A _12804_/Y _12799_/Y _19544_/Q _13531_/X vssd1 vssd1 vccd1 vccd1
+ _13532_/X sky130_fd_sc_hd__a221o_1
X_10744_ _19463_/Q _19301_/Q _18710_/Q _18480_/Q _10614_/X _10682_/X vssd1 vssd1 vccd1
+ vccd1 _10744_/X sky130_fd_sc_hd__mux4_2
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14076__B _16809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16251_ _15718_/X _16250_/Y _16262_/S vssd1 vssd1 vccd1 vccd1 _16251_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14791__S _14797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13463_ _19350_/Q _13245_/X _13099_/X _19540_/Q _13462_/X vssd1 vssd1 vccd1 vccd1
+ _13463_/X sky130_fd_sc_hd__a221o_1
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10675_ _10675_/A vssd1 vssd1 vccd1 vccd1 _10675_/X sky130_fd_sc_hd__buf_4
X_15202_ _15202_/A vssd1 vssd1 vccd1 vccd1 _19130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12414_ _12414_/A vssd1 vssd1 vccd1 vccd1 _12414_/Y sky130_fd_sc_hd__inv_6
X_16182_ _16182_/A vssd1 vssd1 vccd1 vccd1 _19504_/D sky130_fd_sc_hd__clkbuf_1
X_13394_ _18490_/Q _13393_/X _13434_/S vssd1 vssd1 vccd1 vccd1 _13395_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15133_ _19098_/Q vssd1 vssd1 vccd1 vccd1 _15134_/A sky130_fd_sc_hd__clkbuf_1
X_12345_ _17210_/A _12373_/C _12855_/A vssd1 vssd1 vccd1 vccd1 _12345_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10663__S1 _10014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__S _10824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15064_ _14574_/X _19066_/Q _15072_/S vssd1 vssd1 vccd1 vccd1 _15065_/A sky130_fd_sc_hd__mux2_1
X_19941_ _19981_/CLK _19941_/D vssd1 vssd1 vccd1 vccd1 _19941_/Q sky130_fd_sc_hd__dfxtp_1
X_12276_ _19975_/Q _10459_/A _12573_/S vssd1 vssd1 vccd1 vccd1 _17452_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14015_ _14072_/S vssd1 vssd1 vccd1 vccd1 _14024_/S sky130_fd_sc_hd__buf_2
XFILLER_141_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11227_ _18574_/Q _18835_/Q _18734_/Q _19069_/Q _11085_/A _09659_/A vssd1 vssd1 vccd1
+ vccd1 _11227_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10125__A _10846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19872_ _19873_/CLK _19872_/D vssd1 vssd1 vccd1 vccd1 _19872_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16456__B1 _16455_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18823_ _19416_/CLK _18823_/D vssd1 vssd1 vccd1 vccd1 _18823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11158_ _09746_/A _11144_/X _11156_/X _09753_/A _11157_/Y vssd1 vssd1 vccd1 vccd1
+ _12636_/B sky130_fd_sc_hd__o32a_2
XANTENNA__15127__S _15127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10109_ _18694_/Q _19189_/Q _11495_/S vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__mux2_1
X_18754_ _19476_/CLK _18754_/D vssd1 vssd1 vccd1 vccd1 _18754_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14031__S _14035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15966_ _15966_/A vssd1 vssd1 vccd1 vccd1 _19408_/D sky130_fd_sc_hd__clkbuf_1
X_11089_ _10899_/A _11088_/X _10988_/X vssd1 vssd1 vccd1 vccd1 _11089_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10179__S0 _09653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14917_ _18299_/A _14917_/B _15373_/A _14917_/D vssd1 vssd1 vccd1 vccd1 _14974_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17705_ _17705_/A vssd1 vssd1 vccd1 vccd1 _17705_/X sky130_fd_sc_hd__buf_2
XANTENNA__12493__A1 _19843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15897_ _13412_/X _19378_/Q _15901_/S vssd1 vssd1 vccd1 vccd1 _15898_/A sky130_fd_sc_hd__mux2_1
X_18685_ _19406_/CLK _18685_/D vssd1 vssd1 vccd1 vccd1 _18685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13870__S _13878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17636_ _17760_/S vssd1 vssd1 vccd1 vccd1 _17803_/S sky130_fd_sc_hd__clkbuf_2
X_14848_ _14574_/X _18970_/Q _14856_/S vssd1 vssd1 vccd1 vccd1 _14849_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17567_ _17563_/X _17566_/X _17802_/B vssd1 vssd1 vccd1 vccd1 _17567_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14779_ _14779_/A vssd1 vssd1 vccd1 vccd1 _18943_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19306_ _19306_/CLK _19306_/D vssd1 vssd1 vccd1 vccd1 _19306_/Q sky130_fd_sc_hd__dfxtp_1
X_16518_ _19613_/Q _16518_/B _16518_/C vssd1 vssd1 vccd1 vccd1 _16519_/C sky130_fd_sc_hd__and3_1
XANTENNA__11453__C1 _10757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17498_ _12480_/A _17749_/B _17506_/S vssd1 vssd1 vccd1 vccd1 _17498_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19237_ _19402_/CLK _19237_/D vssd1 vssd1 vccd1 vccd1 _19237_/Q sky130_fd_sc_hd__dfxtp_1
X_16449_ _16487_/A vssd1 vssd1 vccd1 vccd1 _16449_/X sky130_fd_sc_hd__buf_2
XFILLER_158_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16482__A _16939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19168_ _19395_/CLK _19168_/D vssd1 vssd1 vccd1 vccd1 _19168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18119_ _17815_/A _12614_/B _17998_/A _18118_/X vssd1 vssd1 vccd1 vccd1 _18119_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19099_ _19734_/CLK _19099_/D vssd1 vssd1 vccd1 vccd1 _19099_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10654__S1 _10645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12234__B _12234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10406__S1 _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10035__A _10751_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20012_ _20020_/CLK _20012_/D vssd1 vssd1 vccd1 vccd1 _20012_/Q sky130_fd_sc_hd__dfxtp_1
X_09823_ _18788_/Q _19059_/Q _19283_/Q _19027_/Q _09812_/X _09822_/X vssd1 vssd1 vccd1
+ vccd1 _09823_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09754_ _10065_/A vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09685_ _10283_/A vssd1 vssd1 vccd1 vccd1 _10188_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14876__S _14878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16657__A _16674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10909__S _10909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11444__C1 _09577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10798__B2 _10063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10460_ _10460_/A _10460_/B vssd1 vssd1 vccd1 vccd1 _11560_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10391_ _10391_/A vssd1 vssd1 vccd1 vccd1 _10391_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14116__S _14120_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12425__A _18333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13020__S _13090_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12130_ _17187_/A _12157_/C vssd1 vssd1 vccd1 vccd1 _12130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17935__B _17937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13955__S _13961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ _19524_/Q _11915_/A _12032_/A vssd1 vssd1 vccd1 vccd1 _12061_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14640__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11012_ _11012_/A _11012_/B _11012_/C vssd1 vssd1 vccd1 vccd1 _11012_/X sky130_fd_sc_hd__or3_2
XFILLER_1_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15820_ _15837_/A _18464_/Q vssd1 vssd1 vccd1 vccd1 _15820_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15661__A1 _13572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _18452_/Q _12853_/X _15750_/X vssd1 vssd1 vccd1 vccd1 _17194_/A sky130_fd_sc_hd__a21oi_4
XFILLER_46_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12963_ _18452_/Q _12959_/X _11411_/A _12962_/X vssd1 vssd1 vccd1 vccd1 _18452_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14786__S _14786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13690__S _13694_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _18905_/Q _14401_/X _14702_/S vssd1 vssd1 vccd1 vccd1 _14703_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _19726_/CLK _18470_/D vssd1 vssd1 vccd1 vccd1 _18470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11914_ _12366_/A _11907_/X _11913_/X _11871_/X vssd1 vssd1 vccd1 vccd1 _11914_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _15814_/A _17160_/A vssd1 vssd1 vccd1 vccd1 _16222_/A sky130_fd_sc_hd__nor2_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _19347_/Q _12802_/A _12704_/A _19537_/Q _12893_/X vssd1 vssd1 vccd1 vccd1
+ _12894_/X sky130_fd_sc_hd__a221o_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17421_/A vssd1 vssd1 vccd1 vccd1 _17749_/B sky130_fd_sc_hd__clkbuf_2
X_14633_ _14633_/A vssd1 vssd1 vccd1 vccd1 _18881_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12227__A1 _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _11958_/B _19820_/Q vssd1 vssd1 vccd1 vccd1 _11845_/X sky130_fd_sc_hd__and2b_1
XFILLER_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output104_A _09209_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _17352_/A vssd1 vssd1 vccd1 vccd1 _19885_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14564_ _13838_/X _18859_/Q _14568_/S vssd1 vssd1 vccd1 vccd1 _14565_/A sky130_fd_sc_hd__mux2_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11776_ _11776_/A vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12319__B _12319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16303_ _16303_/A vssd1 vssd1 vccd1 vccd1 _16303_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13515_ _19353_/Q _13245_/X _13099_/X _19543_/Q _13514_/X vssd1 vssd1 vccd1 vccd1
+ _13515_/X sky130_fd_sc_hd__a221o_1
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17398__A _17507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17283_ _17194_/Y _19865_/Q _17291_/S vssd1 vssd1 vccd1 vccd1 _17284_/A sky130_fd_sc_hd__mux2_1
X_10727_ _10727_/A _12648_/A vssd1 vssd1 vccd1 vccd1 _10728_/B sky130_fd_sc_hd__or2_1
XFILLER_159_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14495_ input49/X vssd1 vssd1 vccd1 vccd1 _14495_/Y sky130_fd_sc_hd__inv_2
X_19022_ _19503_/CLK _19022_/D vssd1 vssd1 vccd1 vccd1 _19022_/Q sky130_fd_sc_hd__dfxtp_1
X_16234_ _16239_/B _16233_/Y _12444_/X vssd1 vssd1 vccd1 vccd1 _16235_/B sky130_fd_sc_hd__a21oi_2
XFILLER_146_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13446_ _19763_/Q _12840_/X _13445_/X _12846_/X vssd1 vssd1 vccd1 vccd1 _13446_/X
+ sky130_fd_sc_hd__a211o_1
X_10658_ _10849_/S vssd1 vssd1 vccd1 vccd1 _10658_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_139_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16165_ _19497_/Q _14618_/A _16167_/S vssd1 vssd1 vccd1 vccd1 _16166_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13377_ _13454_/A vssd1 vssd1 vccd1 vccd1 _13434_/S sky130_fd_sc_hd__buf_2
XFILLER_155_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10589_ _18682_/Q _19177_/Q _10589_/S vssd1 vssd1 vccd1 vccd1 _10590_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15116_ _14653_/X _19090_/Q _15116_/S vssd1 vssd1 vccd1 vccd1 _15117_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12328_ _12328_/A vssd1 vssd1 vccd1 vccd1 _18001_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12950__A2 _12946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16096_ _16096_/A vssd1 vssd1 vccd1 vccd1 _19466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13865__S _13867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10961__B2 _19900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15646__A _15646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15047_ _19059_/Q _14452_/X _15055_/S vssd1 vssd1 vccd1 vccd1 _15048_/A sky130_fd_sc_hd__mux2_1
X_19924_ _19978_/CLK _19924_/D vssd1 vssd1 vccd1 vccd1 _19924_/Q sky130_fd_sc_hd__dfxtp_4
X_12259_ _12259_/A _12259_/B vssd1 vssd1 vccd1 vccd1 _12260_/A sky130_fd_sc_hd__xnor2_4
XFILLER_123_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09644__A _10909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19855_ _19859_/CLK _19855_/D vssd1 vssd1 vccd1 vccd1 _19855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10713__A1 _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18806_ _19369_/CLK _18806_/D vssd1 vssd1 vccd1 vccd1 _18806_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17861__A _17861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19786_ _19805_/CLK _19786_/D vssd1 vssd1 vccd1 vccd1 _19786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16998_ _19757_/Q vssd1 vssd1 vccd1 vccd1 _17005_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18737_ _19200_/CLK _18737_/D vssd1 vssd1 vccd1 vccd1 _18737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15949_ _19401_/Q _15241_/X _15951_/S vssd1 vssd1 vccd1 vccd1 _15950_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14696__S _14702_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16477__A _16487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09470_ _09470_/A vssd1 vssd1 vccd1 vccd1 _10875_/A sky130_fd_sc_hd__clkbuf_2
X_18668_ _19258_/CLK _18668_/D vssd1 vssd1 vccd1 vccd1 _18668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17619_ _17619_/A vssd1 vssd1 vccd1 vccd1 _17619_/X sky130_fd_sc_hd__clkbuf_2
X_18599_ _19574_/CLK _18599_/D vssd1 vssd1 vccd1 vccd1 _18599_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_178_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17157__A1 _13591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18106__B1 _18105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16668__B1 _16667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09806_ _11537_/A _12667_/B vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__and2_1
XFILLER_75_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09737_ _09737_/A vssd1 vssd1 vccd1 vccd1 _09738_/A sky130_fd_sc_hd__buf_2
XFILLER_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09668_ _09929_/A vssd1 vssd1 vccd1 vccd1 _09927_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09599_/A vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _12595_/B _09266_/X _09304_/A vssd1 vssd1 vccd1 vccd1 _11673_/C sky130_fd_sc_hd__a21oi_1
XFILLER_24_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ _11565_/A _11568_/A _11565_/C _10556_/A vssd1 vssd1 vccd1 vccd1 _11561_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ _13371_/A vssd1 vssd1 vccd1 vccd1 _13534_/S sky130_fd_sc_hd__clkbuf_2
X_10512_ _10294_/A _10511_/X _10296_/A vssd1 vssd1 vccd1 vccd1 _10512_/X sky130_fd_sc_hd__a21o_1
X_14280_ _14280_/A vssd1 vssd1 vccd1 vccd1 _18755_/D sky130_fd_sc_hd__clkbuf_1
X_11492_ _09612_/A _11480_/X _11491_/X _09996_/A _19923_/Q vssd1 vssd1 vccd1 vccd1
+ _11520_/A sky130_fd_sc_hd__a32o_4
XFILLER_155_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ _18480_/Q _13230_/X _13278_/S vssd1 vssd1 vccd1 vccd1 _13232_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10443_ _18781_/Q _19052_/Q _19276_/Q _19020_/Q _10390_/S _10333_/A vssd1 vssd1 vccd1
+ vccd1 _10443_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09448__B _18328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12155__A _19527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16659__B1 _16624_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input65_A io_ibus_inst[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13162_ _19650_/Q _12887_/X _12889_/X _19782_/Q vssd1 vssd1 vccd1 vccd1 _15709_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10374_ _18782_/Q _19053_/Q _19277_/Q _19021_/Q _10416_/S _09520_/A vssd1 vssd1 vccd1
+ vccd1 _10374_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12113_ _19590_/Q vssd1 vssd1 vccd1 vccd1 _12119_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17970_ _10506_/Y _17861_/X _17969_/X vssd1 vssd1 vccd1 vccd1 _19910_/D sky130_fd_sc_hd__a21oi_1
X_13093_ _16219_/B _13094_/C _16232_/A vssd1 vssd1 vccd1 vccd1 _13095_/A sky130_fd_sc_hd__a21oi_1
XFILLER_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16921_ _19724_/Q _16921_/B _16921_/C _16921_/D vssd1 vssd1 vccd1 vccd1 _16922_/D
+ sky130_fd_sc_hd__and4_1
X_12044_ _12137_/A _12044_/B vssd1 vssd1 vccd1 vccd1 _12045_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11043__S1 _10974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19640_ _19769_/CLK _19640_/D vssd1 vssd1 vccd1 vccd1 _19640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
X_16852_ _16864_/A _16857_/D _16851_/Y vssd1 vssd1 vccd1 vccd1 _19716_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17623__A2 _17558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15803_ _15811_/A _18462_/Q vssd1 vssd1 vccd1 vccd1 _15803_/Y sky130_fd_sc_hd__nand2_1
X_19571_ _19571_/CLK _19571_/D vssd1 vssd1 vccd1 vccd1 _19571_/Q sky130_fd_sc_hd__dfxtp_1
X_16783_ _16783_/A vssd1 vssd1 vccd1 vccd1 _16818_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12448__A1 _19602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13995_ _13995_/A vssd1 vssd1 vccd1 vccd1 _18632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18522_ _19049_/CLK _18522_/D vssd1 vssd1 vccd1 vccd1 _18522_/Q sky130_fd_sc_hd__dfxtp_1
X_15734_ _15733_/X _19336_/Q _15747_/S vssd1 vssd1 vccd1 vccd1 _15735_/A sky130_fd_sc_hd__mux2_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12946_ _12951_/A vssd1 vssd1 vccd1 vccd1 _12946_/X sky130_fd_sc_hd__clkbuf_8
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _15844_/S vssd1 vssd1 vccd1 vccd1 _15684_/S sky130_fd_sc_hd__clkbuf_2
X_18453_ _19952_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _12884_/A vssd1 vssd1 vccd1 vccd1 _17052_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14616_ _14615_/X _18876_/Q _14622_/S vssd1 vssd1 vccd1 vccd1 _14617_/A sky130_fd_sc_hd__mux2_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17404_ _12617_/A _12620_/A _12620_/B _17403_/X vssd1 vssd1 vccd1 vccd1 _17554_/A
+ sky130_fd_sc_hd__a31o_1
X_11828_ _19517_/Q _11915_/A _11778_/A vssd1 vssd1 vccd1 vccd1 _11828_/X sky130_fd_sc_hd__o21a_1
X_18384_ _18396_/A _18384_/B vssd1 vssd1 vccd1 vccd1 _20030_/D sky130_fd_sc_hd__nor2_1
XANTENNA__17139__A1 _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15596_ _14583_/X _19292_/Q _15600_/S vssd1 vssd1 vccd1 vccd1 _15597_/A sky130_fd_sc_hd__mux2_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17335_ _17395_/A _17335_/B _17335_/C _11895_/C vssd1 vssd1 vccd1 vccd1 _17336_/B
+ sky130_fd_sc_hd__or4b_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14547_ _14547_/A vssd1 vssd1 vccd1 vccd1 _18851_/D sky130_fd_sc_hd__clkbuf_1
X_11759_ _11759_/A _17675_/S vssd1 vssd1 vccd1 vccd1 _11762_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10857__S1 _10010_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09639__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17266_ _17266_/A vssd1 vssd1 vccd1 vccd1 _19857_/D sky130_fd_sc_hd__clkbuf_1
X_14478_ _19323_/D _14478_/B vssd1 vssd1 vccd1 vccd1 _18198_/B sky130_fd_sc_hd__or2_1
XFILLER_174_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19005_ _19487_/CLK _19005_/D vssd1 vssd1 vccd1 vccd1 _19005_/Q sky130_fd_sc_hd__dfxtp_1
X_16217_ _19517_/Q _16216_/X _16223_/S vssd1 vssd1 vccd1 vccd1 _16218_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13429_ _13428_/A _13438_/C _13038_/A vssd1 vssd1 vccd1 vccd1 _13429_/X sky130_fd_sc_hd__o21a_1
XFILLER_162_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17197_ _17197_/A vssd1 vssd1 vccd1 vccd1 _17197_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12923__A2 _12921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16148_ _19489_/Q _14592_/A _16156_/S vssd1 vssd1 vccd1 vccd1 _16149_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10934__A1 _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079_ _16079_/A vssd1 vssd1 vccd1 vccd1 _19458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19907_ _19986_/CLK _19907_/D vssd1 vssd1 vccd1 vccd1 _19907_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11034__S1 _11225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19838_ _19873_/CLK _19838_/D vssd1 vssd1 vccd1 vccd1 _19838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10793__S0 _10849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 io_dbus_rdata[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_8
XFILLER_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19769_ _19769_/CLK _19769_/D vssd1 vssd1 vccd1 vccd1 _19769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09522_ _09809_/A vssd1 vssd1 vccd1 vccd1 _09569_/A sky130_fd_sc_hd__buf_2
XANTENNA__13100__A2 _12992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09453_ _12320_/A _09453_/B _09452_/X vssd1 vssd1 vccd1 vccd1 _12207_/C sky130_fd_sc_hd__or3b_2
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09384_ _09394_/A _13136_/B _18326_/A vssd1 vssd1 vccd1 vccd1 _12693_/C sky130_fd_sc_hd__and3b_1
XFILLER_33_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09549__A _10294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13167__A2 _15709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10386__C1 _09605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15286__A _15286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12703__A _12756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10090_ _11491_/A _10090_/B _10090_/C vssd1 vssd1 vccd1 vccd1 _10090_/X sky130_fd_sc_hd__or3_2
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11319__A _11319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10784__S0 _10751_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16813__B1 _18365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__B2 _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12800_ _19806_/Q _12893_/B vssd1 vssd1 vccd1 vccd1 _12800_/X sky130_fd_sc_hd__and2_1
XFILLER_90_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13780_ _14605_/A vssd1 vssd1 vccd1 vccd1 _13780_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17369__A1 _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10992_ _18642_/Q _19233_/Q _19395_/Q _18610_/Q _10903_/A _10974_/X vssd1 vssd1 vccd1
+ vccd1 _10992_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17369__B2 _19890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _16653_/B _12727_/X _12729_/X _17087_/B vssd1 vssd1 vccd1 vccd1 _13301_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10369__S _10465_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15450_ _19227_/Q _15203_/X _15456_/S vssd1 vssd1 vccd1 vccd1 _15451_/A sky130_fd_sc_hd__mux2_1
X_12662_ _12663_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _12662_/Y sky130_fd_sc_hd__nor2_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14401_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11607_/X _11665_/B _11657_/S vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__mux2_1
X_15381_ _15381_/A vssd1 vssd1 vccd1 vccd1 _19196_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16056__S _16056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10839__S1 _09970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ _12593_/A vssd1 vssd1 vccd1 vccd1 _12593_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__10893__A _11114_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17120_ _19803_/Q _17120_/B _17120_/C vssd1 vssd1 vccd1 vccd1 _17122_/B sky130_fd_sc_hd__and3_1
X_14332_ _14354_/A vssd1 vssd1 vccd1 vccd1 _14341_/S sky130_fd_sc_hd__buf_2
X_11544_ _11544_/A _11544_/B _11544_/C vssd1 vssd1 vccd1 vccd1 _11545_/B sky130_fd_sc_hd__nand3_1
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15895__S _15901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17051_ _17053_/B _17053_/C _17050_/Y vssd1 vssd1 vccd1 vccd1 _19778_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17339__D_N _18328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14263_ _14263_/A vssd1 vssd1 vccd1 vccd1 _18747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11475_ _11475_/A _11475_/B vssd1 vssd1 vccd1 vccd1 _11475_/X sky130_fd_sc_hd__or2_1
XFILLER_143_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11169__A1 _11164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16002_ _16002_/A vssd1 vssd1 vccd1 vccd1 _19424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13214_ _19934_/Q _19935_/Q _13214_/C vssd1 vssd1 vccd1 vccd1 _13225_/B sky130_fd_sc_hd__and3_1
X_10426_ _10426_/A _10426_/B vssd1 vssd1 vccd1 vccd1 _10426_/X sky130_fd_sc_hd__or2_1
XANTENNA__12905__A2 _17220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14194_ _13809_/X _18717_/Q _14196_/S vssd1 vssd1 vccd1 vccd1 _14195_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_126_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13709__A _15273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13145_ _16627_/A _12752_/X _12753_/X _17062_/A _13144_/X vssd1 vssd1 vccd1 vccd1
+ _15701_/B sky130_fd_sc_hd__a221o_1
X_10357_ _18655_/Q _19246_/Q _19408_/Q _18623_/Q _10337_/X _10326_/X vssd1 vssd1 vccd1
+ vccd1 _10357_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14304__S _14308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _19742_/Q vssd1 vssd1 vccd1 vccd1 _16958_/B sky130_fd_sc_hd__clkbuf_2
X_17953_ _17953_/A vssd1 vssd1 vccd1 vccd1 _17953_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10288_ _09750_/A _10277_/X _10286_/X _09757_/A _10287_/Y vssd1 vssd1 vccd1 vccd1
+ _12659_/B sky130_fd_sc_hd__o32a_4
XANTENNA__12332__B _17985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16904_ _16924_/B _16909_/D _16903_/X vssd1 vssd1 vccd1 vccd1 _19732_/D sky130_fd_sc_hd__o21ba_1
X_12027_ _12027_/A hold21/A _12027_/C vssd1 vssd1 vccd1 vccd1 _12086_/C sky130_fd_sc_hd__and3_1
XFILLER_39_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17884_ _17884_/A _17884_/B vssd1 vssd1 vccd1 vccd1 _17885_/D sky130_fd_sc_hd__nor2_1
XFILLER_120_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19623_ _19759_/CLK _19623_/D vssd1 vssd1 vccd1 vccd1 _19623_/Q sky130_fd_sc_hd__dfxtp_1
X_16835_ _16848_/C _16835_/B vssd1 vssd1 vccd1 vccd1 _19711_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19554_ _19555_/CLK _19554_/D vssd1 vssd1 vccd1 vccd1 _19554_/Q sky130_fd_sc_hd__dfxtp_1
X_13978_ _13978_/A vssd1 vssd1 vccd1 vccd1 _18624_/D sky130_fd_sc_hd__clkbuf_1
X_16766_ _16775_/A _16772_/C vssd1 vssd1 vccd1 vccd1 _16766_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18505_ _19745_/CLK _18505_/D vssd1 vssd1 vccd1 vccd1 _18505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15717_ _15737_/A _18446_/Q vssd1 vssd1 vccd1 vccd1 _15717_/Y sky130_fd_sc_hd__nand2_1
X_12929_ _18138_/A vssd1 vssd1 vccd1 vccd1 _18127_/A sky130_fd_sc_hd__clkbuf_4
X_19485_ _19485_/CLK _19485_/D vssd1 vssd1 vccd1 vccd1 _19485_/Q sky130_fd_sc_hd__dfxtp_1
X_16697_ _19779_/Q _19778_/Q _19780_/Q _17047_/A vssd1 vssd1 vccd1 vccd1 _17056_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_34_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18436_ _19892_/CLK input70/X vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_1
X_15648_ _15648_/A vssd1 vssd1 vccd1 vccd1 _19315_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17780__A1 _19899_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15579_ _19285_/Q _15286_/X _15583_/S vssd1 vssd1 vccd1 vccd1 _15580_/A sky130_fd_sc_hd__mux2_1
X_18367_ input61/X vssd1 vssd1 vccd1 vccd1 _18367_/Y sky130_fd_sc_hd__inv_8
XFILLER_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17318_ _17318_/A vssd1 vssd1 vccd1 vccd1 _19881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16335__A2 _15799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18298_ _20031_/Q _18291_/X _18297_/Y _18289_/X vssd1 vssd1 vccd1 vccd1 _19999_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11411__B _12651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17249_ _17317_/S vssd1 vssd1 vccd1 vccd1 _17258_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17296__A0 _15784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14214__S _14218_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12523__A _18343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10978__A _10978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ _09505_/A vssd1 vssd1 vccd1 vccd1 _10245_/S sky130_fd_sc_hd__buf_4
XFILLER_65_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16665__A _16674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ _20051_/Q vssd1 vssd1 vccd1 vccd1 _18347_/A sky130_fd_sc_hd__buf_2
XFILLER_53_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _16808_/A _16808_/B _20018_/Q _20017_/Q vssd1 vssd1 vccd1 vccd1 _12700_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_123_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09298_ _09298_/A vssd1 vssd1 vccd1 vccd1 _17394_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ _11260_/A _11260_/B vssd1 vssd1 vccd1 vccd1 _11260_/X sky130_fd_sc_hd__and2_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17287__A0 _12772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ _19474_/Q _19312_/Q _18721_/Q _18491_/Q _10195_/S _09899_/X vssd1 vssd1 vccd1
+ vccd1 _10212_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09764__A1 _10161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11191_ _18797_/Q _19132_/Q _11191_/S vssd1 vssd1 vccd1 vccd1 _11191_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10142_ _11541_/A _11424_/B _10141_/Y _11544_/B vssd1 vssd1 vccd1 vccd1 _11536_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14950_ _19016_/Q _14417_/X _14950_/S vssd1 vssd1 vccd1 vccd1 _14951_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10073_ _11481_/S vssd1 vssd1 vccd1 vccd1 _10073_/X sky130_fd_sc_hd__buf_4
XANTENNA__11323__A1 _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13901_ _13901_/A vssd1 vssd1 vccd1 vccd1 _18590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14881_ _14624_/X _18985_/Q _14889_/S vssd1 vssd1 vccd1 vccd1 _14882_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input28_A io_dbus_rdata[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11483__S _11483_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13832_ _13832_/A vssd1 vssd1 vccd1 vccd1 _13845_/S sky130_fd_sc_hd__clkbuf_4
X_16620_ _16620_/A vssd1 vssd1 vccd1 vccd1 _16627_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16551_ _19623_/Q _16548_/C _16550_/Y vssd1 vssd1 vccd1 vccd1 _19623_/D sky130_fd_sc_hd__o21a_1
X_13763_ _13763_/A vssd1 vssd1 vccd1 vccd1 _18542_/D sky130_fd_sc_hd__clkbuf_1
X_10975_ _18578_/Q _18839_/Q _18738_/Q _19073_/Q _10018_/A _10974_/X vssd1 vssd1 vccd1
+ vccd1 _10975_/X sky130_fd_sc_hd__mux4_1
XANTENNA__18266__S _18268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11182__S0 _10017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15502_ _15502_/A vssd1 vssd1 vccd1 vccd1 _15511_/S sky130_fd_sc_hd__buf_4
X_12714_ _12714_/A vssd1 vssd1 vccd1 vccd1 _12714_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19270_ _19272_/CLK _19270_/D vssd1 vssd1 vccd1 vccd1 _19270_/Q sky130_fd_sc_hd__dfxtp_1
X_16482_ _16939_/A vssd1 vssd1 vccd1 vccd1 _16482_/X sky130_fd_sc_hd__clkbuf_2
X_13694_ _18526_/Q _13693_/X _13694_/S vssd1 vssd1 vccd1 vccd1 _13695_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_52_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15433_ _14660_/X _19220_/Q _15439_/S vssd1 vssd1 vccd1 vccd1 _15434_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18221_ _18221_/A vssd1 vssd1 vccd1 vccd1 _19966_/D sky130_fd_sc_hd__clkbuf_1
X_12645_ _12651_/B _12645_/B vssd1 vssd1 vccd1 vccd1 _12646_/A sky130_fd_sc_hd__and2b_2
XFILLER_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15364_ _15364_/A vssd1 vssd1 vccd1 vccd1 _19189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18152_ _18152_/A vssd1 vssd1 vccd1 vccd1 _19935_/D sky130_fd_sc_hd__clkbuf_1
X_12576_ _12576_/A _18111_/B vssd1 vssd1 vccd1 vccd1 _12577_/B sky130_fd_sc_hd__or2_1
XFILLER_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10598__C1 _09740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12327__B _12328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17103_ _17104_/B _17104_/C _17102_/Y vssd1 vssd1 vccd1 vccd1 _19796_/D sky130_fd_sc_hd__o21a_1
X_14315_ _18770_/Q _13643_/X _14319_/S vssd1 vssd1 vccd1 vccd1 _14316_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15919__A _15975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11527_ _12606_/A vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__clkbuf_2
X_18083_ _18083_/A _18083_/B vssd1 vssd1 vccd1 vccd1 _18083_/X sky130_fd_sc_hd__or2_1
XFILLER_144_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15295_ _15295_/A vssd1 vssd1 vccd1 vccd1 _15295_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10128__A _11384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17034_ _17046_/A _17034_/B _17034_/C vssd1 vssd1 vccd1 vccd1 _19767_/D sky130_fd_sc_hd__nor3_1
XANTENNA_output96_A _11816_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14246_ _13780_/X _18740_/Q _14246_/S vssd1 vssd1 vccd1 vccd1 _14247_/A sky130_fd_sc_hd__mux2_1
X_11458_ _09707_/A _11448_/Y _11453_/X _11457_/Y _09739_/A vssd1 vssd1 vccd1 vccd1
+ _11458_/X sky130_fd_sc_hd__o311a_1
XANTENNA__17278__A0 _15738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ _10403_/A _10408_/X _10323_/X vssd1 vssd1 vccd1 vccd1 _10409_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_171_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14177_ _13783_/X _18709_/Q _14185_/S vssd1 vssd1 vccd1 vccd1 _14178_/A sky130_fd_sc_hd__mux2_1
X_11389_ _18584_/Q _18845_/Q _18744_/Q _19079_/Q _10640_/S _10637_/A vssd1 vssd1 vccd1
+ vccd1 _11389_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12343__A _19534_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15828__A1 _15818_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _15219_/A vssd1 vssd1 vccd1 vccd1 _13128_/X sky130_fd_sc_hd__clkbuf_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17853__B _17853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18985_ _19305_/CLK _18985_/D vssd1 vssd1 vccd1 vccd1 _18985_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _18930_/Q vssd1 vssd1 vccd1 vccd1 _13351_/A sky130_fd_sc_hd__clkbuf_2
X_17936_ _17865_/S _17935_/X _17723_/X vssd1 vssd1 vccd1 vccd1 _17936_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_2_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_17867_ _17616_/A _17863_/Y _17866_/Y _17827_/A vssd1 vssd1 vccd1 vccd1 _17867_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17450__A0 _17884_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19606_ _19988_/CLK _19606_/D vssd1 vssd1 vccd1 vccd1 _19606_/Q sky130_fd_sc_hd__dfxtp_2
X_16818_ _16818_/A _16841_/A vssd1 vssd1 vccd1 vccd1 _16818_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17798_ _17798_/A vssd1 vssd1 vccd1 vccd1 _18083_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_81_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19537_ _19540_/CLK _19537_/D vssd1 vssd1 vccd1 vccd1 _19537_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__11406__B _12649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16749_ _19687_/Q _19686_/Q _19685_/Q _16749_/D vssd1 vssd1 vccd1 vccd1 _16755_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_59_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13902__A _13913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16916__C _16930_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19468_ _19563_/CLK _19468_/D vssd1 vssd1 vccd1 vccd1 _19468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09221_ _09325_/A _09220_/X input33/X vssd1 vssd1 vccd1 vccd1 _16816_/C sky130_fd_sc_hd__o21bai_2
X_18419_ _12475_/A _18413_/X _18414_/X _18418_/Y vssd1 vssd1 vccd1 vccd1 _18420_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_19399_ _19402_/CLK _19399_/D vssd1 vssd1 vccd1 vccd1 _19399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09994__A1 _10730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16424__S _16426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput70 reset vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_12
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11228__S1 _11179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17269__A0 _15718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10987__S0 _11085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09985_ _09985_/A vssd1 vssd1 vccd1 vccd1 _09985_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_130_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11400__S1 _10054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16395__A _16441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15503__S _15511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13812__A _14637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10760_ _09680_/A _10759_/X _10043_/X vssd1 vssd1 vccd1 vccd1 _10760_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09419_ _18196_/S vssd1 vssd1 vccd1 vccd1 _09419_/X sky130_fd_sc_hd__buf_4
Xclkbuf_4_4_0_clock clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__13531__B _13560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ _10691_/A vssd1 vssd1 vccd1 vccd1 _10691_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12430_ _18046_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _12460_/A sky130_fd_sc_hd__xnor2_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12361_ _12361_/A _12361_/B vssd1 vssd1 vccd1 vccd1 _12362_/A sky130_fd_sc_hd__xnor2_4
XFILLER_165_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14100_ _14146_/S vssd1 vssd1 vccd1 vccd1 _14109_/S sky130_fd_sc_hd__buf_2
X_11312_ _11304_/A _11309_/X _11311_/X vssd1 vssd1 vccd1 vccd1 _11312_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_6_clock _19998_/CLK vssd1 vssd1 vccd1 vccd1 _20032_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09737__A _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15080_ _15080_/A vssd1 vssd1 vccd1 vccd1 _19073_/D sky130_fd_sc_hd__clkbuf_1
X_12292_ _12208_/X _12287_/Y _12290_/X _12291_/X vssd1 vssd1 vccd1 vccd1 _12292_/X
+ sky130_fd_sc_hd__o31a_1
X_14031_ _18647_/Q _13664_/X _14035_/S vssd1 vssd1 vccd1 vccd1 _14032_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13259__A _15241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11243_ _11117_/X _11242_/X _11069_/X vssd1 vssd1 vccd1 vccd1 _11243_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09832__S1 _09822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11174_ _11295_/A _11173_/X _10980_/A vssd1 vssd1 vccd1 vccd1 _11174_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14789__S _14797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10125_ _10846_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10125_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18770_ _19491_/CLK _18770_/D vssd1 vssd1 vccd1 vccd1 _18770_/Q sky130_fd_sc_hd__dfxtp_1
X_15982_ _19416_/Q _15289_/X _15984_/S vssd1 vssd1 vccd1 vccd1 _15983_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09472__A _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17721_ _17721_/A _17721_/B _17721_/C vssd1 vssd1 vccd1 vccd1 _17722_/A sky130_fd_sc_hd__or3_2
X_10056_ _10056_/A vssd1 vssd1 vccd1 vccd1 _10056_/X sky130_fd_sc_hd__clkbuf_4
X_14933_ _19008_/Q _14392_/X _14939_/S vssd1 vssd1 vccd1 vccd1 _14934_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17432__A0 _17702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17652_ _17449_/X _17486_/X _17686_/S vssd1 vssd1 vccd1 vccd1 _17652_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10411__A _19912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14864_ _14864_/A vssd1 vssd1 vccd1 vccd1 _18977_/D sky130_fd_sc_hd__clkbuf_1
X_16603_ _19641_/Q _16601_/B _16577_/X vssd1 vssd1 vccd1 vccd1 _16603_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13815_ _14640_/A vssd1 vssd1 vccd1 vccd1 _13815_/X sky130_fd_sc_hd__clkbuf_1
X_14795_ _18951_/Q _14430_/X _14797_/S vssd1 vssd1 vccd1 vccd1 _14796_/A sky130_fd_sc_hd__mux2_1
X_17583_ _17488_/X _17479_/X _17590_/S vssd1 vssd1 vccd1 vccd1 _17583_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15413__S _15417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13722__A _15283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19322_ _19594_/CLK hold17/X vssd1 vssd1 vccd1 vccd1 _19322_/Q sky130_fd_sc_hd__dfxtp_1
X_16534_ _16538_/B _16538_/C _16533_/X vssd1 vssd1 vccd1 vccd1 _16534_/Y sky130_fd_sc_hd__a21oi_1
X_13746_ _14574_/A vssd1 vssd1 vccd1 vccd1 _13746_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10958_ _11202_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _10958_/X sky130_fd_sc_hd__or2_1
XFILLER_32_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17735__A1 _19897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19253_ _19511_/CLK _19253_/D vssd1 vssd1 vccd1 vccd1 _19253_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14029__S _14035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13677_ _13719_/A vssd1 vssd1 vccd1 vccd1 _13694_/S sky130_fd_sc_hd__clkbuf_4
X_16465_ _18352_/A _16465_/B vssd1 vssd1 vccd1 vccd1 _16466_/A sky130_fd_sc_hd__or2_1
X_10889_ _11478_/A _10889_/B vssd1 vssd1 vccd1 vccd1 _10889_/X sky130_fd_sc_hd__or2_1
X_18204_ _18204_/A vssd1 vssd1 vccd1 vccd1 _19958_/D sky130_fd_sc_hd__clkbuf_1
X_15416_ _15416_/A vssd1 vssd1 vccd1 vccd1 _19212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12628_ _12628_/A _12628_/B vssd1 vssd1 vccd1 vccd1 _12628_/Y sky130_fd_sc_hd__nand2_1
X_19184_ _19412_/CLK _19184_/D vssd1 vssd1 vccd1 vccd1 _19184_/Q sky130_fd_sc_hd__dfxtp_1
X_16396_ _13219_/X _19556_/Q _16404_/S vssd1 vssd1 vccd1 vccd1 _16397_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17499__A0 _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15347_ _15358_/A vssd1 vssd1 vccd1 vccd1 _15356_/S sky130_fd_sc_hd__buf_2
X_18135_ _18135_/A vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__clkbuf_1
XFILLER_145_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12559_ _12559_/A _12559_/B vssd1 vssd1 vccd1 vccd1 _12559_/Y sky130_fd_sc_hd__nor2_8
XFILLER_144_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09647__A _09647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15278_ _15278_/A vssd1 vssd1 vccd1 vccd1 _19154_/D sky130_fd_sc_hd__clkbuf_1
X_18066_ _18068_/A _18068_/B _18088_/S vssd1 vssd1 vccd1 vccd1 _18066_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14229_ _13755_/X _18732_/Q _14235_/S vssd1 vssd1 vccd1 vccd1 _14230_/A sky130_fd_sc_hd__mux2_1
X_17017_ _17027_/D vssd1 vssd1 vccd1 vccd1 _17025_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09823__S1 _09822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09770_ _09567_/A _09767_/X _09769_/X _09580_/X vssd1 vssd1 vccd1 vccd1 _09771_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ _19671_/CLK _18968_/D vssd1 vssd1 vccd1 vccd1 _18968_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _17919_/A _17919_/B _17919_/C _17919_/D vssd1 vssd1 vccd1 vccd1 _17919_/X
+ sky130_fd_sc_hd__or4_1
X_18899_ _19487_/CLK _18899_/D vssd1 vssd1 vccd1 vccd1 _18899_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11394__S0 _10640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16943__A _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ _11648_/A vssd1 vssd1 vccd1 vccd1 _12601_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13212__A1 _15722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18151__A1 _19967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10577__A2 _10567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__A _10606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15993__S _16001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09968_ _10675_/A vssd1 vssd1 vccd1 vccd1 _10735_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__14402__S _14402_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09899_ _09899_/A vssd1 vssd1 vccd1 vccd1 _09899_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11324__A1_N _11313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11930_ _17772_/A _11930_/B vssd1 vssd1 vccd1 vccd1 _11932_/A sky130_fd_sc_hd__xnor2_2
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ _11861_/A _11861_/B vssd1 vssd1 vccd1 vccd1 _11933_/A sky130_fd_sc_hd__nor2_2
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _18468_/Q _13600_/B vssd1 vssd1 vccd1 vccd1 _13600_/X sky130_fd_sc_hd__or2_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _18805_/Q _19140_/Q _10812_/S vssd1 vssd1 vccd1 vccd1 _10813_/B sky130_fd_sc_hd__mux2_1
XANTENNA__17014__A _17046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14580_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11792_ _19580_/Q _11792_/B vssd1 vssd1 vccd1 vccd1 _11792_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13451__A1 _13054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13531_ _19880_/Q _13560_/A vssd1 vssd1 vccd1 vccd1 _13531_/X sky130_fd_sc_hd__and2_1
X_10743_ _11440_/A _10743_/B vssd1 vssd1 vccd1 vccd1 _10743_/X sky130_fd_sc_hd__or2_1
XANTENNA__11462__B1 _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17949__A _17949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16250_ _16255_/B _16250_/B vssd1 vssd1 vccd1 vccd1 _16250_/Y sky130_fd_sc_hd__nand2_1
X_13462_ _19876_/Q _12992_/X _13205_/X _19843_/Q vssd1 vssd1 vccd1 vccd1 _13462_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10674_ _11569_/A vssd1 vssd1 vccd1 vccd1 _10674_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ _19130_/Q _15197_/X _15213_/S vssd1 vssd1 vccd1 vccd1 _15202_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12413_ _12413_/A _12413_/B vssd1 vssd1 vccd1 vccd1 _12414_/A sky130_fd_sc_hd__xnor2_2
X_16181_ _19504_/Q _14640_/A _16189_/S vssd1 vssd1 vccd1 vccd1 _16182_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15469__A _15515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13393_ _15267_/A vssd1 vssd1 vccd1 vccd1 _13393_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14373__A _14472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18142__A1 _19963_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_154_clock clkbuf_opt_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19718_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15132_ _15132_/A vssd1 vssd1 vccd1 vccd1 _19097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12344_ _19837_/Q vssd1 vssd1 vccd1 vccd1 _17210_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15063_ _15131_/S vssd1 vssd1 vccd1 vccd1 _15072_/S sky130_fd_sc_hd__clkbuf_4
X_19940_ _19987_/CLK _19940_/D vssd1 vssd1 vccd1 vccd1 _19940_/Q sky130_fd_sc_hd__dfxtp_1
X_12275_ _12303_/S vssd1 vssd1 vccd1 vccd1 _12573_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11517__A1 _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ _14014_/A vssd1 vssd1 vccd1 vccd1 _18639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11226_ _10969_/A _11223_/Y _11225_/Y _10899_/A vssd1 vssd1 vccd1 vccd1 _11226_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19871_ _19873_/CLK _19871_/D vssd1 vssd1 vccd1 vccd1 _19871_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_169_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19988_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13717__A _15279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18822_ _19478_/CLK _18822_/D vssd1 vssd1 vccd1 vccd1 _18822_/Q sky130_fd_sc_hd__dfxtp_1
X_11157_ _19897_/Q vssd1 vssd1 vccd1 vccd1 _11157_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10108_ _10665_/A vssd1 vssd1 vccd1 vccd1 _11387_/A sky130_fd_sc_hd__buf_4
X_18753_ _19476_/CLK _18753_/D vssd1 vssd1 vccd1 vccd1 _18753_/Q sky130_fd_sc_hd__dfxtp_1
X_15965_ _19408_/Q _15263_/X _15973_/S vssd1 vssd1 vccd1 vccd1 _15966_/A sky130_fd_sc_hd__mux2_1
X_11088_ _19103_/Q _18869_/Q _19551_/Q _19199_/Q _10017_/A _10917_/A vssd1 vssd1 vccd1
+ vccd1 _11088_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10179__S1 _09929_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11376__S0 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17704_ _17794_/A vssd1 vssd1 vccd1 vccd1 _17705_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10039_ _10039_/A vssd1 vssd1 vccd1 vccd1 _10652_/A sky130_fd_sc_hd__clkbuf_2
X_14916_ _14916_/A vssd1 vssd1 vccd1 vccd1 _19001_/D sky130_fd_sc_hd__clkbuf_1
X_18684_ _19051_/CLK _18684_/D vssd1 vssd1 vccd1 vccd1 _18684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15896_ _15896_/A vssd1 vssd1 vccd1 vccd1 _19377_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17956__A1 _19909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17635_ _17675_/S vssd1 vssd1 vccd1 vccd1 _17760_/S sky130_fd_sc_hd__clkbuf_2
X_14847_ _14915_/S vssd1 vssd1 vccd1 vccd1 _14856_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_63_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14548__A _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17566_ _17564_/X _17565_/X _17802_/D vssd1 vssd1 vccd1 vccd1 _17566_/X sky130_fd_sc_hd__mux2_1
X_14778_ _18943_/Q _14404_/X _14786_/S vssd1 vssd1 vccd1 vccd1 _14779_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_107_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19398_/CLK sky130_fd_sc_hd__clkbuf_16
X_19305_ _19305_/CLK _19305_/D vssd1 vssd1 vccd1 vccd1 _19305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15719__A0 _19902_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16517_ _16518_/B _16518_/C _19613_/Q vssd1 vssd1 vccd1 vccd1 _16519_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__13171__B _13299_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13729_ _13729_/A vssd1 vssd1 vccd1 vccd1 _18534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17497_ _17495_/X _17496_/X _17500_/S vssd1 vssd1 vccd1 vccd1 _17497_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19236_ _19268_/CLK _19236_/D vssd1 vssd1 vccd1 vccd1 _19236_/Q sky130_fd_sc_hd__dfxtp_1
X_16448_ _16448_/A vssd1 vssd1 vccd1 vccd1 _19579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19167_ _19391_/CLK _19167_/D vssd1 vssd1 vccd1 vccd1 _19167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16379_ _16379_/A vssd1 vssd1 vccd1 vccd1 _19548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09377__A _13527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12953__B1 _10869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18118_ _18118_/A _18118_/B vssd1 vssd1 vccd1 vccd1 _18118_/X sky130_fd_sc_hd__or2_1
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19098_ _19290_/CLK _19098_/D vssd1 vssd1 vccd1 vccd1 _19098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17892__A0 _19905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18049_ _17971_/A _17806_/B _18048_/X _17796_/X vssd1 vssd1 vccd1 vccd1 _18049_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_160_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11508__A1 _10039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_174_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15826__B _18465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12181__A1 _19528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09822_ _09822_/A vssd1 vssd1 vccd1 vccd1 _09822_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20011_ _20020_/CLK _20011_/D vssd1 vssd1 vccd1 vccd1 _20011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14222__S _14222_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16003__A _16060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09753_ _09753_/A vssd1 vssd1 vccd1 vccd1 _10065_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11367__S0 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__A _11147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ _09884_/A vssd1 vssd1 vccd1 vccd1 _10283_/A sky130_fd_sc_hd__buf_2
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11119__S0 _11004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15053__S _15055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10247__A1 _10196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15988__S _15988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14892__S _14900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_99_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_71_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19313_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15289__A _15289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10390_ _18686_/Q _19181_/Q _10390_/S vssd1 vssd1 vccd1 vccd1 _10391_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_86_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19557_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09799__S0 _09726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ _12153_/A _11976_/B _12059_/X _11825_/A vssd1 vssd1 vccd1 vccd1 _12060_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_151_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15736__B _15736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11011_ _11016_/A _11008_/X _11010_/X _10949_/X vssd1 vssd1 vccd1 vccd1 _11012_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15752__A _15806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15750_ _18452_/Q _13289_/X _15749_/Y _15700_/X vssd1 vssd1 vccd1 vccd1 _15750_/X
+ sky130_fd_sc_hd__o211a_1
X_12962_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12962_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17938__A1 _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A io_dbus_rdata[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09340__A2 _16809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _12240_/B _12153_/B _12153_/A _11913_/D vssd1 vssd1 vccd1 vccd1 _11913_/X
+ sky130_fd_sc_hd__and4b_1
X_14701_ _14701_/A vssd1 vssd1 vccd1 vccd1 _18904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19405_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09971__S0 _10735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _12893_/A _12893_/B vssd1 vssd1 vccd1 vccd1 _12893_/X sky130_fd_sc_hd__and2_1
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15681_ _13580_/X _15679_/X _15680_/Y _13577_/A _18441_/Q vssd1 vssd1 vccd1 vccd1
+ _17160_/A sky130_fd_sc_hd__a32oi_4
XFILLER_61_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _17729_/B _12501_/A _17450_/S vssd1 vssd1 vccd1 vccd1 _17420_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14632_ _14631_/X _18881_/Q _14638_/S vssd1 vssd1 vccd1 vccd1 _14633_/A sky130_fd_sc_hd__mux2_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _11843_/A _11843_/B _11843_/C vssd1 vssd1 vccd1 vccd1 _11844_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14563_/A vssd1 vssd1 vccd1 vccd1 _18858_/D sky130_fd_sc_hd__clkbuf_1
X_17351_ _17355_/A _17351_/B vssd1 vssd1 vccd1 vccd1 _17352_/A sky130_fd_sc_hd__and2_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _19817_/Q _13604_/A vssd1 vssd1 vccd1 vccd1 _11776_/A sky130_fd_sc_hd__and2_1
XANTENNA__16583__A _16629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16301_/A _16301_/C _16301_/B vssd1 vssd1 vccd1 vccd1 _16302_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19053_/CLK sky130_fd_sc_hd__clkbuf_16
X_13514_ _19879_/Q _12699_/A _13205_/X _19846_/Q vssd1 vssd1 vccd1 vccd1 _13514_/X
+ sky130_fd_sc_hd__a22o_1
X_10726_ _10727_/A _12648_/A vssd1 vssd1 vccd1 vccd1 _10728_/A sky130_fd_sc_hd__nand2_1
X_17282_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17291_/S sky130_fd_sc_hd__buf_2
X_14494_ _14828_/A _18410_/B vssd1 vssd1 vccd1 vccd1 _18829_/D sky130_fd_sc_hd__nor2_4
Xclkbuf_3_1_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_19021_ _19439_/CLK _19021_/D vssd1 vssd1 vccd1 vccd1 _19021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15199__A hold10/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13445_ _19349_/Q _13245_/X _13099_/X _19539_/Q _13444_/X vssd1 vssd1 vccd1 vccd1
+ _13445_/X sky130_fd_sc_hd__a221o_1
X_16233_ _16232_/A _16232_/C _13115_/A vssd1 vssd1 vccd1 vccd1 _16233_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_173_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10657_ _10642_/X _10647_/Y _10651_/Y _10656_/Y _09739_/A vssd1 vssd1 vccd1 vccd1
+ _10657_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11520__A _11520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16164_ _16164_/A vssd1 vssd1 vccd1 vccd1 _19496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13376_ _15263_/A vssd1 vssd1 vccd1 vccd1 _13376_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10588_ _10588_/A _10588_/B vssd1 vssd1 vccd1 vccd1 _10588_/Y sky130_fd_sc_hd__nor2_1
X_15115_ _15115_/A vssd1 vssd1 vccd1 vccd1 _19089_/D sky130_fd_sc_hd__clkbuf_1
X_12327_ _12329_/A _12328_/A vssd1 vssd1 vccd1 vccd1 _12330_/A sky130_fd_sc_hd__and2_1
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16095_ _13277_/X _19466_/Q _16095_/S vssd1 vssd1 vccd1 vccd1 _16096_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10136__A _10137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14831__A _14831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18303__A _18341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15046_ _15046_/A vssd1 vssd1 vccd1 vccd1 _15055_/S sky130_fd_sc_hd__buf_4
X_19923_ _19978_/CLK _19923_/D vssd1 vssd1 vccd1 vccd1 _19923_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12258_ _12228_/A _17949_/A _12232_/A _12232_/B vssd1 vssd1 vccd1 vccd1 _12259_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11209_ _09472_/A _11202_/X _11204_/X _11208_/X _09600_/A vssd1 vssd1 vccd1 vccd1
+ _11209_/X sky130_fd_sc_hd__a311o_2
XANTENNA__14042__S _14046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19854_ _19881_/CLK _19854_/D vssd1 vssd1 vccd1 vccd1 _19854_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12351__A _12429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ _12189_/A vssd1 vssd1 vccd1 vccd1 _17334_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18805_ _19366_/CLK _18805_/D vssd1 vssd1 vccd1 vccd1 _18805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19785_ _19805_/CLK _19785_/D vssd1 vssd1 vccd1 vccd1 _19785_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14977__S _14983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16997_ _19756_/Q _16993_/C _16996_/Y vssd1 vssd1 vccd1 vccd1 _19756_/D sky130_fd_sc_hd__o21a_1
XFILLER_95_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13881__S _13889_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18736_ _19551_/CLK _18736_/D vssd1 vssd1 vccd1 vccd1 _18736_/Q sky130_fd_sc_hd__dfxtp_1
X_15948_ _15948_/A vssd1 vssd1 vccd1 vccd1 _19400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11123__C1 _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18667_ _19258_/CLK _18667_/D vssd1 vssd1 vccd1 vccd1 _18667_/Q sky130_fd_sc_hd__dfxtp_1
X_15879_ _13277_/X _19370_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15880_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12871__C1 _12870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17618_ _17940_/A vssd1 vssd1 vccd1 vccd1 _17619_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13316__D_N _12764_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18598_ _19573_/CLK _18598_/D vssd1 vssd1 vccd1 vccd1 _18598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17549_ _17549_/A _17549_/B vssd1 vssd1 vccd1 vccd1 _17940_/A sky130_fd_sc_hd__nor2_2
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18354__B2 input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16365__A0 _19544_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19219_ _19313_/CLK _19219_/D vssd1 vssd1 vccd1 vccd1 _19219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18106__A1 _12559_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09835__A _10559_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17617__B1 _17533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13357__A _15260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input2_A io_dbus_rdata[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _09750_/X _09794_/X _09803_/X _09757_/X _09804_/Y vssd1 vssd1 vccd1 vccd1
+ _12667_/B sky130_fd_sc_hd__o32a_4
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14887__S _14889_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13791__S _13797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09736_ _09736_/A vssd1 vssd1 vccd1 vccd1 _09737_/A sky130_fd_sc_hd__buf_2
XFILLER_86_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10468__A1 _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _09667_/A vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__buf_2
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09598_ _18969_/Q vssd1 vssd1 vccd1 vccd1 _09599_/A sky130_fd_sc_hd__inv_2
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15511__S _15511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11560_ _11560_/A _11563_/A _11560_/C vssd1 vssd1 vccd1 vccd1 _11560_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__12090__B1 _12855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10511_ _18683_/Q _19178_/Q _10560_/S vssd1 vssd1 vccd1 vccd1 _10511_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14127__S _14131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ _11491_/A _11491_/B _11491_/C vssd1 vssd1 vccd1 vccd1 _11491_/X sky130_fd_sc_hd__or3_2
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13031__S _13554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ _15235_/A vssd1 vssd1 vccd1 vccd1 _13230_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10442_ _18589_/Q _18850_/Q _18749_/Q _19084_/Q _10337_/X _10326_/X vssd1 vssd1 vccd1
+ vccd1 _10442_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13966__S _13972_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09794__C1 _09741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13161_ _16864_/C _12719_/X _12723_/X _16737_/B _13160_/X vssd1 vssd1 vccd1 vccd1
+ _15709_/B sky130_fd_sc_hd__a221o_2
X_10373_ _10373_/A _10373_/B vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__or2_1
XFILLER_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12112_ _12112_/A vssd1 vssd1 vccd1 vccd1 _12117_/B sky130_fd_sc_hd__inv_6
XANTENNA__09745__A _09745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input58_A io_ibus_inst[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _19930_/Q vssd1 vssd1 vccd1 vccd1 _16232_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10390__S _10390_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16920_ _19721_/Q _16920_/B _16920_/C vssd1 vssd1 vccd1 vccd1 _16921_/D sky130_fd_sc_hd__and3_1
X_12043_ _12104_/A _12104_/C vssd1 vssd1 vccd1 vccd1 _12044_/B sky130_fd_sc_hd__nor2_1
XFILLER_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16851_ _16864_/A _16857_/D _16768_/X vssd1 vssd1 vccd1 vccd1 _16851_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14797__S _14797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15802_ _15802_/A vssd1 vssd1 vccd1 vccd1 _19348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19570_ _19570_/CLK _19570_/D vssd1 vssd1 vccd1 vccd1 _19570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16782_ _16874_/A _16782_/B _16784_/B vssd1 vssd1 vccd1 vccd1 _19698_/D sky130_fd_sc_hd__nor3_1
XANTENNA__12448__A2 _11771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13994_ _18632_/Q _13735_/X _13994_/S vssd1 vssd1 vccd1 vccd1 _13995_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18521_ _19498_/CLK _18521_/D vssd1 vssd1 vccd1 vccd1 _18521_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _19905_/Q _12874_/X _15757_/S vssd1 vssd1 vccd1 vccd1 _15733_/X sky130_fd_sc_hd__mux2_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _18028_/A vssd1 vssd1 vccd1 vccd1 _12951_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _19952_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _15808_/A vssd1 vssd1 vccd1 vccd1 _15844_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_122_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _16528_/A _19773_/Q _17129_/S _12875_/X vssd1 vssd1 vccd1 vccd1 _19773_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _18121_/A _12615_/B _17387_/Y _17388_/X _17966_/A vssd1 vssd1 vccd1 vccd1
+ _17403_/X sky130_fd_sc_hd__a41o_1
X_14615_ _14615_/A vssd1 vssd1 vccd1 vccd1 _14615_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _11827_/A vssd1 vssd1 vccd1 vccd1 _11915_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18383_ _20030_/Q _18373_/X _18374_/X _18382_/Y vssd1 vssd1 vccd1 vccd1 _18384_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15595_ _15595_/A vssd1 vssd1 vccd1 vccd1 _19291_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11959__A1 _16226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13730__A _15289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17334_ _18118_/A _17334_/B _17333_/X vssd1 vssd1 vccd1 vccd1 _17335_/C sky130_fd_sc_hd__or3b_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _13812_/X _18851_/Q _14546_/S vssd1 vssd1 vccd1 vccd1 _14547_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11758_ _11849_/C vssd1 vssd1 vccd1 vccd1 _17675_/S sky130_fd_sc_hd__buf_2
XANTENNA__17544__C1 _17543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ _18583_/Q _18844_/Q _18743_/Q _19078_/Q _10653_/X _10665_/X vssd1 vssd1 vccd1
+ vccd1 _10709_/X sky130_fd_sc_hd__mux4_2
X_17265_ _17141_/A _19857_/Q _17269_/S vssd1 vssd1 vccd1 vccd1 _17266_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14477_ _14477_/A _14477_/B _14477_/C _11792_/B vssd1 vssd1 vccd1 vccd1 _14478_/B
+ sky130_fd_sc_hd__or4b_1
X_11689_ _11699_/A vssd1 vssd1 vccd1 vccd1 _11894_/A sky130_fd_sc_hd__clkbuf_2
X_19004_ _19484_/CLK _19004_/D vssd1 vssd1 vccd1 vccd1 _19004_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11250__A _11250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16216_ _16213_/X _16215_/Y _13597_/B vssd1 vssd1 vccd1 vccd1 _16216_/X sky130_fd_sc_hd__a21o_1
XFILLER_139_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13428_ _13428_/A _13438_/C vssd1 vssd1 vccd1 vccd1 _13428_/Y sky130_fd_sc_hd__nand2_1
X_17196_ _17194_/Y _17182_/X _17195_/X _17185_/X vssd1 vssd1 vccd1 vccd1 _19832_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13876__S _13878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ _13359_/A vssd1 vssd1 vccd1 vccd1 _18488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16147_ _16204_/S vssd1 vssd1 vccd1 vccd1 _16156_/S sky130_fd_sc_hd__buf_2
XFILLER_127_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16078_ _13128_/X _19458_/Q _16084_/S vssd1 vssd1 vccd1 vccd1 _16079_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_47_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15029_ _19051_/Q _14427_/X _15033_/S vssd1 vssd1 vccd1 vccd1 _15030_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19906_ _19906_/CLK _19906_/D vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_4
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10242__S0 _09902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19837_ _19837_/CLK _19837_/D vssd1 vssd1 vccd1 vccd1 _19837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10793__S1 _11496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16919__C _16955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 io_dbus_rdata[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_6
X_19768_ _19768_/CLK _19768_/D vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfxtp_1
XFILLER_110_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09521_ _09822_/A vssd1 vssd1 vccd1 vccd1 _09809_/A sky130_fd_sc_hd__clkbuf_4
X_18719_ _19311_/CLK _18719_/D vssd1 vssd1 vccd1 vccd1 _18719_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09935__S0 _10218_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19699_ _19737_/CLK _19699_/D vssd1 vssd1 vccd1 vccd1 _19699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09452_ _17338_/A _18343_/A _17339_/A vssd1 vssd1 vccd1 vccd1 _09452_/X sky130_fd_sc_hd__and3_1
XFILLER_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09383_ _12702_/A vssd1 vssd1 vccd1 vccd1 _18326_/A sky130_fd_sc_hd__inv_2
XFILLER_52_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18327__A1 _17339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10622__A1 _11440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16951__A _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13815__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10784__S1 _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09719_ _09719_/A vssd1 vssd1 vccd1 vccd1 _09719_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10991_ _11025_/A _10991_/B vssd1 vssd1 vccd1 vccd1 _10991_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17369__A2 _18301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _19790_/Q vssd1 vssd1 vccd1 vccd1 _17087_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12661_ _12663_/A _12661_/B vssd1 vssd1 vccd1 vccd1 _12661_/Y sky130_fd_sc_hd__nor2_8
XFILLER_15_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18118__A _18118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _18138_/A vssd1 vssd1 vccd1 vccd1 _11657_/S sky130_fd_sc_hd__buf_6
X_14400_ _14400_/A vssd1 vssd1 vccd1 vccd1 _18803_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15380_ _14583_/X _19196_/Q _15384_/S vssd1 vssd1 vccd1 vccd1 _15381_/A sky130_fd_sc_hd__mux2_1
X_12592_ _12188_/X _12670_/B _12319_/B vssd1 vssd1 vccd1 vccd1 _18118_/B sky130_fd_sc_hd__a21bo_1
XFILLER_129_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11810__A0 _19960_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14331_ _14331_/A vssd1 vssd1 vccd1 vccd1 _18777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11543_ _11543_/A vssd1 vssd1 vccd1 vccd1 _11544_/C sky130_fd_sc_hd__inv_2
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14262_ _13803_/X _18747_/Q _14268_/S vssd1 vssd1 vccd1 vccd1 _14263_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17050_ _17053_/B _17053_/C _17021_/X vssd1 vssd1 vccd1 vccd1 _17050_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11474_ _19514_/Q _18926_/Q _18963_/Q _18537_/Q _09532_/A _09514_/A vssd1 vssd1 vccd1
+ vccd1 _11475_/B sky130_fd_sc_hd__mux4_1
XFILLER_167_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16001_ _13089_/X _19424_/Q _16001_/S vssd1 vssd1 vccd1 vccd1 _16002_/A sky130_fd_sc_hd__mux2_1
X_13213_ _13191_/A _13214_/C _19935_/Q vssd1 vssd1 vccd1 vccd1 _13215_/B sky130_fd_sc_hd__a21oi_1
X_10425_ _19502_/Q _18914_/Q _18951_/Q _18525_/Q _10367_/S _10291_/X vssd1 vssd1 vccd1
+ vccd1 _10426_/B sky130_fd_sc_hd__mux4_1
XFILLER_109_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14193_ _14193_/A vssd1 vssd1 vccd1 vccd1 _18716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09475__A _09475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13144_ _13143_/X _19713_/Q _13144_/S vssd1 vssd1 vccd1 vccd1 _13144_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10356_ _10448_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output164_A _11799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12613__B _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _19778_/Q vssd1 vssd1 vccd1 vccd1 _17053_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17952_ _17765_/X _17931_/X _17951_/X _17940_/X vssd1 vssd1 vccd1 vccd1 _17952_/X
+ sky130_fd_sc_hd__a211o_1
X_10287_ _19914_/Q vssd1 vssd1 vccd1 vccd1 _10287_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16903_ _16924_/B _16924_/C _16906_/D _16875_/X vssd1 vssd1 vccd1 vccd1 _16903_/X
+ sky130_fd_sc_hd__a31o_1
X_12026_ _12214_/A vssd1 vssd1 vccd1 vccd1 _12026_/X sky130_fd_sc_hd__clkbuf_4
X_17883_ _17917_/A _17883_/B vssd1 vssd1 vccd1 vccd1 _17885_/C sky130_fd_sc_hd__nor2_1
X_19622_ _19759_/CLK _19622_/D vssd1 vssd1 vccd1 vccd1 _19622_/Q sky130_fd_sc_hd__dfxtp_1
X_16834_ _19711_/Q _16829_/B _16833_/X vssd1 vssd1 vccd1 vccd1 _16835_/B sky130_fd_sc_hd__o21ai_1
XFILLER_38_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09917__S0 _10245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19553_ _19553_/CLK _19553_/D vssd1 vssd1 vccd1 vccd1 _19553_/Q sky130_fd_sc_hd__dfxtp_1
X_16765_ _19693_/Q _16765_/B vssd1 vssd1 vccd1 vccd1 _16772_/C sky130_fd_sc_hd__and2_1
X_13977_ _18624_/Q _13702_/X _13983_/S vssd1 vssd1 vccd1 vccd1 _13978_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18504_ _19745_/CLK _18504_/D vssd1 vssd1 vccd1 vccd1 _18504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15716_ _18446_/Q _15716_/B vssd1 vssd1 vccd1 vccd1 _15716_/X sky130_fd_sc_hd__or2_1
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19484_ _19484_/CLK _19484_/D vssd1 vssd1 vccd1 vccd1 _19484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _18311_/A _11324_/X _12942_/S vssd1 vssd1 vccd1 vccd1 _12928_/X sky130_fd_sc_hd__mux2_2
X_16696_ _19774_/Q _19775_/Q _19777_/Q _19776_/Q vssd1 vssd1 vccd1 vccd1 _17047_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18435_ _18435_/A _18435_/B vssd1 vssd1 vccd1 vccd1 _20052_/D sky130_fd_sc_hd__nor2_1
X_15647_ _14656_/X _19315_/Q _15655_/S vssd1 vssd1 vccd1 vccd1 _15648_/A sky130_fd_sc_hd__mux2_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _16315_/A _12854_/X _12856_/X _17319_/B _12893_/A vssd1 vssd1 vccd1 vccd1
+ _12859_/X sky130_fd_sc_hd__o32a_1
XFILLER_22_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13460__A _16347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18366_ _18366_/A vssd1 vssd1 vccd1 vccd1 _20025_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11899__B _11899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15578_ _15578_/A vssd1 vssd1 vccd1 vccd1 _19284_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17317_ _13603_/B _19881_/Q _17317_/S vssd1 vssd1 vccd1 vccd1 _17318_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14529_ _13787_/X _18843_/Q _14535_/S vssd1 vssd1 vccd1 vccd1 _14530_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10295__S _10417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18297_ _18297_/A _18326_/B vssd1 vssd1 vccd1 vccd1 _18297_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12076__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17248_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17317_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17179_ _15718_/X _17167_/X _17178_/X _17171_/X vssd1 vssd1 vccd1 vccd1 _19826_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10463__S0 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10135__A3 _10133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13635__A _13744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16946__A _16946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ _10466_/S vssd1 vssd1 vccd1 vccd1 _09505_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09435_ _20052_/Q vssd1 vssd1 vccd1 vccd1 _18349_/A sky130_fd_sc_hd__buf_2
XFILLER_80_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10994__A _10994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09366_ _20012_/Q _20011_/Q _20009_/Q _20010_/Q vssd1 vssd1 vccd1 vccd1 _12804_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09297_ _11704_/B _11809_/A _09296_/X vssd1 vssd1 vccd1 vccd1 _09297_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_138_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10210_ _18657_/Q _19248_/Q _19410_/Q _18625_/Q _10162_/S _10196_/A vssd1 vssd1 vccd1
+ vccd1 _10210_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ _11190_/A _11190_/B vssd1 vssd1 vccd1 vccd1 _11190_/X sky130_fd_sc_hd__and2_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10141_ _11544_/A _11543_/A vssd1 vssd1 vccd1 vccd1 _10141_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_clock clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__10206__S0 _10160_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10072_ _09515_/A _10071_/X _10606_/A vssd1 vssd1 vccd1 vccd1 _10072_/X sky130_fd_sc_hd__a21o_1
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11323__A2 _11322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ _13812_/X _18590_/Q _13900_/S vssd1 vssd1 vccd1 vccd1 _13901_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14140__S _14142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14880_ _14902_/A vssd1 vssd1 vccd1 vccd1 _14889_/S sky130_fd_sc_hd__buf_2
X_13831_ _14656_/A vssd1 vssd1 vccd1 vccd1 _13831_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11065__A _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16550_ _16550_/A _16555_/C vssd1 vssd1 vccd1 vccd1 _16550_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13762_ _13761_/X _18542_/Q _13765_/S vssd1 vssd1 vccd1 vccd1 _13763_/A sky130_fd_sc_hd__mux2_1
X_10974_ _10974_/A vssd1 vssd1 vccd1 vccd1 _10974_/X sky130_fd_sc_hd__buf_2
X_15501_ _15501_/A vssd1 vssd1 vccd1 vccd1 _19250_/D sky130_fd_sc_hd__clkbuf_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11182__S1 _10917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12713_ _12995_/A vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16481_ _12340_/A _12537_/X _12347_/X _16480_/X vssd1 vssd1 vccd1 vccd1 _19598_/D
+ sky130_fd_sc_hd__o211a_1
X_13693_ _14637_/A vssd1 vssd1 vccd1 vccd1 _13693_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16067__S _16073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18220_ _19966_/Q hold21/X _18220_/S vssd1 vssd1 vccd1 vccd1 _18221_/A sky130_fd_sc_hd__mux2_1
X_15432_ _15432_/A vssd1 vssd1 vccd1 vccd1 _19219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12644_ _12644_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _12644_/Y sky130_fd_sc_hd__nor2_8
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18151_ _19935_/Q _19967_/Q _18159_/S vssd1 vssd1 vccd1 vccd1 _18152_/A sky130_fd_sc_hd__mux2_1
X_12575_ _12576_/A _18111_/B vssd1 vssd1 vccd1 vccd1 _12618_/A sky130_fd_sc_hd__nand2_2
X_15363_ _19189_/Q _15286_/X _15367_/S vssd1 vssd1 vccd1 vccd1 _15364_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16591__A _16629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17102_ _17104_/B _17104_/C _17101_/X vssd1 vssd1 vccd1 vccd1 _17102_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11004__S _11004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14314_ _14314_/A vssd1 vssd1 vccd1 vccd1 _18769_/D sky130_fd_sc_hd__clkbuf_1
X_11526_ _11645_/B vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__buf_2
X_18082_ _17971_/A _17717_/X _18081_/X _17646_/A vssd1 vssd1 vccd1 vccd1 _18082_/X
+ sky130_fd_sc_hd__a211o_1
X_15294_ _15294_/A vssd1 vssd1 vccd1 vccd1 _19159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17033_ _19767_/Q _19766_/Q _17033_/C vssd1 vssd1 vccd1 vccd1 _17034_/C sky130_fd_sc_hd__and3_1
XFILLER_172_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11457_ _11460_/A _11454_/X _11456_/X vssd1 vssd1 vccd1 vccd1 _11457_/Y sky130_fd_sc_hd__o21ai_1
X_14245_ _14245_/A vssd1 vssd1 vccd1 vccd1 _18739_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14315__S _14319_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10408_ _19471_/Q _19309_/Q _18718_/Q _18488_/Q _10268_/S _10440_/A vssd1 vssd1 vccd1
+ vccd1 _10408_/X sky130_fd_sc_hd__mux4_1
X_14176_ _14222_/S vssd1 vssd1 vccd1 vccd1 _14185_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA_output89_A _12485_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ _10665_/X _11385_/Y _11387_/Y _10648_/A vssd1 vssd1 vccd1 vccd1 _11388_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15828__A2 _18465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16486__C1 _16480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10339_ _10339_/A vssd1 vssd1 vccd1 vccd1 _10588_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13127_ input29/X _12988_/A _13126_/X _13036_/X vssd1 vssd1 vccd1 vccd1 _15219_/A
+ sky130_fd_sc_hd__a22o_2
X_18984_ _19575_/CLK _18984_/D vssd1 vssd1 vccd1 vccd1 _18984_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18311__A _18311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18227__A0 _19969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _13058_/A vssd1 vssd1 vccd1 vccd1 _18471_/D sky130_fd_sc_hd__clkbuf_1
X_17935_ _17933_/B _17937_/A vssd1 vssd1 vccd1 vccd1 _17935_/X sky130_fd_sc_hd__and2b_1
XFILLER_87_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12009_ _12005_/Y _12007_/X _12008_/X vssd1 vssd1 vccd1 vccd1 _12009_/X sky130_fd_sc_hd__o21a_1
X_17866_ _17866_/A _17866_/B vssd1 vssd1 vccd1 vccd1 _17866_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17450__A1 _17985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16817_ _16832_/C vssd1 vssd1 vccd1 vccd1 _16841_/A sky130_fd_sc_hd__clkbuf_1
X_19605_ _19988_/CLK _19605_/D vssd1 vssd1 vccd1 vccd1 _19605_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17797_ _17781_/X _18050_/B _17795_/X _17796_/X vssd1 vssd1 vccd1 vccd1 _17797_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14985__S _14987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19536_ _19988_/CLK _19536_/D vssd1 vssd1 vccd1 vccd1 _19536_/Q sky130_fd_sc_hd__dfxtp_1
X_16748_ _16773_/A _16748_/B _16748_/C vssd1 vssd1 vccd1 vccd1 _19686_/D sky130_fd_sc_hd__nor3_1
XFILLER_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17202__A1 _12741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11173__S1 _10978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19467_ _19561_/CLK _19467_/D vssd1 vssd1 vccd1 vccd1 _19467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16679_ _16898_/A vssd1 vssd1 vccd1 vccd1 _16728_/A sky130_fd_sc_hd__buf_2
XFILLER_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09220_ _19892_/Q _19891_/Q vssd1 vssd1 vccd1 vccd1 _09220_/X sky130_fd_sc_hd__or2_1
XANTENNA__17753__A2 _17743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18418_ input52/X vssd1 vssd1 vccd1 vccd1 _18418_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19398_ _19398_/CLK _19398_/D vssd1 vssd1 vccd1 vccd1 _19398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18349_ _18349_/A _18349_/B vssd1 vssd1 vccd1 vccd1 _18349_/X sky130_fd_sc_hd__or2_1
XFILLER_148_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10684__S0 _10617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17910__C1 _11657_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10753__S _10753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput60 io_ibus_inst[4] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10987__S1 _09659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09984_ _10812_/S vssd1 vssd1 vccd1 vccd1 _09984_/X sky130_fd_sc_hd__buf_4
XFILLER_104_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18218__A0 _19965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17992__A2 _17877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10277__C1 _09741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_169_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12018__A0 _19966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _18138_/A vssd1 vssd1 vccd1 vccd1 _18196_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_10690_ _10826_/S vssd1 vssd1 vccd1 vccd1 _10690_/X sky130_fd_sc_hd__buf_4
XFILLER_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09349_ _09349_/A _09349_/B vssd1 vssd1 vccd1 vccd1 _09350_/A sky130_fd_sc_hd__nor2_1
XFILLER_139_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12360_ _12335_/A _12335_/B _12330_/A vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__a21oi_2
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11311_ _10941_/X _11310_/X _09574_/A vssd1 vssd1 vccd1 vccd1 _11311_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12291_ _19532_/Q _11782_/X _12314_/A vssd1 vssd1 vccd1 vccd1 _12291_/X sky130_fd_sc_hd__o21a_1
X_14030_ _14030_/A vssd1 vssd1 vccd1 vccd1 _18646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10427__S0 _10367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11242_ _18766_/Q _19037_/Q _19261_/Q _19005_/Q _11057_/S _10943_/X vssd1 vssd1 vccd1
+ vccd1 _11242_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12741__B2 _18453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ _18573_/Q _18834_/Q _18733_/Q _19068_/Q _11329_/S _10978_/A vssd1 vssd1 vccd1
+ vccd1 _11173_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18209__A0 _19961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ _19383_/Q _18997_/Q _19447_/Q _18566_/Q _10753_/S _10014_/A vssd1 vssd1 vccd1
+ vccd1 _10125_/B sky130_fd_sc_hd__mux4_1
XANTENNA_input40_A io_ibus_inst[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15981_ _15981_/A vssd1 vssd1 vccd1 vccd1 _19415_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10899__A _10899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17720_ _17627_/X _17871_/A _17719_/X vssd1 vssd1 vccd1 vccd1 _18083_/B sky130_fd_sc_hd__a21oi_2
X_10055_ _19510_/Q _18922_/Q _18959_/Q _18533_/Q _10053_/X _10054_/X vssd1 vssd1 vccd1
+ vccd1 _10055_/X sky130_fd_sc_hd__mux4_1
X_14932_ _14932_/A vssd1 vssd1 vccd1 vccd1 _19007_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17432__A1 _12529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17651_ _17651_/A vssd1 vssd1 vccd1 vccd1 _17651_/Y sky130_fd_sc_hd__inv_2
X_14863_ _14599_/X _18977_/Q _14867_/S vssd1 vssd1 vccd1 vccd1 _14864_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output127_A _12665_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16602_ _19640_/Q _16600_/B _16601_/Y vssd1 vssd1 vccd1 vccd1 _19640_/D sky130_fd_sc_hd__o21a_1
X_13814_ _13814_/A vssd1 vssd1 vccd1 vccd1 _18558_/D sky130_fd_sc_hd__clkbuf_1
X_17582_ _17485_/X _17487_/X _17582_/S vssd1 vssd1 vccd1 vccd1 _17582_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14794_ _14794_/A vssd1 vssd1 vccd1 vccd1 _18950_/D sky130_fd_sc_hd__clkbuf_1
X_19321_ _19577_/CLK _19321_/D vssd1 vssd1 vccd1 vccd1 _19321_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10807__A1 _10746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16533_ _18281_/B vssd1 vssd1 vccd1 vccd1 _16533_/X sky130_fd_sc_hd__buf_2
XFILLER_17_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ _13745_/A vssd1 vssd1 vccd1 vccd1 _18538_/D sky130_fd_sc_hd__clkbuf_1
X_10957_ _19459_/Q _19297_/Q _18706_/Q _18476_/Q _10937_/S _09954_/A vssd1 vssd1 vccd1
+ vccd1 _10958_/B sky130_fd_sc_hd__mux4_1
XANTENNA__17735__A2 _09419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19252_ _19510_/CLK _19252_/D vssd1 vssd1 vccd1 vccd1 _19252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16464_ _16875_/A vssd1 vssd1 vccd1 vccd1 _18352_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15746__A1 _19907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13676_ _14624_/A vssd1 vssd1 vccd1 vccd1 _13676_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10888_ _19492_/Q _18904_/Q _18941_/Q _18515_/Q _09983_/A _10084_/A vssd1 vssd1 vccd1
+ vccd1 _10889_/B sky130_fd_sc_hd__mux4_1
X_18203_ _19958_/Q _19579_/Q _18209_/S vssd1 vssd1 vccd1 vccd1 _18204_/A sky130_fd_sc_hd__mux2_1
X_15415_ _14634_/X _19212_/Q _15417_/S vssd1 vssd1 vccd1 vccd1 _15416_/A sky130_fd_sc_hd__mux2_1
X_19183_ _19409_/CLK _19183_/D vssd1 vssd1 vccd1 vccd1 _19183_/Q sky130_fd_sc_hd__dfxtp_1
X_12627_ _19848_/Q _17240_/A _12588_/B _12626_/Y _12026_/X vssd1 vssd1 vccd1 vccd1
+ _12628_/B sky130_fd_sc_hd__a311o_1
X_16395_ _16441_/S vssd1 vssd1 vccd1 vccd1 _16404_/S sky130_fd_sc_hd__buf_6
XANTENNA__10139__A _10139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18134_ _16219_/A _19960_/Q _18136_/S vssd1 vssd1 vccd1 vccd1 _18135_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17499__A1 _17729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15346_ _15346_/A vssd1 vssd1 vccd1 vccd1 _19181_/D sky130_fd_sc_hd__clkbuf_1
X_12558_ _12532_/A _12535_/A _12555_/Y _12556_/Y vssd1 vssd1 vccd1 vccd1 _12559_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_157_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18065_ _18068_/A _18068_/B vssd1 vssd1 vccd1 vccd1 _18065_/Y sky130_fd_sc_hd__nand2_1
X_11509_ _19482_/Q _19320_/Q _18729_/Q _18499_/Q _10119_/X _10112_/A vssd1 vssd1 vccd1
+ vccd1 _11510_/B sky130_fd_sc_hd__mux4_1
XFILLER_145_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15277_ _19154_/Q _15276_/X _15277_/S vssd1 vssd1 vccd1 vccd1 _15278_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12489_ _19540_/Q _12120_/X _12314_/A vssd1 vssd1 vccd1 vccd1 _12489_/X sky130_fd_sc_hd__o21a_1
X_17016_ _19762_/Q _19761_/Q _17016_/C _17016_/D vssd1 vssd1 vccd1 vccd1 _17027_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_7_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14228_ _14228_/A vssd1 vssd1 vccd1 vccd1 _18731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _13758_/X _18701_/Q _14163_/S vssd1 vssd1 vccd1 vccd1 _14160_/A sky130_fd_sc_hd__mux2_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09663__A _10703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17671__A1 _17670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ _19671_/CLK _18967_/D vssd1 vssd1 vccd1 vccd1 _18967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17918_ _17914_/B _17918_/B vssd1 vssd1 vccd1 vccd1 _17919_/D sky130_fd_sc_hd__and2b_1
XANTENNA__10602__A _10813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18898_ _19486_/CLK _18898_/D vssd1 vssd1 vccd1 vccd1 _18898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11394__S1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17849_ _17849_/A _17853_/A vssd1 vssd1 vccd1 vccd1 _17849_/X sky130_fd_sc_hd__or2_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13913__A _13913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12248__B1 _12494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19519_ _19542_/CLK _19519_/D vssd1 vssd1 vccd1 vccd1 _19519_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12529__A _12529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_170_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16934__B1 _16833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09203_ _09275_/B vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16435__S _16437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09838__A _09904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10577__A3 _10576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12971__A1 _18458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13794__S _13797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16170__S _16178_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_95_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09967_ _09967_/A vssd1 vssd1 vccd1 vccd1 _10675_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15673__A0 _15672_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09292__B _14074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09898_ _09901_/A vssd1 vssd1 vccd1 vccd1 _10197_/S sky130_fd_sc_hd__buf_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14919__A _14987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11860_ _11860_/A _17418_/A vssd1 vssd1 vccd1 vccd1 _11861_/B sky130_fd_sc_hd__nor2_1
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _18677_/Q _19172_/Q _10811_/S vssd1 vssd1 vccd1 vccd1 _10811_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _19580_/Q _11792_/B vssd1 vssd1 vccd1 vccd1 _11868_/C sky130_fd_sc_hd__and2_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13034__S _13090_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11462__A1 _11464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13530_ _19354_/Q _13154_/Y _13155_/Y vssd1 vssd1 vccd1 vccd1 _13530_/X sky130_fd_sc_hd__o21a_1
X_10742_ _19495_/Q _18907_/Q _18944_/Q _18518_/Q _10608_/X _10609_/X vssd1 vssd1 vccd1
+ vccd1 _10743_/B sky130_fd_sc_hd__mux4_2
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10673_ _10673_/A _10673_/B vssd1 vssd1 vccd1 vccd1 _11569_/A sky130_fd_sc_hd__or2_1
XANTENNA__09407__A1 _19813_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13461_ _13491_/C _13460_/Y _11607_/X vssd1 vssd1 vccd1 vccd1 _13461_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09407__B2 _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15200_ _15299_/S vssd1 vssd1 vccd1 vccd1 _15213_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_138_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12412_ _12390_/A _12391_/A _12390_/B _12388_/A vssd1 vssd1 vccd1 vccd1 _12413_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11214__A1 _11141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16180_ _16191_/A vssd1 vssd1 vccd1 vccd1 _16189_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_127_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09748__A _09748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ _13382_/X _13390_/Y _13391_/Y vssd1 vssd1 vccd1 vccd1 _15267_/A sky130_fd_sc_hd__a21oi_4
XFILLER_127_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15131_ _14675_/X _19097_/Q _15131_/S vssd1 vssd1 vccd1 vccd1 _15132_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12343_ _19534_/Q _12584_/B vssd1 vssd1 vccd1 vccd1 _12343_/X sky130_fd_sc_hd__or2_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15062_ _15118_/A vssd1 vssd1 vccd1 vccd1 _15131_/S sky130_fd_sc_hd__buf_4
X_12274_ _17977_/B _12274_/B vssd1 vssd1 vccd1 vccd1 _12278_/A sky130_fd_sc_hd__xnor2_1
XFILLER_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11517__A2 _12668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14013_ _18639_/Q _13630_/X _14013_/S vssd1 vssd1 vccd1 vccd1 _14014_/A sky130_fd_sc_hd__mux2_1
X_11225_ _11225_/A _11225_/B vssd1 vssd1 vccd1 vccd1 _11225_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17102__B1 _17101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19870_ _19873_/CLK _19870_/D vssd1 vssd1 vccd1 vccd1 _19870_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10725__B1 _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09483__A _11014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18821_ _19478_/CLK _18821_/D vssd1 vssd1 vccd1 vccd1 _18821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11156_ _10920_/X _11151_/X _11153_/Y _11155_/Y _09736_/A vssd1 vssd1 vccd1 vccd1
+ _11156_/X sky130_fd_sc_hd__o221a_4
XFILLER_110_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10107_ _10648_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10107_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18752_ _19570_/CLK _18752_/D vssd1 vssd1 vccd1 vccd1 _18752_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11518__A _12593_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15964_ _15975_/A vssd1 vssd1 vccd1 vccd1 _15973_/S sky130_fd_sc_hd__buf_2
XFILLER_110_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11087_ _11032_/A _11083_/X _11086_/Y _10976_/X vssd1 vssd1 vccd1 vccd1 _11087_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17703_ _17616_/A _17698_/Y _17702_/Y vssd1 vssd1 vccd1 vccd1 _17703_/Y sky130_fd_sc_hd__a21oi_1
X_10038_ _18597_/Q _18858_/Q _18757_/Q _19092_/Q _10640_/S _10037_/X vssd1 vssd1 vccd1
+ vccd1 _10038_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11376__S1 _09957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14915_ _14675_/X _19001_/Q _14915_/S vssd1 vssd1 vccd1 vccd1 _14916_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18683_ _19501_/CLK _18683_/D vssd1 vssd1 vccd1 vccd1 _18683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15895_ _13393_/X _19377_/Q _15901_/S vssd1 vssd1 vccd1 vccd1 _15896_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14829__A _16875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__B1 _11170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15424__S _15428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17634_ _17794_/A vssd1 vssd1 vccd1 vccd1 _17634_/X sky130_fd_sc_hd__clkbuf_2
X_14846_ _14902_/A vssd1 vssd1 vccd1 vccd1 _14915_/S sky130_fd_sc_hd__buf_4
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17565_ _17435_/X _17430_/X _17565_/S vssd1 vssd1 vccd1 vccd1 _17565_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14777_ _14823_/S vssd1 vssd1 vccd1 vccd1 _14786_/S sky130_fd_sc_hd__buf_2
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12349__A _20042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ _12042_/A vssd1 vssd1 vccd1 vccd1 _17820_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19304_ _19560_/CLK _19304_/D vssd1 vssd1 vccd1 vccd1 _19304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16516_ _16518_/B _16518_/C _16515_/Y vssd1 vssd1 vccd1 vccd1 _19612_/D sky130_fd_sc_hd__o21a_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13728_ _18534_/Q _13727_/X _13736_/S vssd1 vssd1 vccd1 vccd1 _13729_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15719__A1 _15718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17496_ _12455_/A _11969_/A _17506_/S vssd1 vssd1 vccd1 vccd1 _17496_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19235_ _19493_/CLK _19235_/D vssd1 vssd1 vccd1 vccd1 _19235_/Q sky130_fd_sc_hd__dfxtp_1
X_16447_ _17185_/A _16447_/B vssd1 vssd1 vccd1 vccd1 _16448_/A sky130_fd_sc_hd__and2_1
X_13659_ _15235_/A vssd1 vssd1 vccd1 vccd1 _14612_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19166_ _19391_/CLK _19166_/D vssd1 vssd1 vccd1 vccd1 _19166_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09658__A _09658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16378_ _13056_/X _19548_/Q _16382_/S vssd1 vssd1 vccd1 vccd1 _16379_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18117_ _19923_/Q _17558_/X _18116_/X vssd1 vssd1 vccd1 vccd1 _19923_/D sky130_fd_sc_hd__o21a_1
X_15329_ _15329_/A vssd1 vssd1 vccd1 vccd1 _19173_/D sky130_fd_sc_hd__clkbuf_1
X_19097_ _19129_/CLK _19097_/D vssd1 vssd1 vccd1 vccd1 _19097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18048_ _17785_/X _18045_/X _18047_/Y _17794_/X vssd1 vssd1 vccd1 vccd1 _18048_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_117_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20010_ _20020_/CLK _20010_/D vssd1 vssd1 vccd1 vccd1 _20010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09821_ _09809_/X _09811_/X _09819_/X _10156_/A _09820_/X vssd1 vssd1 vccd1 vccd1
+ _09828_/B sky130_fd_sc_hd__o221a_1
XFILLER_59_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19999_ _20000_/CLK _19999_/D vssd1 vssd1 vccd1 vccd1 _19999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12469__B1 _19842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _09752_/A vssd1 vssd1 vccd1 vccd1 _09753_/A sky130_fd_sc_hd__buf_2
XFILLER_100_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11367__S1 _10609_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09683_ _10407_/A vssd1 vssd1 vccd1 vccd1 _09884_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13643__A _14599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_clock _19998_/CLK vssd1 vssd1 vccd1 vccd1 _19888_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11119__S1 _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16165__S _16167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14474__A _16875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09568__A _09761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15509__S _15511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09799__S1 _09730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12722__A _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ _11202_/A _11010_/B vssd1 vssd1 vccd1 vccd1 _11010_/X sky130_fd_sc_hd__or2_1
XFILLER_78_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10802__S0 _10617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11380__B1 _09612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13121__A1 _19744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15752__B _17194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ _18451_/Q _12959_/X _10672_/A _12954_/X vssd1 vssd1 vccd1 vccd1 _18451_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _18904_/Q _14398_/X _14702_/S vssd1 vssd1 vccd1 vccd1 _14701_/A sky130_fd_sc_hd__mux2_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _19583_/Q _11912_/B vssd1 vssd1 vccd1 vccd1 _11913_/D sky130_fd_sc_hd__or2_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _15680_/A _18441_/Q vssd1 vssd1 vccd1 vccd1 _15680_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11683__A1 _12600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09971__S1 _09970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12892_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14631_ _14631_/A vssd1 vssd1 vccd1 vccd1 _14631_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _11843_/A _11843_/B _11843_/C vssd1 vssd1 vccd1 vccd1 _11843_/X sky130_fd_sc_hd__or3_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__A2 _10227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17350_ _17323_/A _12601_/Y _12824_/A _17358_/A _15819_/B vssd1 vssd1 vccd1 vccd1
+ _17351_/B sky130_fd_sc_hd__a32o_1
X_14562_ _13835_/X _18858_/Q _14568_/S vssd1 vssd1 vccd1 vccd1 _14563_/A sky130_fd_sc_hd__mux2_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11774_/A vssd1 vssd1 vccd1 vccd1 _13604_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16301_ _16301_/A _16301_/B _16301_/C vssd1 vssd1 vccd1 vccd1 _16308_/B sky130_fd_sc_hd__or3_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13699__S _13715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13513_ _13511_/Y _13536_/B _11607_/X vssd1 vssd1 vccd1 vccd1 _13513_/Y sky130_fd_sc_hd__o21ai_1
X_10725_ _09748_/A _10713_/X _10723_/X _09755_/A _10724_/Y vssd1 vssd1 vccd1 vccd1
+ _12648_/A sky130_fd_sc_hd__o32a_4
X_17281_ _17281_/A vssd1 vssd1 vccd1 vccd1 _19864_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _18328_/A _14485_/X _14486_/X _14492_/Y vssd1 vssd1 vccd1 vccd1 _18410_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_19020_ _19051_/CLK _19020_/D vssd1 vssd1 vccd1 vccd1 _19020_/Q sky130_fd_sc_hd__dfxtp_1
X_16232_ _16232_/A _19931_/Q _16232_/C vssd1 vssd1 vccd1 vccd1 _16239_/B sky130_fd_sc_hd__or3_1
XFILLER_146_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13444_ _19875_/Q _12992_/X _13205_/X _19842_/Q vssd1 vssd1 vccd1 vccd1 _13444_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10656_ _10768_/A _10654_/X _10655_/X vssd1 vssd1 vccd1 vccd1 _10656_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16163_ _19496_/Q _14615_/A _16167_/S vssd1 vssd1 vccd1 vccd1 _16164_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11520__B _12669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10587_ _19113_/Q _18879_/Q _19561_/Q _19209_/Q _10533_/S _09665_/A vssd1 vssd1 vccd1
+ vccd1 _10588_/B sky130_fd_sc_hd__mux4_1
XFILLER_103_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13375_ _13363_/X _13373_/Y _13374_/Y vssd1 vssd1 vccd1 vccd1 _15263_/A sky130_fd_sc_hd__a21oi_4
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15114_ _14650_/X _19089_/Q _15116_/S vssd1 vssd1 vccd1 vccd1 _15115_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12326_ _19977_/Q _10363_/A _12528_/S vssd1 vssd1 vccd1 vccd1 _12328_/A sky130_fd_sc_hd__mux2_2
X_16094_ _16094_/A vssd1 vssd1 vccd1 vccd1 _19465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10136__B _12666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15045_ _15045_/A vssd1 vssd1 vccd1 vccd1 _19058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19922_ _19978_/CLK _19922_/D vssd1 vssd1 vccd1 vccd1 _19922_/Q sky130_fd_sc_hd__dfxtp_4
X_12257_ _12257_/A vssd1 vssd1 vccd1 vccd1 _17949_/A sky130_fd_sc_hd__buf_2
XANTENNA__12632__A _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output71_A _12675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12163__A2 _12650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _11202_/A _11205_/X _11207_/X _09574_/A vssd1 vssd1 vccd1 vccd1 _11208_/X
+ sky130_fd_sc_hd__o211a_1
X_19853_ _19857_/CLK _19853_/D vssd1 vssd1 vccd1 vccd1 _19853_/Q sky130_fd_sc_hd__dfxtp_1
X_12188_ _12188_/A vssd1 vssd1 vccd1 vccd1 _12188_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18804_ _19204_/CLK _18804_/D vssd1 vssd1 vccd1 vccd1 _18804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11139_ _10976_/X _11138_/X _10988_/X vssd1 vssd1 vccd1 vccd1 _11139_/Y sky130_fd_sc_hd__o21ai_1
X_16996_ _17007_/A _17003_/C vssd1 vssd1 vccd1 vccd1 _16996_/Y sky130_fd_sc_hd__nor2_1
X_19784_ _19805_/CLK _19784_/D vssd1 vssd1 vccd1 vccd1 _19784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15947_ _19400_/Q _15238_/X _15951_/S vssd1 vssd1 vccd1 vccd1 _15948_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18735_ _19292_/CLK _18735_/D vssd1 vssd1 vccd1 vccd1 _18735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14559__A _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18051__B2 _12436_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18666_ _19952_/CLK _18666_/D vssd1 vssd1 vccd1 vccd1 _18666_/Q sky130_fd_sc_hd__dfxtp_1
X_15878_ _15878_/A vssd1 vssd1 vccd1 vccd1 _19369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17617_ _17608_/A _17610_/B _17533_/X _17613_/X _17616_/Y vssd1 vssd1 vccd1 vccd1
+ _17617_/X sky130_fd_sc_hd__o2111a_1
X_14829_ _16875_/A vssd1 vssd1 vccd1 vccd1 _18401_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18597_ _19573_/CLK _18597_/D vssd1 vssd1 vccd1 vccd1 _18597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17548_ _12673_/A _12673_/B _17976_/A vssd1 vssd1 vccd1 vccd1 _17548_/X sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_43_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18354__A2 _14476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17479_ _12328_/A _17866_/B _17488_/S vssd1 vssd1 vccd1 vccd1 _17479_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19218_ _19314_/CLK _19218_/D vssd1 vssd1 vccd1 vccd1 _19218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19149_ _19407_/CLK _19149_/D vssd1 vssd1 vccd1 vccd1 _19149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13638__A _15219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14233__S _14235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__S0 _11035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16014__A _16060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12154__A2 _12148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ _19921_/Q vssd1 vssd1 vccd1 vccd1 _09804_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18290__A1 _14501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09851__A _10392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _09735_/A vssd1 vssd1 vccd1 vccd1 _09736_/A sky130_fd_sc_hd__buf_2
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15064__S _15072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18042__A1 _19916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_153_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19720_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09666_ _10534_/A vssd1 vssd1 vccd1 vccd1 _09667_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15999__S _16001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09773_/A _09596_/X _09580_/X vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__o21a_1
XANTENNA__15800__A0 _19917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_168_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19956_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12090__A1 _19525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16356__A1 _19542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11621__A _17379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ _10510_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10510_/X sky130_fd_sc_hd__and2_1
XFILLER_128_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11490_ _11475_/A _11487_/X _11489_/X _09976_/A vssd1 vssd1 vccd1 vccd1 _11491_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ _10335_/A _10438_/Y _10440_/Y _10500_/A vssd1 vssd1 vccd1 vccd1 _10441_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10237__A _19915_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18404__A _18404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10372_ _18590_/Q _18851_/Q _18750_/Q _19085_/Q _10416_/S _09520_/A vssd1 vssd1 vccd1
+ vccd1 _10373_/B sky130_fd_sc_hd__mux4_1
XFILLER_108_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13160_ _13156_/X _13157_/X _13158_/X _12891_/X _16538_/B vssd1 vssd1 vccd1 vccd1
+ _13160_/X sky130_fd_sc_hd__o32a_1
XFILLER_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12111_ _12111_/A _12111_/B vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__xnor2_2
XFILLER_163_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13091_ _13091_/A vssd1 vssd1 vccd1 vccd1 _18473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12042_ _12042_/A _17832_/A vssd1 vssd1 vccd1 vccd1 _12104_/C sky130_fd_sc_hd__or2_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_106_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19203_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11353__B1 _11082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16850_ _19715_/Q _16845_/B _16849_/Y vssd1 vssd1 vccd1 vccd1 _19715_/D sky130_fd_sc_hd__o21a_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16292__A0 _12741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15801_ _15800_/X _19348_/Q _15801_/S vssd1 vssd1 vccd1 vccd1 _15802_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16781_ _19698_/Q _19697_/Q _16781_/C vssd1 vssd1 vccd1 vccd1 _16784_/B sky130_fd_sc_hd__and3_1
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13993_ _13993_/A vssd1 vssd1 vccd1 vccd1 _18631_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11105__B1 _10980_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18520_ _19559_/CLK _18520_/D vssd1 vssd1 vccd1 vccd1 _18520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _15732_/A vssd1 vssd1 vccd1 vccd1 _19335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12944_ _12944_/A vssd1 vssd1 vccd1 vccd1 _18441_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _19954_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _11952_/D _15662_/X _13563_/Y vssd1 vssd1 vccd1 vccd1 _15808_/A sky130_fd_sc_hd__a21o_2
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _16315_/A _12856_/X _12874_/X _17319_/B _12914_/A vssd1 vssd1 vccd1 vccd1
+ _12875_/X sky130_fd_sc_hd__o32a_1
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _17721_/A _17538_/C vssd1 vssd1 vccd1 vccd1 _17966_/A sky130_fd_sc_hd__or2_2
X_14614_ _14614_/A vssd1 vssd1 vccd1 vccd1 _18875_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18382_ input65/X vssd1 vssd1 vccd1 vccd1 _18382_/Y sky130_fd_sc_hd__clkinv_4
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _11870_/C _12088_/B _11823_/X _11977_/A vssd1 vssd1 vccd1 vccd1 _11826_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _14580_/X _19291_/Q _15600_/S vssd1 vssd1 vccd1 vccd1 _15595_/A sky130_fd_sc_hd__mux2_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17333_ _17327_/A _12610_/A _11648_/C _17331_/X _17332_/X vssd1 vssd1 vccd1 vccd1
+ _17333_/X sky130_fd_sc_hd__o311a_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14545_ _14545_/A vssd1 vssd1 vccd1 vccd1 _18850_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11757_ _11856_/S _12633_/B _11756_/Y vssd1 vssd1 vccd1 vccd1 _11849_/C sky130_fd_sc_hd__o21ai_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10708_ _10764_/A _10708_/B vssd1 vssd1 vccd1 vccd1 _10708_/Y sky130_fd_sc_hd__nor2_1
X_17264_ _17264_/A vssd1 vssd1 vccd1 vccd1 _19856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14476_ _14476_/A vssd1 vssd1 vccd1 vccd1 _16811_/A sky130_fd_sc_hd__buf_2
XFILLER_174_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11688_ _11688_/A vssd1 vssd1 vccd1 vccd1 _11928_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19003_ _19485_/CLK _19003_/D vssd1 vssd1 vccd1 vccd1 _19003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16215_ _16219_/A _16219_/C vssd1 vssd1 vccd1 vccd1 _16215_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_174_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13030__A0 _09345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13427_ _19949_/Q vssd1 vssd1 vccd1 vccd1 _13428_/A sky130_fd_sc_hd__clkbuf_2
X_10639_ _10639_/A vssd1 vssd1 vccd1 vccd1 _10639_/Y sky130_fd_sc_hd__inv_2
X_17195_ _19832_/Q _17195_/B vssd1 vssd1 vccd1 vccd1 _17195_/X sky130_fd_sc_hd__or2_1
XFILLER_155_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16146_ _16146_/A vssd1 vssd1 vccd1 vccd1 _19488_/D sky130_fd_sc_hd__clkbuf_1
X_13358_ _18488_/Q _13357_/X _13358_/S vssd1 vssd1 vccd1 vccd1 _13359_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11019__S0 _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12309_ _12309_/A vssd1 vssd1 vccd1 vccd1 _12309_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16077_ _16077_/A vssd1 vssd1 vccd1 vccd1 _19457_/D sky130_fd_sc_hd__clkbuf_1
X_13289_ _19657_/Q _12887_/A _12889_/A _19789_/Q _13288_/X vssd1 vssd1 vccd1 vccd1
+ _13289_/X sky130_fd_sc_hd__a221o_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15028_ _15028_/A vssd1 vssd1 vccd1 vccd1 _19050_/D sky130_fd_sc_hd__clkbuf_1
X_19905_ _19986_/CLK _19905_/D vssd1 vssd1 vccd1 vccd1 _19905_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13892__S _13900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19836_ _19836_/CLK _19836_/D vssd1 vssd1 vccd1 vccd1 _19836_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10242__S1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_70_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19569_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19767_ _19768_/CLK _19767_/D vssd1 vssd1 vccd1 vccd1 _19767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 io_dbus_rdata[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
X_16979_ _17007_/A _16981_/B vssd1 vssd1 vccd1 vccd1 _16979_/Y sky130_fd_sc_hd__nor2_1
X_09520_ _09520_/A vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__buf_2
XANTENNA__14833__B2 _14832_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18718_ _19564_/CLK _18718_/D vssd1 vssd1 vccd1 vccd1 _18718_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09935__S1 _09929_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19698_ _19737_/CLK _19698_/D vssd1 vssd1 vccd1 vccd1 _19698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11425__B _12667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09451_ _20049_/Q vssd1 vssd1 vccd1 vccd1 _18343_/A sky130_fd_sc_hd__clkbuf_4
X_18649_ _19464_/CLK _18649_/D vssd1 vssd1 vccd1 vccd1 _18649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_85_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19301_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09382_ _20010_/Q vssd1 vssd1 vccd1 vccd1 _12702_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18327__A2 _18291_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15848__A _15916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19407_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11583__B1 _11324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15059__S _15059_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14898__S _14900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19439_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16813__A2 _16812_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09718_ _09718_/A vssd1 vssd1 vccd1 vccd1 _09719_/A sky130_fd_sc_hd__clkbuf_2
X_10990_ _19459_/Q _19297_/Q _18706_/Q _18476_/Q _10018_/A _11225_/A vssd1 vssd1 vccd1
+ vccd1 _10991_/B sky130_fd_sc_hd__mux4_1
XFILLER_55_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09649_ _10591_/S vssd1 vssd1 vccd1 vccd1 _10496_/S sky130_fd_sc_hd__buf_2
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12663_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _12660_/Y sky130_fd_sc_hd__nor2_8
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _14477_/C vssd1 vssd1 vccd1 vccd1 _11665_/B sky130_fd_sc_hd__buf_4
XFILLER_24_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12591_ _12532_/A _12535_/A _12555_/A _12556_/Y _12579_/A vssd1 vssd1 vccd1 vccd1
+ _12618_/B sky130_fd_sc_hd__a311o_1
XANTENNA__14138__S _14142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14330_ _18777_/Q _13672_/X _14330_/S vssd1 vssd1 vccd1 vccd1 _14331_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11542_ _11550_/A _11548_/C _11540_/Y _11541_/Y vssd1 vssd1 vccd1 vccd1 _11545_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_51_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11810__A1 _11808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17957__B _17957_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ _14261_/A vssd1 vssd1 vccd1 vccd1 _18746_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11249__S0 _11057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11473_ _11473_/A _11473_/B vssd1 vssd1 vccd1 vccd1 _11473_/X sky130_fd_sc_hd__or2_1
XFILLER_109_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16000_ _16000_/A vssd1 vssd1 vccd1 vccd1 _19423_/D sky130_fd_sc_hd__clkbuf_1
X_13212_ _19903_/Q _15722_/B _13468_/S vssd1 vssd1 vccd1 vccd1 _13212_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input70_A reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10424_ _10314_/X _10415_/X _10419_/X _10423_/X _10519_/A vssd1 vssd1 vccd1 vccd1
+ _10424_/X sky130_fd_sc_hd__a311o_1
XANTENNA__09756__A _09756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14192_ _13806_/X _18716_/Q _14196_/S vssd1 vssd1 vccd1 vccd1 _14193_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12497__A2_N _12666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13143_ _19681_/Q _13342_/A _13141_/X _13142_/X vssd1 vssd1 vccd1 vccd1 _13143_/X
+ sky130_fd_sc_hd__a22o_1
X_10355_ _19472_/Q _19310_/Q _18719_/Q _18489_/Q _09651_/A _10440_/A vssd1 vssd1 vccd1
+ vccd1 _10356_/B sky130_fd_sc_hd__mux4_1
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10279_/Y _10281_/Y _10283_/Y _10285_/Y _09719_/A vssd1 vssd1 vccd1 vccd1
+ _10286_/X sky130_fd_sc_hd__o221a_1
XFILLER_112_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _19646_/Q vssd1 vssd1 vccd1 vccd1 _16617_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17951_ _17946_/X _17948_/Y _17950_/X vssd1 vssd1 vccd1 vccd1 _17951_/X sky130_fd_sc_hd__o21a_1
XFILLER_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output157_A _12424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16902_ _19732_/Q vssd1 vssd1 vccd1 vccd1 _16924_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_12025_ hold21/A _12150_/B vssd1 vssd1 vccd1 vccd1 _12037_/A sky130_fd_sc_hd__or2_1
X_17882_ _17725_/A _17883_/B _17881_/Y _17722_/A vssd1 vssd1 vccd1 vccd1 _17885_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12910__A _12989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19621_ _19762_/CLK _19621_/D vssd1 vssd1 vccd1 vccd1 _19621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16833_ _16939_/A vssd1 vssd1 vccd1 vccd1 _16833_/X sky130_fd_sc_hd__buf_2
XFILLER_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16764_ _16773_/A _16764_/B _16765_/B vssd1 vssd1 vccd1 vccd1 _19692_/D sky130_fd_sc_hd__nor3_1
X_19552_ _19552_/CLK _19552_/D vssd1 vssd1 vccd1 vccd1 _19552_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09917__S1 _09899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ _13976_/A vssd1 vssd1 vccd1 vccd1 _18623_/D sky130_fd_sc_hd__clkbuf_1
X_15715_ _15715_/A vssd1 vssd1 vccd1 vccd1 _19332_/D sky130_fd_sc_hd__clkbuf_1
X_18503_ _19852_/CLK _18503_/D vssd1 vssd1 vccd1 vccd1 _18503_/Q sky130_fd_sc_hd__dfxtp_1
X_12927_ _12914_/A _12908_/X _12880_/X _12883_/X _12926_/X vssd1 vssd1 vccd1 vccd1
+ _19771_/D sky130_fd_sc_hd__o32a_1
XFILLER_62_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16695_ _16507_/B _16692_/B _16694_/Y vssd1 vssd1 vccd1 vccd1 _19673_/D sky130_fd_sc_hd__o21a_1
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19483_ _19576_/CLK _19483_/D vssd1 vssd1 vccd1 vccd1 _19483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15646_ _15646_/A vssd1 vssd1 vccd1 vccd1 _15655_/S sky130_fd_sc_hd__buf_4
XANTENNA__17213__A _17242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18434_ _18349_/A _17138_/B _14486_/X _18433_/Y vssd1 vssd1 vccd1 vccd1 _18435_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ _14476_/A _16268_/A vssd1 vssd1 vccd1 vccd1 _17319_/B sky130_fd_sc_hd__nand2_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ _18365_/A _18365_/B vssd1 vssd1 vccd1 vccd1 _18366_/A sky130_fd_sc_hd__or2_1
X_11809_ _11809_/A vssd1 vssd1 vccd1 vccd1 _11966_/A sky130_fd_sc_hd__buf_2
X_15577_ _19284_/Q _15283_/X _15583_/S vssd1 vssd1 vccd1 vccd1 _15578_/A sky130_fd_sc_hd__mux2_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11488__S0 _09967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12789_ _13587_/A _12787_/X _12788_/Y _12903_/A _18455_/Q vssd1 vssd1 vccd1 vccd1
+ _15764_/A sky130_fd_sc_hd__a32oi_4
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17316_/A vssd1 vssd1 vccd1 vccd1 _19880_/D sky130_fd_sc_hd__clkbuf_1
X_14528_ _14528_/A vssd1 vssd1 vccd1 vccd1 _18842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18296_ _20030_/Q _18291_/X _18295_/Y _18289_/X vssd1 vssd1 vccd1 vccd1 _19998_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18190__A0 _19953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13887__S _13889_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17247_ _17247_/A _17247_/B _17247_/C _17247_/D vssd1 vssd1 vccd1 vccd1 _17304_/A
+ sky130_fd_sc_hd__or4_4
X_14459_ _14663_/A vssd1 vssd1 vccd1 vccd1 _14459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17178_ _19826_/Q _17180_/B vssd1 vssd1 vccd1 vccd1 _17178_/X sky130_fd_sc_hd__or2_1
XFILLER_127_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16129_ _16129_/A vssd1 vssd1 vccd1 vccd1 _19481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12820__A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14511__S _14513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19819_ _19852_/CLK _19819_/D vssd1 vssd1 vccd1 vccd1 _19819_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09503_ _10560_/S vssd1 vssd1 vccd1 vccd1 _10466_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17756__B1 _09464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13651__A _14605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17123__A _17123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ _20045_/Q vssd1 vssd1 vccd1 vccd1 _18333_/A sky130_fd_sc_hd__buf_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _12711_/A _12689_/B _09375_/A vssd1 vssd1 vccd1 vccd1 _13527_/B sky130_fd_sc_hd__nor3_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09296_ _09608_/A _09282_/X _09287_/X _09295_/X vssd1 vssd1 vccd1 vccd1 _09296_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13797__S _13797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09576__A _10621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12348__A2 _11771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ _11543_/A _10140_/B _10139_/X vssd1 vssd1 vccd1 vccd1 _11424_/B sky130_fd_sc_hd__or3b_1
XFILLER_161_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_165_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput170 _16458_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[6] sky130_fd_sc_hd__buf_2
XFILLER_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10071_ _18822_/Q _19157_/Q _10675_/A vssd1 vssd1 vccd1 vccd1 _10071_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10206__S1 _10196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13830_ _13830_/A vssd1 vssd1 vccd1 vccd1 _18563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ _14586_/A vssd1 vssd1 vccd1 vccd1 _13761_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10973_ _11179_/A vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__14657__A _14657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15252__S _15261_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15500_ _19250_/Q _15276_/X _15500_/S vssd1 vssd1 vccd1 vccd1 _15501_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12712_ _12837_/A _12837_/B vssd1 vssd1 vccd1 vccd1 _12995_/A sky130_fd_sc_hd__nor2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _17185_/A vssd1 vssd1 vccd1 vccd1 _16480_/X sky130_fd_sc_hd__clkbuf_4
X_13692_ _15260_/A vssd1 vssd1 vccd1 vccd1 _14637_/A sky130_fd_sc_hd__buf_2
XFILLER_44_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15431_ _14656_/X _19219_/Q _15439_/S vssd1 vssd1 vccd1 vccd1 _15432_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12036__A1 _12026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13233__A0 _19905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ _12643_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _12643_/Y sky130_fd_sc_hd__nor2_4
XFILLER_62_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18150_ _18183_/A vssd1 vssd1 vccd1 vccd1 _18159_/S sky130_fd_sc_hd__clkbuf_2
X_15362_ _15362_/A vssd1 vssd1 vccd1 vccd1 _19188_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11244__C1 _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12574_ _12574_/A vssd1 vssd1 vccd1 vccd1 _18111_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17101_ _17101_/A vssd1 vssd1 vccd1 vccd1 _17101_/X sky130_fd_sc_hd__buf_4
X_14313_ _18769_/Q _13639_/X _14319_/S vssd1 vssd1 vccd1 vccd1 _14314_/A sky130_fd_sc_hd__mux2_1
X_18081_ _17543_/X _18078_/X _18080_/Y _17794_/X vssd1 vssd1 vccd1 vccd1 _18081_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11525_ _11534_/A _11534_/B _11524_/Y vssd1 vssd1 vccd1 vccd1 _11530_/B sky130_fd_sc_hd__a21oi_1
X_15293_ _19159_/Q _15292_/X hold9/X vssd1 vssd1 vccd1 vccd1 _15294_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14392__A _14596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17032_ _19766_/Q _17033_/C _19767_/Q vssd1 vssd1 vccd1 vccd1 _17034_/B sky130_fd_sc_hd__a21oi_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09486__A _10840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14244_ _13777_/X _18739_/Q _14246_/S vssd1 vssd1 vccd1 vccd1 _14245_/A sky130_fd_sc_hd__mux2_1
X_11456_ _10052_/X _11455_/X _09706_/A vssd1 vssd1 vccd1 vccd1 _11456_/X sky130_fd_sc_hd__o21a_1
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10407_ _10407_/A _10407_/B vssd1 vssd1 vccd1 vccd1 _10407_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14175_ _14175_/A vssd1 vssd1 vccd1 vccd1 _18708_/D sky130_fd_sc_hd__clkbuf_1
X_11387_ _11387_/A _11387_/B vssd1 vssd1 vccd1 vccd1 _11387_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13126_ _13066_/X _13114_/X _13115_/Y _13125_/X vssd1 vssd1 vccd1 vccd1 _13126_/X
+ sky130_fd_sc_hd__a31o_1
X_10338_ _18783_/Q _19054_/Q _19278_/Q _19022_/Q _10337_/X _09667_/A vssd1 vssd1 vccd1
+ vccd1 _10338_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15828__A3 _15819_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18983_ _19369_/CLK _18983_/D vssd1 vssd1 vccd1 vccd1 _18983_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10770__A1 _10757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10144__B _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _18471_/Q _13056_/X _13090_/S vssd1 vssd1 vccd1 vccd1 _13058_/A sky130_fd_sc_hd__mux2_1
X_17934_ _11625_/B _17937_/A _17814_/X _17933_/Y vssd1 vssd1 vccd1 vccd1 _17934_/X
+ sky130_fd_sc_hd__o211a_1
X_10269_ _10269_/A vssd1 vssd1 vccd1 vccd1 _10269_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ _19522_/Q _11915_/A _11778_/A vssd1 vssd1 vccd1 vccd1 _12008_/X sky130_fd_sc_hd__o21a_1
XFILLER_120_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17865_ _17863_/Y _17864_/X _17865_/S vssd1 vssd1 vccd1 vccd1 _17865_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19604_ _19987_/CLK _19604_/D vssd1 vssd1 vccd1 vccd1 _19604_/Q sky130_fd_sc_hd__dfxtp_2
X_16816_ _16815_/Y _17346_/A _16816_/C _16816_/D vssd1 vssd1 vccd1 vccd1 _16832_/C
+ sky130_fd_sc_hd__and4b_4
XFILLER_54_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17796_ _17940_/A vssd1 vssd1 vccd1 vccd1 _17796_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19535_ _19988_/CLK _19535_/D vssd1 vssd1 vccd1 vccd1 _19535_/Q sky130_fd_sc_hd__dfxtp_2
X_13959_ _18616_/Q _13668_/X _13961_/S vssd1 vssd1 vccd1 vccd1 _13960_/A sky130_fd_sc_hd__mux2_1
X_16747_ _19686_/Q _16747_/B _16747_/C vssd1 vssd1 vccd1 vccd1 _16748_/C sky130_fd_sc_hd__and3_1
XFILLER_59_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13471__A _15283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19466_ _19560_/CLK _19466_/D vssd1 vssd1 vccd1 vccd1 _19466_/Q sky130_fd_sc_hd__dfxtp_1
X_16678_ _16678_/A vssd1 vssd1 vccd1 vccd1 _16898_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10381__S0 _10416_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18417_ _18426_/A _18417_/B vssd1 vssd1 vccd1 vccd1 _20046_/D sky130_fd_sc_hd__nor2_1
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15629_ _14631_/X _19307_/Q _15633_/S vssd1 vssd1 vccd1 vccd1 _15630_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19397_ _19514_/CLK _19397_/D vssd1 vssd1 vccd1 vccd1 _19397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18348_ _16808_/B _18302_/B _18347_/X _18341_/X vssd1 vssd1 vccd1 vccd1 _20019_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18279_ _18279_/A _18311_/B vssd1 vssd1 vccd1 vccd1 _18279_/X sky130_fd_sc_hd__or2_1
XANTENNA__10684__S1 _10682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12815__A _13578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput50 io_ibus_inst[24] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
Xinput61 io_ibus_inst[5] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10335__A _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09983_ _09983_/A vssd1 vssd1 vccd1 vccd1 _10812_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_88_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15337__S _15345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13646__A _15225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10070__A _11482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13463__B1 _13099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15072__S _15072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__S0 _10416_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09417_ input70/X _17346_/B vssd1 vssd1 vccd1 vccd1 _18138_/A sky130_fd_sc_hd__nor2_2
XANTENNA__12018__A1 _10869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_91_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11226__C1 _10899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09348_ _19888_/Q vssd1 vssd1 vccd1 vccd1 _09349_/A sky130_fd_sc_hd__inv_2
XANTENNA__10124__S0 _10753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09279_ _20036_/Q vssd1 vssd1 vccd1 vccd1 _09608_/A sky130_fd_sc_hd__buf_2
XFILLER_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11310_ _18763_/Q _19034_/Q _19258_/Q _19002_/Q _11114_/S _11260_/A vssd1 vssd1 vccd1
+ vccd1 _11310_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12290_ _12365_/D _12395_/S _12290_/C vssd1 vssd1 vccd1 vccd1 _12290_/X sky130_fd_sc_hd__and3b_1
XFILLER_147_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11241_ _11250_/A _11241_/B vssd1 vssd1 vccd1 vccd1 _11241_/X sky130_fd_sc_hd__or2_1
XANTENNA__10427__S1 _10291_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18412__A _18412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11172_ _11280_/S vssd1 vssd1 vccd1 vccd1 _11329_/S sky130_fd_sc_hd__buf_2
XFILLER_122_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10123_ _09706_/A _10107_/Y _10115_/X _10122_/Y _09738_/A vssd1 vssd1 vccd1 vccd1
+ _10123_/X sky130_fd_sc_hd__o311a_1
XANTENNA__17028__A _17066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15980_ _19415_/Q _15286_/X _15984_/S vssd1 vssd1 vccd1 vccd1 _15981_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A io_dbus_valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10054_ _10054_/A vssd1 vssd1 vccd1 vccd1 _10054_/X sky130_fd_sc_hd__buf_4
X_14931_ _19007_/Q _14388_/X _14939_/S vssd1 vssd1 vccd1 vccd1 _14932_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13990__S _13994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17650_ _17647_/X _17648_/X _17800_/S vssd1 vssd1 vccd1 vccd1 _17651_/A sky130_fd_sc_hd__mux2_1
X_14862_ _14862_/A vssd1 vssd1 vccd1 vccd1 _18976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13813_ _13812_/X _18558_/Q _13813_/S vssd1 vssd1 vccd1 vccd1 _13814_/A sky130_fd_sc_hd__mux2_1
X_16601_ _16631_/A _16601_/B vssd1 vssd1 vccd1 vccd1 _16601_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17581_ _17579_/X _17580_/X _17581_/S vssd1 vssd1 vccd1 vccd1 _17581_/X sky130_fd_sc_hd__mux2_1
X_14793_ _18950_/Q _14427_/X _14797_/S vssd1 vssd1 vccd1 vccd1 _14794_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19320_ _19482_/CLK _19320_/D vssd1 vssd1 vccd1 vccd1 _19320_/Q sky130_fd_sc_hd__dfxtp_1
X_16532_ _19617_/Q _16528_/C _16531_/Y vssd1 vssd1 vccd1 vccd1 _19617_/D sky130_fd_sc_hd__o21a_1
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13744_ _18538_/Q _13743_/X _13744_/S vssd1 vssd1 vccd1 vccd1 _13745_/A sky130_fd_sc_hd__mux2_1
X_10956_ _18642_/Q _19233_/Q _19395_/Q _18610_/Q _10893_/X _09512_/A vssd1 vssd1 vccd1
+ vccd1 _10956_/X sky130_fd_sc_hd__mux4_1
X_19251_ _19569_/CLK _19251_/D vssd1 vssd1 vccd1 vccd1 _19251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16463_ _12037_/A _12037_/B _16455_/X vssd1 vssd1 vccd1 vccd1 _19587_/D sky130_fd_sc_hd__a21o_1
X_13675_ _15247_/A vssd1 vssd1 vccd1 vccd1 _14624_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13206__B1 _13205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887_ _11489_/A _10887_/B vssd1 vssd1 vccd1 vccd1 _10887_/X sky130_fd_sc_hd__or2_1
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ _15414_/A vssd1 vssd1 vccd1 vccd1 _19211_/D sky130_fd_sc_hd__clkbuf_1
X_18202_ _18202_/A vssd1 vssd1 vccd1 vccd1 _19957_/D sky130_fd_sc_hd__clkbuf_1
X_19182_ _19409_/CLK _19182_/D vssd1 vssd1 vccd1 vccd1 _19182_/Q sky130_fd_sc_hd__dfxtp_1
X_12626_ _17240_/A _12588_/B _19848_/Q vssd1 vssd1 vccd1 vccd1 _12626_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_169_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16394_ _16394_/A vssd1 vssd1 vccd1 vccd1 _19555_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10139__B _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18133_ _18133_/A vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__clkbuf_1
X_15345_ _19181_/Q _15260_/X _15345_/S vssd1 vssd1 vccd1 vccd1 _15346_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _12555_/Y _12556_/Y _12532_/A _12535_/A vssd1 vssd1 vccd1 vccd1 _12559_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10666__S1 _10665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12635__A _12635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13509__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ _10039_/A _11507_/X _10056_/A vssd1 vssd1 vccd1 vccd1 _11508_/Y sky130_fd_sc_hd__o21ai_1
X_18064_ _19918_/Q _18019_/X _18063_/X vssd1 vssd1 vccd1 vccd1 _19918_/D sky130_fd_sc_hd__o21a_1
XFILLER_172_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15276_ _15276_/A vssd1 vssd1 vccd1 vccd1 _15276_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12488_ _12485_/Y _12487_/Y _12583_/S vssd1 vssd1 vccd1 vccd1 _12488_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17015_ _17073_/A vssd1 vssd1 vccd1 vccd1 _17066_/A sky130_fd_sc_hd__buf_2
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14227_ _13746_/X _18731_/Q _14235_/S vssd1 vssd1 vccd1 vccd1 _14228_/A sky130_fd_sc_hd__mux2_1
X_11439_ _19513_/Q _18925_/Q _18962_/Q _18536_/Q _10690_/X _10691_/X vssd1 vssd1 vccd1
+ vccd1 _11440_/B sky130_fd_sc_hd__mux4_1
XFILLER_99_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09944__A _19917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14158_ _14158_/A vssd1 vssd1 vccd1 vccd1 _18700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _15215_/A vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ _19666_/CLK _18966_/D vssd1 vssd1 vccd1 vccd1 _18966_/Q sky130_fd_sc_hd__dfxtp_2
X_14089_ _14146_/S vssd1 vssd1 vccd1 vccd1 _14098_/S sky130_fd_sc_hd__buf_2
XFILLER_26_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _17917_/A _17917_/B vssd1 vssd1 vccd1 vccd1 _17919_/C sky130_fd_sc_hd__nor2_1
XANTENNA__14996__S _15000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18897_ _19485_/CLK _18897_/D vssd1 vssd1 vccd1 vccd1 _18897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17848_ _17600_/X _17742_/A _17632_/X vssd1 vssd1 vccd1 vccd1 _17848_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_94_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13445__B1 _13099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17779_ _11940_/Y _17755_/X _17777_/X _17778_/X vssd1 vssd1 vccd1 vccd1 _17779_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19518_ _19831_/CLK _19518_/D vssd1 vssd1 vccd1 vccd1 _19518_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_clkbuf_leaf_113_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19449_ _19449_/CLK _19449_/D vssd1 vssd1 vccd1 vccd1 _19449_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15620__S _15622_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _09215_/A vssd1 vssd1 vccd1 vccd1 _09202_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__17401__A _17542_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18136__A0 _16219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10106__S0 _11449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12545__A _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10065__A _10065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11931__A0 _19963_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13376__A _15263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_38_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _11475_/A vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__buf_2
XFILLER_103_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09897_ _10373_/A vssd1 vssd1 vccd1 vccd1 _10254_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09352__A1 _19894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15591__A _15659_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _11378_/A _10810_/B vssd1 vssd1 vccd1 vccd1 _10810_/X sky130_fd_sc_hd__or2_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11790_ _11790_/A _11790_/B vssd1 vssd1 vccd1 vccd1 _11792_/B sky130_fd_sc_hd__or2_2
XFILLER_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ _11362_/A _10741_/B vssd1 vssd1 vccd1 vccd1 _10741_/X sky130_fd_sc_hd__or2_1
XFILLER_14_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10670__B1 _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13460_ _16347_/A _13460_/B vssd1 vssd1 vccd1 vccd1 _13460_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10672_ _10672_/A _12650_/A vssd1 vssd1 vccd1 vccd1 _10673_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12411_ _12411_/A _12411_/B vssd1 vssd1 vccd1 vccd1 _12413_/A sky130_fd_sc_hd__nor2_1
XFILLER_166_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14146__S _14146_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ input14/X _13353_/X _13354_/X vssd1 vssd1 vccd1 vccd1 _13391_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__12455__A _12455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15130_ _15130_/A vssd1 vssd1 vccd1 vccd1 _19096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12342_ _11745_/X _12336_/Y _12341_/X vssd1 vssd1 vccd1 vccd1 _12342_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15061_ _15061_/A _18297_/A _15373_/A _15373_/B vssd1 vssd1 vccd1 vccd1 _15118_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_142_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12273_ _17389_/A _12300_/B vssd1 vssd1 vccd1 vccd1 _12274_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14012_ _14012_/A vssd1 vssd1 vccd1 vccd1 _18638_/D sky130_fd_sc_hd__clkbuf_1
X_11224_ _18798_/Q _19133_/Q _11224_/S vssd1 vssd1 vccd1 vccd1 _11225_/B sky130_fd_sc_hd__mux2_1
XFILLER_122_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10725__A1 _09748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12902__B _18460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__B2 _10724_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18820_ _19287_/CLK _18820_/D vssd1 vssd1 vccd1 vccd1 _18820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11155_ _11141_/A _11154_/X _09703_/A vssd1 vssd1 vccd1 vccd1 _11155_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10703__A _10703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10106_ _19125_/Q _18891_/Q _19573_/Q _19221_/Q _11449_/S _10718_/A vssd1 vssd1 vccd1
+ vccd1 _10107_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16861__B1 _16860_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18751_ _19565_/CLK _18751_/D vssd1 vssd1 vccd1 vccd1 _18751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11518__B _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15963_ _15963_/A vssd1 vssd1 vccd1 vccd1 _19407_/D sky130_fd_sc_hd__clkbuf_1
X_11086_ _10914_/X _11084_/Y _11085_/Y _09659_/A vssd1 vssd1 vccd1 vccd1 _11086_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17702_ _17702_/A _17702_/B vssd1 vssd1 vccd1 vccd1 _17702_/Y sky130_fd_sc_hd__nor2_1
X_10037_ _10037_/A vssd1 vssd1 vccd1 vccd1 _10037_/X sky130_fd_sc_hd__buf_4
X_14914_ _14914_/A vssd1 vssd1 vccd1 vccd1 _19000_/D sky130_fd_sc_hd__clkbuf_1
X_15894_ _15894_/A vssd1 vssd1 vccd1 vccd1 _19376_/D sky130_fd_sc_hd__clkbuf_1
X_18682_ _19049_/CLK _18682_/D vssd1 vssd1 vccd1 vccd1 _18682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11150__A1 _10024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17633_ _17627_/X _17906_/A _17632_/X vssd1 vssd1 vccd1 vccd1 _17633_/Y sky130_fd_sc_hd__a21oi_1
X_14845_ _15445_/B _15990_/B vssd1 vssd1 vccd1 vccd1 _14902_/A sky130_fd_sc_hd__or2_4
XANTENNA__10849__S _10849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17564_ _17432_/X _17420_/X _17565_/S vssd1 vssd1 vccd1 vccd1 _17564_/X sky130_fd_sc_hd__mux2_1
X_14776_ _14776_/A vssd1 vssd1 vccd1 vccd1 _18942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11988_ _12069_/A _12643_/A _12039_/C _20049_/Q vssd1 vssd1 vccd1 vccd1 _12042_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12349__B _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19303_ _19369_/CLK _19303_/D vssd1 vssd1 vccd1 vccd1 _19303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13727_ _14663_/A vssd1 vssd1 vccd1 vccd1 _13727_/X sky130_fd_sc_hd__clkbuf_2
X_16515_ _16518_/B _16518_/C _12908_/X vssd1 vssd1 vccd1 vccd1 _16515_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10939_ _11191_/S vssd1 vssd1 vccd1 vccd1 _11237_/S sky130_fd_sc_hd__buf_4
X_17495_ _12432_/A _17792_/B _17504_/S vssd1 vssd1 vccd1 vccd1 _17495_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18317__A _18341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19234_ _19490_/CLK _19234_/D vssd1 vssd1 vccd1 vccd1 _19234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13658_ _13658_/A vssd1 vssd1 vccd1 vccd1 _18517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16446_ _17319_/A vssd1 vssd1 vccd1 vccd1 _17185_/A sky130_fd_sc_hd__clkbuf_2
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _17391_/B _12609_/B _12609_/C _12609_/D vssd1 vssd1 vccd1 vccd1 _12611_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__12402__A1 _17338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16377_ _16377_/A vssd1 vssd1 vccd1 vccd1 _19547_/D sky130_fd_sc_hd__clkbuf_1
X_19165_ _19391_/CLK _19165_/D vssd1 vssd1 vccd1 vccd1 _19165_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09803__C1 _09719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13589_ _15783_/A _18439_/Q vssd1 vssd1 vccd1 vccd1 _13589_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15328_ _19173_/Q _15235_/X _15334_/S vssd1 vssd1 vccd1 vccd1 _15329_/A sky130_fd_sc_hd__mux2_1
X_18116_ _12579_/X _17755_/A _18115_/X _12951_/A vssd1 vssd1 vccd1 vccd1 _18116_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_144_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09377__C _12888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19096_ _19299_/CLK _19096_/D vssd1 vssd1 vccd1 vccd1 _19096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15259_ _15259_/A vssd1 vssd1 vccd1 vccd1 _19148_/D sky130_fd_sc_hd__clkbuf_1
X_18047_ _17791_/X _18043_/Y _18046_/Y vssd1 vssd1 vccd1 vccd1 _18047_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_160_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09820_ _09820_/A vssd1 vssd1 vccd1 vccd1 _09820_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19998_ _19998_/CLK _19998_/D vssd1 vssd1 vccd1 vccd1 _19998_/Q sky130_fd_sc_hd__dfxtp_2
X_09751_ _09751_/A _09751_/B _09751_/C vssd1 vssd1 vccd1 vccd1 _09752_/A sky130_fd_sc_hd__or3_4
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18949_ _19500_/CLK _18949_/D vssd1 vssd1 vccd1 vccd1 _18949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09682_ _10548_/A vssd1 vssd1 vccd1 vccd1 _10407_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10327__S0 _10325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10101__C1 _10621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14755__A _14823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16181__S _16189_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14490__A _16678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09584__A _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11904__A0 _19962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10802__S1 _10682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09949_ _11491_/A vssd1 vssd1 vccd1 vccd1 _10834_/A sky130_fd_sc_hd__buf_2
XFILLER_77_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12960_ _18450_/Q _12959_/X _11406_/A _12954_/X vssd1 vssd1 vccd1 vccd1 _18450_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16210__A _16299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11911_ _11911_/A vssd1 vssd1 vccd1 vccd1 _12153_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _13204_/A vssd1 vssd1 vccd1 vccd1 _12891_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14630_/A vssd1 vssd1 vccd1 vccd1 _18880_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _19820_/Q _11842_/B vssd1 vssd1 vccd1 vccd1 _11843_/C sky130_fd_sc_hd__xnor2_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10318__S0 _09505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14561_/A vssd1 vssd1 vccd1 vccd1 _18857_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__A3 _10236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ _19813_/Q _19808_/Q _11772_/Y _11837_/A vssd1 vssd1 vccd1 vccd1 _11773_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16300_ _16300_/A vssd1 vssd1 vccd1 vccd1 _16300_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _19954_/Q _13512_/B vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__and2_1
X_10724_ _19905_/Q vssd1 vssd1 vccd1 vccd1 _10724_/Y sky130_fd_sc_hd__inv_2
X_17280_ _17191_/Y _19864_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17281_/A sky130_fd_sc_hd__mux2_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ input48/X vssd1 vssd1 vccd1 vccd1 _14492_/Y sky130_fd_sc_hd__inv_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ _16231_/A vssd1 vssd1 vccd1 vccd1 _19519_/D sky130_fd_sc_hd__clkbuf_1
X_13443_ _19731_/Q vssd1 vssd1 vccd1 vccd1 _16924_/C sky130_fd_sc_hd__clkbuf_2
X_10655_ _10655_/A vssd1 vssd1 vccd1 vccd1 _10655_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17976__A _17976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16162_ _16162_/A vssd1 vssd1 vccd1 vccd1 _19495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13374_ input13/X _13353_/X _13354_/X vssd1 vssd1 vccd1 vccd1 _13374_/Y sky130_fd_sc_hd__a21oi_2
X_10586_ _10579_/Y _10581_/Y _10583_/Y _10585_/Y _09718_/A vssd1 vssd1 vccd1 vccd1
+ _10586_/X sky130_fd_sc_hd__o221a_1
XFILLER_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15113_ _15113_/A vssd1 vssd1 vccd1 vccd1 _19088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12325_ _12573_/S vssd1 vssd1 vccd1 vccd1 _12528_/S sky130_fd_sc_hd__buf_2
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16091__S _16095_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16093_ _13259_/X _19465_/Q _16095_/S vssd1 vssd1 vccd1 vccd1 _16094_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12913__A _12992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15044_ _19058_/Q _14449_/X _15044_/S vssd1 vssd1 vccd1 vccd1 _15045_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09494__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19921_ _19986_/CLK _19921_/D vssd1 vssd1 vccd1 vccd1 _19921_/Q sky130_fd_sc_hd__dfxtp_4
X_12256_ _12256_/A _17445_/A vssd1 vssd1 vccd1 vccd1 _12259_/A sky130_fd_sc_hd__xor2_4
XFILLER_141_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12632__B _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11207_ _11315_/A _11207_/B vssd1 vssd1 vccd1 vccd1 _11207_/X sky130_fd_sc_hd__or2_1
XANTENNA__18284__C1 _17243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19852_ _19852_/CLK _19852_/D vssd1 vssd1 vccd1 vccd1 _19852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12187_ hold18/A _11920_/X _12182_/X _12186_/X vssd1 vssd1 vccd1 vccd1 _16471_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_68_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16834__B1 _16833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18803_ _19493_/CLK _18803_/D vssd1 vssd1 vccd1 vccd1 _18803_/Q sky130_fd_sc_hd__dfxtp_1
X_11138_ _19488_/Q _18900_/Q _18937_/Q _18511_/Q _10017_/A _10917_/A vssd1 vssd1 vccd1
+ vccd1 _11138_/X sky130_fd_sc_hd__mux4_1
X_19783_ _19783_/CLK _19783_/D vssd1 vssd1 vccd1 vccd1 _19783_/Q sky130_fd_sc_hd__dfxtp_1
X_16995_ _17005_/D vssd1 vssd1 vccd1 vccd1 _17003_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15435__S _15439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18734_ _18836_/CLK _18734_/D vssd1 vssd1 vccd1 vccd1 _18734_/Q sky130_fd_sc_hd__dfxtp_1
X_15946_ _15946_/A vssd1 vssd1 vccd1 vccd1 _19399_/D sky130_fd_sc_hd__clkbuf_1
X_11069_ _18968_/Q vssd1 vssd1 vccd1 vccd1 _11069_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11123__A1 _10875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10557__S0 _10560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18665_ _19418_/CLK _18665_/D vssd1 vssd1 vccd1 vccd1 _18665_/Q sky130_fd_sc_hd__dfxtp_1
X_15877_ _13259_/X _19369_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15878_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17616_ _17616_/A _17616_/B vssd1 vssd1 vccd1 vccd1 _17616_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14828_ _14828_/A _18402_/B vssd1 vssd1 vccd1 vccd1 _18965_/D sky130_fd_sc_hd__nor2_4
X_18596_ _19571_/CLK _18596_/D vssd1 vssd1 vccd1 vccd1 _18596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12623__A1 _12395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17547_ _17917_/A vssd1 vssd1 vccd1 vccd1 _17976_/A sky130_fd_sc_hd__buf_2
X_14759_ _14759_/A vssd1 vssd1 vccd1 vccd1 _18934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10634__B1 _09577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09669__A _09927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17478_ _17507_/S vssd1 vssd1 vccd1 vccd1 _17488_/S sky130_fd_sc_hd__buf_2
XFILLER_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19217_ _19313_/CLK _19217_/D vssd1 vssd1 vccd1 vccd1 _19217_/Q sky130_fd_sc_hd__dfxtp_1
X_16429_ _13453_/X _19571_/Q _16437_/S vssd1 vssd1 vccd1 vccd1 _16430_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10608__A _10824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19148_ _19406_/CLK _19148_/D vssd1 vssd1 vccd1 vccd1 _19148_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11285__S1 _10978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19079_ _19559_/CLK _19079_/D vssd1 vssd1 vccd1 vccd1 _19079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11037__S1 _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17617__A2 _17610_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09803_ _09796_/Y _09798_/Y _09800_/Y _09802_/Y _09719_/X vssd1 vssd1 vccd1 vccd1
+ _09803_/X sky130_fd_sc_hd__o221a_1
XFILLER_141_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15345__S _15345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13654__A _15231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _18831_/Q vssd1 vssd1 vccd1 vccd1 _09735_/A sky130_fd_sc_hd__inv_2
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09665_ _09665_/A vssd1 vssd1 vccd1 vccd1 _10534_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17250__A0 _13572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09596_ _19483_/Q _19321_/Q _18730_/Q _18500_/Q _09542_/S _09526_/X vssd1 vssd1 vccd1
+ vccd1 _09596_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16176__S _16178_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09579__A _09826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10440_ _10440_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10440_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ _10380_/A _10366_/X _10368_/X _10370_/X vssd1 vssd1 vccd1 vccd1 _10371_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12110_ _12055_/A _12055_/B _12083_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _12111_/B
+ sky130_fd_sc_hd__a31o_2
X_13090_ _18473_/Q _13089_/X _13090_/S vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12041_ _17853_/A vssd1 vssd1 vccd1 vccd1 _12045_/A sky130_fd_sc_hd__inv_2
XFILLER_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11353__A1 _10961_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__B2 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15255__S _15261_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15800_ _19917_/Q _15799_/Y _15800_/S vssd1 vssd1 vccd1 vccd1 _15800_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13992_ _18631_/Q _13731_/X _13994_/S vssd1 vssd1 vccd1 vccd1 _13993_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16780_ _19697_/Q _16781_/C _19698_/Q vssd1 vssd1 vccd1 vccd1 _16782_/B sky130_fd_sc_hd__a21oi_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ _15730_/X _19335_/Q _15747_/S vssd1 vssd1 vccd1 vccd1 _15732_/A sky130_fd_sc_hd__mux2_1
X_12943_ _18441_/Q _12942_/X _17808_/S vssd1 vssd1 vccd1 vccd1 _12944_/A sky130_fd_sc_hd__mux2_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16875__A _16875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10864__B1 _09706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18450_ _19954_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _15662_/A _15662_/B _13562_/B vssd1 vssd1 vccd1 vccd1 _15662_/X sky130_fd_sc_hd__or3b_1
X_12874_ _12735_/X _12872_/X _12873_/Y _12853_/X _18449_/Q vssd1 vssd1 vccd1 vccd1
+ _12874_/X sky130_fd_sc_hd__a32o_4
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17542_/D _17465_/S vssd1 vssd1 vccd1 vccd1 _17538_/C sky130_fd_sc_hd__or2b_1
X_14613_ _14612_/X _18875_/Q _14622_/S vssd1 vssd1 vccd1 vccd1 _14614_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11825_ _11825_/A vssd1 vssd1 vccd1 vccd1 _11977_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15593_ _15593_/A vssd1 vssd1 vccd1 vccd1 _19290_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output102_A _12024_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18381_ _18401_/A vssd1 vssd1 vccd1 vccd1 _18396_/A sky130_fd_sc_hd__buf_2
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14395__A _14599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12908__A _18281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _13809_/X _18850_/Q _14546_/S vssd1 vssd1 vccd1 vccd1 _14545_/A sky130_fd_sc_hd__mux2_1
X_17332_ _12610_/B _09426_/B _11638_/A _12610_/A vssd1 vssd1 vccd1 vccd1 _17332_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _20030_/Q _11854_/B _11894_/A _12320_/B _11755_/X vssd1 vssd1 vccd1 vccd1
+ _11756_/Y sky130_fd_sc_hd__o2111ai_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10707_ _19110_/Q _18876_/Q _19558_/Q _19206_/Q _10644_/X _10645_/X vssd1 vssd1 vccd1
+ vccd1 _10708_/B sky130_fd_sc_hd__mux4_1
X_17263_ _17166_/Y _19856_/Q _17269_/S vssd1 vssd1 vccd1 vccd1 _17264_/A sky130_fd_sc_hd__mux2_1
X_14475_ _18404_/A vssd1 vssd1 vccd1 vccd1 _17041_/B sky130_fd_sc_hd__buf_4
XFILLER_174_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11687_ _11901_/A _11901_/B _17397_/B _11901_/D vssd1 vssd1 vccd1 vccd1 _11688_/A
+ sky130_fd_sc_hd__nor4_2
XFILLER_128_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19002_ _19484_/CLK _19002_/D vssd1 vssd1 vccd1 vccd1 _19002_/Q sky130_fd_sc_hd__dfxtp_1
X_16214_ _16206_/A _19322_/Q vssd1 vssd1 vccd1 vccd1 _16219_/C sky130_fd_sc_hd__nand2b_1
X_13426_ input17/X _13318_/X _13354_/A vssd1 vssd1 vccd1 vccd1 _13432_/A sky130_fd_sc_hd__a21o_1
X_10638_ _18681_/Q _19176_/Q _11386_/S vssd1 vssd1 vccd1 vccd1 _10639_/A sky130_fd_sc_hd__mux2_1
X_17194_ _17194_/A vssd1 vssd1 vccd1 vccd1 _17194_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16145_ _19488_/Q _14589_/A _16145_/S vssd1 vssd1 vccd1 vccd1 _16146_/A sky130_fd_sc_hd__mux2_1
X_13357_ _15260_/A vssd1 vssd1 vccd1 vccd1 _13357_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10569_ _10569_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10569_/X sky130_fd_sc_hd__or2_1
XANTENNA__12643__A _12643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_clock _19998_/CLK vssd1 vssd1 vccd1 vccd1 _19892_/CLK sky130_fd_sc_hd__clkbuf_16
X_12308_ _12308_/A _12308_/B vssd1 vssd1 vccd1 vccd1 _12309_/A sky130_fd_sc_hd__xnor2_1
XFILLER_114_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16076_ _13109_/X _19457_/Q _16084_/S vssd1 vssd1 vccd1 vccd1 _16077_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13288_ _19721_/Q _13144_/S _12723_/A _19689_/Q _13287_/X vssd1 vssd1 vccd1 vccd1
+ _13288_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11019__S1 _10083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15027_ _19050_/Q _14424_/X _15033_/S vssd1 vssd1 vccd1 vccd1 _15028_/A sky130_fd_sc_hd__mux2_1
X_19904_ _19906_/CLK _19904_/D vssd1 vssd1 vccd1 vccd1 _19904_/Q sky130_fd_sc_hd__dfxtp_4
X_12239_ _12240_/B _12240_/C _16474_/A vssd1 vssd1 vccd1 vccd1 _12241_/B sky130_fd_sc_hd__a21oi_1
XFILLER_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19835_ _19836_/CLK _19835_/D vssd1 vssd1 vccd1 vccd1 _19835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17480__A0 _12356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19766_ _19768_/CLK _19766_/D vssd1 vssd1 vccd1 vccd1 _19766_/Q sky130_fd_sc_hd__dfxtp_1
X_16978_ _19751_/Q _19750_/Q _16978_/C vssd1 vssd1 vccd1 vccd1 _16981_/B sky130_fd_sc_hd__and3_1
Xinput4 io_dbus_rdata[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
XFILLER_65_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18717_ _19308_/CLK _18717_/D vssd1 vssd1 vccd1 vccd1 _18717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15929_ _19392_/Q _15212_/X _15929_/S vssd1 vssd1 vccd1 vccd1 _15930_/A sky130_fd_sc_hd__mux2_1
X_19697_ _19737_/CLK _19697_/D vssd1 vssd1 vccd1 vccd1 _19697_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12844__B2 _19525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16785__A _16818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09450_ _20050_/Q vssd1 vssd1 vccd1 vccd1 _17338_/A sky130_fd_sc_hd__clkbuf_4
X_18648_ _18845_/CLK _18648_/D vssd1 vssd1 vccd1 vccd1 _18648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09381_ _09398_/B vssd1 vssd1 vccd1 vccd1 _13136_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14509__S _14513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18579_ _19074_/CLK _18579_/D vssd1 vssd1 vccd1 vccd1 _18579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12818__A _17247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14244__S _14246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16025__A _16047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12553__A _12553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11583__A1 _11302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11583__B2 _12631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10769__S0 _11451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13088__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10801__A _10805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13088__B2 _13007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ _09717_/A vssd1 vssd1 vccd1 vccd1 _09718_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09648_ _10589_/S vssd1 vssd1 vccd1 vccd1 _10591_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_43_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15785__A0 _19914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _09826_/A vssd1 vssd1 vccd1 vccd1 _09580_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12728__A _12888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17918__A_N _17914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_161_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11610_ _11619_/A _17394_/B vssd1 vssd1 vccd1 vccd1 _14477_/C sky130_fd_sc_hd__nand2_1
XFILLER_24_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12590_ _19608_/Q _12537_/X _12585_/X _12589_/X vssd1 vssd1 vccd1 vccd1 _12590_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11541_ _11541_/A vssd1 vssd1 vccd1 vccd1 _11541_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14260_ _13799_/X _18746_/Q _14268_/S vssd1 vssd1 vccd1 vccd1 _14261_/A sky130_fd_sc_hd__mux2_1
X_11472_ _19386_/Q _19000_/Q _19450_/Q _18569_/Q _09532_/A _09985_/A vssd1 vssd1 vccd1
+ vccd1 _11473_/B sky130_fd_sc_hd__mux4_1
XFILLER_13_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11249__S1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ _16636_/B _13116_/X _13117_/X _17070_/B _13210_/X vssd1 vssd1 vccd1 vccd1
+ _15722_/B sky130_fd_sc_hd__a221o_2
X_10423_ _10426_/A _10420_/X _10422_/X _10307_/X vssd1 vssd1 vccd1 vccd1 _10423_/X
+ sky130_fd_sc_hd__o211a_1
X_14191_ _14191_/A vssd1 vssd1 vccd1 vccd1 _18715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13142_ _19617_/Q _13142_/B vssd1 vssd1 vccd1 vccd1 _13142_/X sky130_fd_sc_hd__or2_1
XANTENNA_input63_A io_ibus_inst[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10354_ _10534_/A vssd1 vssd1 vccd1 vccd1 _10440_/A sky130_fd_sc_hd__buf_2
XFILLER_151_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17973__B _17973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _16219_/B _13094_/C vssd1 vssd1 vccd1 vccd1 _13073_/X sky130_fd_sc_hd__xor2_1
X_17950_ _18000_/A _17947_/X _17949_/X _17533_/A vssd1 vssd1 vccd1 vccd1 _17950_/X
+ sky130_fd_sc_hd__o211a_1
X_10285_ _10264_/A _10284_/X _09711_/A vssd1 vssd1 vccd1 vccd1 _10285_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16901_ _16919_/A _16901_/B _16909_/D vssd1 vssd1 vccd1 vccd1 _19731_/D sky130_fd_sc_hd__nor3_1
X_12024_ _12024_/A vssd1 vssd1 vccd1 vccd1 _12024_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_86_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17881_ _17998_/A _17881_/B vssd1 vssd1 vccd1 vccd1 _17881_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13294__A _13454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19620_ _19620_/CLK _19620_/D vssd1 vssd1 vccd1 vccd1 _19620_/Q sky130_fd_sc_hd__dfxtp_1
X_16832_ _19709_/Q _19708_/Q _16832_/C _16863_/D vssd1 vssd1 vccd1 vccd1 _16848_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18006__A2 _09464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19551_ _19551_/CLK _19551_/D vssd1 vssd1 vccd1 vccd1 _19551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16763_ _19692_/Q _19691_/Q _16763_/C vssd1 vssd1 vccd1 vccd1 _16765_/B sky130_fd_sc_hd__and3_1
XFILLER_76_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13975_ _18623_/Q _13697_/X _13983_/S vssd1 vssd1 vccd1 vccd1 _13976_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18502_ _19852_/CLK _18502_/D vssd1 vssd1 vccd1 vccd1 _18502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15714_ _15713_/X _19332_/Q _15720_/S vssd1 vssd1 vccd1 vccd1 _15715_/A sky130_fd_sc_hd__mux2_1
X_19482_ _19482_/CLK _19482_/D vssd1 vssd1 vccd1 vccd1 _19482_/Q sky130_fd_sc_hd__dfxtp_1
X_12926_ _19773_/Q _14752_/B _12909_/X _12925_/Y vssd1 vssd1 vccd1 vccd1 _12926_/X
+ sky130_fd_sc_hd__o22a_1
X_16694_ _16507_/B _16692_/B _16667_/X vssd1 vssd1 vccd1 vccd1 _16694_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18433_ input58/X vssd1 vssd1 vccd1 vccd1 _18433_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15645_ _15645_/A vssd1 vssd1 vccd1 vccd1 _19314_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _12857_/A vssd1 vssd1 vccd1 vccd1 _14476_/A sky130_fd_sc_hd__buf_2
XFILLER_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18364_ _12606_/D _14476_/A _18414_/A input60/X vssd1 vssd1 vccd1 vccd1 _18365_/B
+ sky130_fd_sc_hd__o22a_1
X_11808_ _09614_/A _11244_/X _11253_/X _09621_/A _19896_/Q vssd1 vssd1 vccd1 vccd1
+ _11808_/X sky130_fd_sc_hd__a32o_4
X_15576_ _15576_/A vssd1 vssd1 vccd1 vccd1 _19283_/D sky130_fd_sc_hd__clkbuf_1
X_12788_ _15702_/A _18455_/Q vssd1 vssd1 vccd1 vccd1 _12788_/Y sky130_fd_sc_hd__nand2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _15839_/X _19880_/Q _17317_/S vssd1 vssd1 vccd1 vccd1 _17316_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14527_ _13783_/X _18842_/Q _14535_/S vssd1 vssd1 vccd1 vccd1 _14528_/A sky130_fd_sc_hd__mux2_1
X_11739_ _11739_/A _12674_/A vssd1 vssd1 vccd1 vccd1 _11740_/A sky130_fd_sc_hd__xnor2_4
X_18295_ _18295_/A _18326_/B vssd1 vssd1 vccd1 vccd1 _18295_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17246_ _17246_/A vssd1 vssd1 vccd1 vccd1 _19849_/D sky130_fd_sc_hd__clkbuf_1
X_14458_ _14458_/A vssd1 vssd1 vccd1 vccd1 _18821_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13409_ _13337_/X _13408_/X _13351_/X vssd1 vssd1 vccd1 vccd1 _13409_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__14064__S _14068_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17177_ _17175_/Y _17167_/X _17176_/X _17171_/X vssd1 vssd1 vccd1 vccd1 _19825_/D
+ sky130_fd_sc_hd__o211a_1
X_14389_ _14472_/S vssd1 vssd1 vccd1 vccd1 _14402_/S sky130_fd_sc_hd__buf_2
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_152_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19721_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16128_ _13523_/X _19481_/Q _16128_/S vssd1 vssd1 vccd1 vccd1 _16129_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16059_ _16059_/A vssd1 vssd1 vccd1 vccd1 _19450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_167_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19938_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17453__A0 _17899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19818_ _19852_/CLK _19818_/D vssd1 vssd1 vccd1 vccd1 _19818_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10621__A _10621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19749_ _19756_/CLK _19749_/D vssd1 vssd1 vccd1 vccd1 _19749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09502_ _11428_/S vssd1 vssd1 vccd1 vccd1 _10560_/S sky130_fd_sc_hd__buf_2
XFILLER_53_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13490__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17756__A1 _11907_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09433_ _20050_/Q _20049_/Q vssd1 vssd1 vccd1 vccd1 _11723_/B sky130_fd_sc_hd__or2_1
XFILLER_25_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12548__A _17338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _20016_/Q _20015_/Q _20014_/Q _20013_/Q vssd1 vssd1 vccd1 vccd1 _09375_/A
+ sky130_fd_sc_hd__or4_4
Xclkbuf_leaf_105_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19288_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_123_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15859__A _15916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09997__B2 _19919_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09295_ _18313_/A _14148_/A _09290_/X _09292_/Y _09294_/Y vssd1 vssd1 vccd1 vccd1
+ _09295_/X sky130_fd_sc_hd__o2111a_1
XANTENNA__10068__A _10139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11005__B1 _11204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11100__S0 _10017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_108_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput160 _12495_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[26] sky130_fd_sc_hd__buf_2
XANTENNA__14702__S _14702_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__A1 _11482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput171 _11987_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[7] sky130_fd_sc_hd__buf_2
X_10070_ _11482_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10070_/X sky130_fd_sc_hd__and2_1
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09921__B2 _19917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14003__A _14059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12808__B2 _19820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15533__S _15539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13760_ _13760_/A vssd1 vssd1 vccd1 vccd1 _18541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10972_ _11032_/A _10967_/Y _10969_/Y _11221_/A vssd1 vssd1 vccd1 vccd1 _10972_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17747__A1 _17749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12711_ _12711_/A vssd1 vssd1 vccd1 vccd1 _12837_/A sky130_fd_sc_hd__clkbuf_4
X_13691_ _13691_/A vssd1 vssd1 vccd1 vccd1 _18525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15430_ _15430_/A vssd1 vssd1 vccd1 vccd1 _15439_/S sky130_fd_sc_hd__buf_4
X_12642_ _12651_/B vssd1 vssd1 vccd1 vccd1 _12649_/B sky130_fd_sc_hd__buf_8
XFILLER_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_6_0_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__13988__S _13994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15361_ _19188_/Q _15283_/X _15367_/S vssd1 vssd1 vccd1 vccd1 _15362_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12573_ _19987_/Q _11520_/A _12573_/S vssd1 vssd1 vccd1 vccd1 _12574_/A sky130_fd_sc_hd__mux2_4
XFILLER_8_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17100_ _19795_/Q _17097_/B _17099_/Y vssd1 vssd1 vccd1 vccd1 _19795_/D sky130_fd_sc_hd__o21a_1
XANTENNA__11795__A1 _11745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11524_ _18302_/A _17381_/A vssd1 vssd1 vccd1 vccd1 _11524_/Y sky130_fd_sc_hd__nor2_1
X_14312_ _14312_/A vssd1 vssd1 vccd1 vccd1 _18768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15292_ _15292_/A vssd1 vssd1 vccd1 vccd1 _15292_/X sky130_fd_sc_hd__clkbuf_1
X_18080_ _17791_/X _18076_/Y _18079_/Y vssd1 vssd1 vccd1 vccd1 _18080_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17031_ _19766_/Q _17033_/C _17030_/Y vssd1 vssd1 vccd1 vccd1 _19766_/D sky130_fd_sc_hd__o21a_1
XFILLER_7_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14243_ _14243_/A vssd1 vssd1 vccd1 vccd1 _18738_/D sky130_fd_sc_hd__clkbuf_1
X_11455_ _18792_/Q _19063_/Q _19287_/Q _19031_/Q _10053_/X _10054_/X vssd1 vssd1 vccd1
+ vccd1 _11455_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10406_ _18654_/Q _19245_/Q _19407_/Q _18622_/Q _10268_/S _10335_/A vssd1 vssd1 vccd1
+ vccd1 _10407_/B sky130_fd_sc_hd__mux4_1
X_14174_ _13780_/X _18708_/Q _14174_/S vssd1 vssd1 vccd1 vccd1 _14175_/A sky130_fd_sc_hd__mux2_1
X_11386_ _18808_/Q _19143_/Q _11386_/S vssd1 vssd1 vccd1 vccd1 _11387_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10755__C1 _10846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16486__A1 _19602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13125_ _13316_/A _15693_/B _15693_/C _13124_/X _13147_/S vssd1 vssd1 vccd1 vccd1
+ _13125_/X sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_84_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19431_/CLK sky130_fd_sc_hd__clkbuf_16
X_10337_ _10337_/A vssd1 vssd1 vccd1 vccd1 _10337_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18982_ _19464_/CLK _18982_/D vssd1 vssd1 vccd1 vccd1 _18982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13056_ _15206_/A vssd1 vssd1 vccd1 vccd1 _13056_/X sky130_fd_sc_hd__clkbuf_1
X_17933_ _17945_/A _17933_/B vssd1 vssd1 vccd1 vccd1 _17933_/Y sky130_fd_sc_hd__nand2_1
X_10268_ _18688_/Q _19183_/Q _10268_/S vssd1 vssd1 vccd1 vccd1 _10269_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17435__A0 _17610_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ _11870_/C _12153_/B _12006_/X _11977_/A vssd1 vssd1 vccd1 vccd1 _12007_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17864_ _17866_/A _17866_/B _18109_/S vssd1 vssd1 vccd1 vccd1 _17864_/X sky130_fd_sc_hd__mux2_1
X_10199_ _19120_/Q _18886_/Q _19568_/Q _19216_/Q _09812_/X _09822_/X vssd1 vssd1 vccd1
+ vccd1 _10199_/X sky130_fd_sc_hd__mux4_2
XFILLER_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_99_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19430_/CLK sky130_fd_sc_hd__clkbuf_16
X_19603_ _19987_/CLK _19603_/D vssd1 vssd1 vccd1 vccd1 _19603_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_120_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16815_ _19707_/Q _19706_/Q vssd1 vssd1 vccd1 vccd1 _16815_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__18965__D _18965_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17795_ _17785_/X _17790_/X _17793_/Y _17794_/X vssd1 vssd1 vccd1 vccd1 _17795_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15443__S _15443_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13752__A _13851_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19534_ _19988_/CLK _19534_/D vssd1 vssd1 vccd1 vccd1 _19534_/Q sky130_fd_sc_hd__dfxtp_1
X_16746_ _16747_/B _16747_/C _19686_/Q vssd1 vssd1 vccd1 vccd1 _16748_/B sky130_fd_sc_hd__a21oi_1
X_13958_ _13958_/A vssd1 vssd1 vccd1 vccd1 _18615_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19465_ _19497_/CLK _19465_/D vssd1 vssd1 vccd1 vccd1 _19465_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_22_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19919_/CLK sky130_fd_sc_hd__clkbuf_16
X_12909_ _12914_/A _16678_/A _12829_/X vssd1 vssd1 vccd1 vccd1 _12909_/X sky130_fd_sc_hd__o21a_1
X_16677_ _16680_/A _16680_/C _16676_/Y vssd1 vssd1 vccd1 vccd1 _19667_/D sky130_fd_sc_hd__o21a_1
X_13889_ _13796_/X _18585_/Q _13889_/S vssd1 vssd1 vccd1 vccd1 _13890_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10381__S1 _09520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18416_ _18336_/A _18413_/X _18414_/X _18415_/Y vssd1 vssd1 vccd1 vccd1 _18417_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15628_ _15628_/A vssd1 vssd1 vccd1 vccd1 _19306_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19396_ _19514_/CLK _19396_/D vssd1 vssd1 vccd1 vccd1 _19396_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13898__S _13900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18347_ _18347_/A _18349_/B vssd1 vssd1 vccd1 vccd1 _18347_/X sky130_fd_sc_hd__or2_1
X_15559_ _19276_/Q _15257_/X _15561_/S vssd1 vssd1 vccd1 vccd1 _15560_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_37_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19502_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12983__B1 _11520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__A _11141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18278_ _18335_/A vssd1 vssd1 vccd1 vccd1 _18311_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput40 io_ibus_inst[15] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
X_17229_ _17229_/A vssd1 vssd1 vccd1 vccd1 _17229_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput51 io_ibus_inst[25] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 io_ibus_inst[6] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15618__S _15622_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09982_ _11305_/S vssd1 vssd1 vccd1 vccd1 _09983_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__14522__S _14524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16303__A _16303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17134__A input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13463__B2 _19540_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14477__B _14477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10372__S1 _09520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _17247_/C vssd1 vssd1 vccd1 vccd1 _17346_/B sky130_fd_sc_hd__buf_4
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14412__A0 _18807_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09347_ _19890_/Q _13173_/B _19888_/Q vssd1 vssd1 vccd1 vccd1 _09347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10124__S1 _10014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11910__A _11910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09587__A _10519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09278_ _11624_/A _17336_/A _11624_/C _09278_/D vssd1 vssd1 vccd1 vccd1 _11809_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_21_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_3_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ _18574_/Q _18835_/Q _18734_/Q _19069_/Q _11129_/X _11115_/A vssd1 vssd1 vccd1
+ vccd1 _11241_/B sky130_fd_sc_hd__mux4_1
XFILLER_146_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11171_ _18765_/Q _19036_/Q _19260_/Q _19004_/Q _11147_/A _10007_/A vssd1 vssd1 vccd1
+ vccd1 _11171_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10122_ _10846_/A _10118_/X _10121_/X vssd1 vssd1 vccd1 vccd1 _10122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_103_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10053_ _10847_/S vssd1 vssd1 vccd1 vccd1 _10053_/X sky130_fd_sc_hd__buf_6
XFILLER_48_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14930_ _14987_/S vssd1 vssd1 vccd1 vccd1 _14939_/S sky130_fd_sc_hd__buf_2
XFILLER_76_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input26_A io_dbus_rdata[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14861_ _14596_/X _18976_/Q _14867_/S vssd1 vssd1 vccd1 vccd1 _14862_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16600_ _19640_/Q _16600_/B vssd1 vssd1 vccd1 vccd1 _16601_/B sky130_fd_sc_hd__and2_1
XFILLER_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13812_ _14637_/A vssd1 vssd1 vccd1 vccd1 _13812_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17580_ _17480_/X _17474_/X _17586_/S vssd1 vssd1 vccd1 vccd1 _17580_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14792_ _14792_/A vssd1 vssd1 vccd1 vccd1 _18949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16531_ _16550_/A _16538_/C vssd1 vssd1 vccd1 vccd1 _16531_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10955_ _10955_/A _10955_/B vssd1 vssd1 vccd1 vccd1 _10955_/X sky130_fd_sc_hd__or2_1
X_13743_ _14675_/A vssd1 vssd1 vccd1 vccd1 _13743_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19250_ _19412_/CLK _19250_/D vssd1 vssd1 vccd1 vccd1 _19250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16462_ _16462_/A vssd1 vssd1 vccd1 vccd1 _19586_/D sky130_fd_sc_hd__clkbuf_1
X_13674_ _13674_/A vssd1 vssd1 vccd1 vccd1 _18521_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17698__B _17702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10886_ _19364_/Q _18978_/Q _19428_/Q _18547_/Q _09983_/A _09513_/A vssd1 vssd1 vccd1
+ vccd1 _10887_/B sky130_fd_sc_hd__mux4_1
XFILLER_32_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18201_ _19957_/Q _19578_/Q _18209_/S vssd1 vssd1 vccd1 vccd1 _18202_/A sky130_fd_sc_hd__mux2_1
X_15413_ _14631_/X _19211_/Q _15417_/S vssd1 vssd1 vccd1 vccd1 _15414_/A sky130_fd_sc_hd__mux2_1
X_19181_ _19407_/CLK _19181_/D vssd1 vssd1 vccd1 vccd1 _19181_/Q sky130_fd_sc_hd__dfxtp_1
X_12625_ _12621_/X _12623_/Y _12624_/Y vssd1 vssd1 vccd1 vccd1 _12625_/Y sky130_fd_sc_hd__a21oi_1
X_16393_ _13195_/X _19555_/Q _16393_/S vssd1 vssd1 vccd1 vccd1 _16394_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18132_ _16206_/A _19959_/Q _18136_/S vssd1 vssd1 vccd1 vccd1 _18133_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09497__A _10937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12965__B1 _11562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15344_ _15344_/A vssd1 vssd1 vccd1 vccd1 _19180_/D sky130_fd_sc_hd__clkbuf_1
X_12556_ _12556_/A _18097_/B vssd1 vssd1 vccd1 vccd1 _12556_/Y sky130_fd_sc_hd__nor2_2
XFILLER_106_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ _19514_/Q _18926_/Q _18963_/Q _18537_/Q _11384_/S _10105_/A vssd1 vssd1 vccd1
+ vccd1 _11507_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13509__A2 _13353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18063_ _12463_/Y _18007_/X _18062_/X _18028_/X vssd1 vssd1 vccd1 vccd1 _18063_/X
+ sky130_fd_sc_hd__a211o_1
X_15275_ _15275_/A vssd1 vssd1 vccd1 vccd1 _19153_/D sky130_fd_sc_hd__clkbuf_1
X_12487_ _12487_/A _12511_/C vssd1 vssd1 vccd1 vccd1 _12487_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_156_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11031__S _11083_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17014_ _17046_/A _17014_/B _17014_/C vssd1 vssd1 vccd1 vccd1 _19761_/D sky130_fd_sc_hd__nor3_1
X_11438_ _11438_/A _11438_/B vssd1 vssd1 vccd1 vccd1 _11438_/X sky130_fd_sc_hd__or2_1
XFILLER_144_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14226_ _14294_/S vssd1 vssd1 vccd1 vccd1 _14235_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA_output94_A _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14157_ _13755_/X _18700_/Q _14163_/S vssd1 vssd1 vccd1 vccd1 _14158_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13747__A _14074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ _11362_/Y _11364_/Y _11366_/Y _11368_/Y _10834_/A vssd1 vssd1 vccd1 vccd1
+ _11369_/X sky130_fd_sc_hd__o221a_2
XANTENNA__12651__A _12651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ input28/X _12988_/X _13107_/X _13007_/X vssd1 vssd1 vccd1 vccd1 _15215_/A
+ sky130_fd_sc_hd__a22o_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18965_ _19666_/CLK _18965_/D vssd1 vssd1 vccd1 vccd1 _18965_/Q sky130_fd_sc_hd__dfxtp_2
X_14088_ _14088_/A vssd1 vssd1 vccd1 vccd1 _18671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13039_ _19708_/Q vssd1 vssd1 vccd1 vccd1 _16840_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17916_ _17725_/A _17917_/B _17915_/X _17722_/A vssd1 vssd1 vccd1 vccd1 _17919_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18896_ _19484_/CLK _18896_/D vssd1 vssd1 vccd1 vccd1 _18896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09992__S0 _10824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17847_ _17666_/S _17744_/Y _17846_/X vssd1 vssd1 vccd1 vccd1 _17847_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17778_ _18028_/A vssd1 vssd1 vccd1 vccd1 _17778_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13445__B2 _19539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19517_ _19831_/CLK _19517_/D vssd1 vssd1 vccd1 vccd1 _19517_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__11456__B1 _09706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16729_ _19681_/Q _19680_/Q _19679_/Q _16729_/D vssd1 vssd1 vccd1 vccd1 _16740_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_81_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16793__A _16818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15901__S _15901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19448_ _19510_/CLK _19448_/D vssd1 vssd1 vccd1 vccd1 _19448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09201_ _09201_/A vssd1 vssd1 vccd1 vccd1 _09215_/A sky130_fd_sc_hd__clkbuf_4
X_19379_ _19443_/CLK _19379_/D vssd1 vssd1 vccd1 vccd1 _19379_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18136__A1 _19961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10106__S1 _10718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11303__S0 _11004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12956__B1 _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13381__B1 _13054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11931__A1 _11352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09965_ _09952_/X _09962_/X _09963_/X _10840_/A _09964_/X vssd1 vssd1 vccd1 vccd1
+ _09978_/B sky130_fd_sc_hd__o221a_1
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10081__A _11483_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09896_ _09947_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _09896_/Y sky130_fd_sc_hd__nand2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10498__A1 _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10042__S0 _10700_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_10_0_clock_A clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10740_ _19367_/Q _18981_/Q _19431_/Q _18550_/Q _10608_/X _10682_/X vssd1 vssd1 vccd1
+ vccd1 _10741_/B sky130_fd_sc_hd__mux4_2
XFILLER_129_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10020__S _11384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11998__B2 _17412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10670__A1 _09748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ _10672_/A _12650_/A vssd1 vssd1 vccd1 vccd1 _10673_/A sky130_fd_sc_hd__and2_1
XFILLER_167_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12736__A _13578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ _12410_/A _18036_/B vssd1 vssd1 vccd1 vccd1 _12411_/B sky130_fd_sc_hd__and2_1
XFILLER_139_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ _13337_/X _13389_/X _13351_/X vssd1 vssd1 vccd1 vccd1 _13390_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_166_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12341_ _11818_/X _11819_/X _12340_/X _11977_/X vssd1 vssd1 vccd1 vccd1 _12341_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_166_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15060_ _15060_/A vssd1 vssd1 vccd1 vccd1 _19065_/D sky130_fd_sc_hd__clkbuf_1
X_12272_ _12196_/B _12272_/B _17964_/B _12272_/D vssd1 vssd1 vccd1 vccd1 _12300_/B
+ sky130_fd_sc_hd__and4b_1
X_14011_ _18638_/Q _13626_/X _14013_/S vssd1 vssd1 vccd1 vccd1 _14012_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13372__A0 _19913_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15258__S _15261_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _11223_/A vssd1 vssd1 vccd1 vccd1 _11223_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10186__B1 _09696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11922__A1 _11890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11154_ _18767_/Q _19038_/Q _19262_/Q _19006_/Q _11224_/S _11330_/A vssd1 vssd1 vccd1
+ vccd1 _11154_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_7_0_clock_A clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10105_ _10105_/A vssd1 vssd1 vccd1 vccd1 _10718_/A sky130_fd_sc_hd__buf_4
X_18750_ _19564_/CLK _18750_/D vssd1 vssd1 vccd1 vccd1 _18750_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15782__A _18458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15962_ _19407_/Q _15260_/X _15962_/S vssd1 vssd1 vccd1 vccd1 _15963_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11085_ _11085_/A _18672_/Q vssd1 vssd1 vccd1 vccd1 _11085_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17701_ _17698_/Y _17700_/X _17748_/S vssd1 vssd1 vccd1 vccd1 _17701_/X sky130_fd_sc_hd__mux2_1
X_10036_ _10041_/A vssd1 vssd1 vccd1 vccd1 _10037_/A sky130_fd_sc_hd__buf_2
X_14913_ _14672_/X _19000_/Q _14915_/S vssd1 vssd1 vccd1 vccd1 _14914_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09343__A2 _09342_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18681_ _19272_/CLK _18681_/D vssd1 vssd1 vccd1 vccd1 _18681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16089__S _16095_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15893_ _13376_/X _19376_/Q _15901_/S vssd1 vssd1 vccd1 vccd1 _15894_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output132_A _12669_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14398__A _14602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17632_ _17719_/A vssd1 vssd1 vccd1 vccd1 _17632_/X sky130_fd_sc_hd__clkbuf_2
X_14844_ _18299_/A _14917_/B _14844_/C _14844_/D vssd1 vssd1 vccd1 vccd1 _15990_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17563_ _17561_/X _17562_/X _17685_/S vssd1 vssd1 vccd1 vccd1 _17563_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11534__B _11534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14775_ _18942_/Q _14401_/X _14775_/S vssd1 vssd1 vccd1 vccd1 _14776_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11987_ _11987_/A vssd1 vssd1 vccd1 vccd1 _11987_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19302_ _19302_/CLK _19302_/D vssd1 vssd1 vccd1 vccd1 _19302_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11026__S _11026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16514_ _19611_/Q _16508_/C _16513_/Y vssd1 vssd1 vccd1 vccd1 _19611_/D sky130_fd_sc_hd__o21a_1
X_13726_ _15286_/A vssd1 vssd1 vccd1 vccd1 _14663_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17494_ _17675_/S vssd1 vssd1 vccd1 vccd1 _17799_/S sky130_fd_sc_hd__clkbuf_2
X_10938_ _11001_/A _10938_/B vssd1 vssd1 vccd1 vccd1 _10938_/X sky130_fd_sc_hd__and2_1
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19233_ _19395_/CLK _19233_/D vssd1 vssd1 vccd1 vccd1 _19233_/Q sky130_fd_sc_hd__dfxtp_1
X_16445_ _16445_/A vssd1 vssd1 vccd1 vccd1 _19578_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14337__S _14341_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13657_ _18517_/Q _13655_/X _13673_/S vssd1 vssd1 vccd1 vccd1 _13658_/A sky130_fd_sc_hd__mux2_1
X_10869_ _10869_/A _12644_/A vssd1 vssd1 vccd1 vccd1 _11578_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12646__A _12646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12938__B1 _11348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19164_ _19392_/CLK _19164_/D vssd1 vssd1 vccd1 vccd1 _19164_/Q sky130_fd_sc_hd__dfxtp_1
X_12608_ _18302_/A _12601_/A _12605_/X _12607_/X vssd1 vssd1 vccd1 vccd1 _12609_/D
+ sky130_fd_sc_hd__o31ai_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12402__A2 _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16376_ _13033_/X _19547_/Q _16382_/S vssd1 vssd1 vccd1 vccd1 _16377_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17326__C1 _12651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ _18439_/Q _13588_/B vssd1 vssd1 vccd1 vccd1 _13588_/X sky130_fd_sc_hd__or2_1
XFILLER_118_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18115_ _18054_/X _17606_/Y _18072_/X _18114_/X vssd1 vssd1 vccd1 vccd1 _18115_/X
+ sky130_fd_sc_hd__o211a_1
X_15327_ _15327_/A vssd1 vssd1 vccd1 vccd1 _19172_/D sky130_fd_sc_hd__clkbuf_1
X_19095_ _19575_/CLK _19095_/D vssd1 vssd1 vccd1 vccd1 _19095_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10166__A _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12539_ _19606_/Q _12540_/B vssd1 vssd1 vccd1 vccd1 _12539_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18333__A _18333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09377__D _12989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18046_ _18046_/A _18046_/B vssd1 vssd1 vccd1 vccd1 _18046_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09955__A _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15258_ _19148_/Q _15257_/X _15261_/S vssd1 vssd1 vccd1 vccd1 _15259_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14209_ _14209_/A vssd1 vssd1 vccd1 vccd1 _14218_/S sky130_fd_sc_hd__buf_4
XFILLER_99_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14072__S _14072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15189_ _19126_/Q vssd1 vssd1 vccd1 vccd1 _15190_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_99_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19997_ _19997_/CLK _19997_/D vssd1 vssd1 vccd1 vccd1 _19997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09750_ _09750_/A vssd1 vssd1 vccd1 vccd1 _09750_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__14800__S _14808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18948_ _19500_/CLK _18948_/D vssd1 vssd1 vccd1 vccd1 _18948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09681_ _11464_/A vssd1 vssd1 vccd1 vccd1 _10548_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18879_ _19305_/CLK _18879_/D vssd1 vssd1 vccd1 vccd1 _18879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10327__S1 _10326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15631__S _15633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17412__A _17412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16368__B1 _13604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11460__A _11460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10076__A _11014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10168__B1 _09580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11904__A1 _11082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10263__S0 _10216_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13106__A0 _19898_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ _09896_/Y _10145_/A _10143_/A vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__a21o_1
XFILLER_161_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09879_ _10229_/A _09875_/X _09878_/X vssd1 vssd1 vccd1 vccd1 _09879_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15107__A _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _11910_/A vssd1 vssd1 vccd1 vccd1 _12153_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_161_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _19729_/Q vssd1 vssd1 vccd1 vccd1 _16923_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _09407_/X _11950_/B _11840_/Y vssd1 vssd1 vccd1 vccd1 _11842_/B sky130_fd_sc_hd__a21oi_2
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18418__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16359__A0 _19543_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _13831_/X _18857_/Q _14568_/S vssd1 vssd1 vccd1 vccd1 _14561_/A sky130_fd_sc_hd__mux2_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _19814_/Q _19809_/Q vssd1 vssd1 vccd1 vccd1 _11772_/Y sky130_fd_sc_hd__nand2_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _10715_/Y _10717_/Y _10720_/Y _10722_/Y _09717_/A vssd1 vssd1 vccd1 vccd1
+ _10723_/X sky130_fd_sc_hd__o221a_2
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _16361_/A _13512_/B vssd1 vssd1 vccd1 vccd1 _13511_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17041__B _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14157__S _14163_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14491_ _17123_/A vssd1 vssd1 vccd1 vccd1 _14828_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16230_ _19519_/Q _16227_/X _16252_/S vssd1 vssd1 vccd1 vccd1 _16231_/A sky130_fd_sc_hd__mux2_1
X_10654_ _18777_/Q _19048_/Q _19272_/Q _19016_/Q _10653_/X _10645_/X vssd1 vssd1 vccd1
+ vccd1 _10654_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13442_ _19799_/Q vssd1 vssd1 vccd1 vccd1 _17112_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13996__S _13998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16161_ _19495_/Q _14612_/A _16167_/S vssd1 vssd1 vccd1 vccd1 _16162_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13373_ _13337_/X _13372_/X _13351_/X vssd1 vssd1 vccd1 vccd1 _13373_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__17859__B1 _17857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10585_ _10339_/A _10584_/X _10322_/A vssd1 vssd1 vccd1 vccd1 _10585_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14681__A _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15112_ _14647_/X _19088_/Q _15116_/S vssd1 vssd1 vccd1 vccd1 _15113_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15334__A1 _15244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12324_ _18001_/A _12324_/B vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__xor2_1
X_16092_ _16092_/A vssd1 vssd1 vccd1 vccd1 _19464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15043_ _15043_/A vssd1 vssd1 vccd1 vccd1 _19057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12255_ _19974_/Q _11562_/A _12303_/S vssd1 vssd1 vccd1 vccd1 _17445_/A sky130_fd_sc_hd__mux2_2
X_19920_ _19978_/CLK _19920_/D vssd1 vssd1 vccd1 vccd1 _19920_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_170_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_3_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ _18637_/Q _19228_/Q _19390_/Q _18605_/Q _11259_/S _10082_/A vssd1 vssd1 vccd1
+ vccd1 _11207_/B sky130_fd_sc_hd__mux4_1
X_19851_ _19852_/CLK _19851_/D vssd1 vssd1 vccd1 vccd1 _19851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_156_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12186_ _16226_/A _12184_/X _12185_/Y _11668_/X vssd1 vssd1 vccd1 vccd1 _12186_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11137_ _11153_/A _11137_/B vssd1 vssd1 vccd1 vccd1 _11137_/Y sky130_fd_sc_hd__nor2_1
X_18802_ _19042_/CLK _18802_/D vssd1 vssd1 vccd1 vccd1 _18802_/Q sky130_fd_sc_hd__dfxtp_1
X_19782_ _19782_/CLK _19782_/D vssd1 vssd1 vccd1 vccd1 _19782_/Q sky130_fd_sc_hd__dfxtp_1
X_16994_ _19756_/Q _19755_/Q _16994_/C _16994_/D vssd1 vssd1 vccd1 vccd1 _17005_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18733_ _19734_/CLK _18733_/D vssd1 vssd1 vccd1 vccd1 _18733_/Q sky130_fd_sc_hd__dfxtp_1
X_15945_ _19399_/Q _15235_/X _15951_/S vssd1 vssd1 vccd1 vccd1 _15946_/A sky130_fd_sc_hd__mux2_1
X_11068_ _11274_/A _11068_/B vssd1 vssd1 vccd1 vccd1 _11068_/X sky130_fd_sc_hd__or2_1
XFILLER_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13236__S _13299_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _10040_/A vssd1 vssd1 vccd1 vccd1 _11384_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_77_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18664_ _19063_/CLK _18664_/D vssd1 vssd1 vccd1 vccd1 _18664_/Q sky130_fd_sc_hd__dfxtp_1
X_15876_ _15876_/A vssd1 vssd1 vccd1 vccd1 _19368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17615_ _17791_/A vssd1 vssd1 vccd1 vccd1 _17616_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14827_ _18311_/A _14485_/X _14825_/X _14826_/Y vssd1 vssd1 vccd1 vccd1 _18402_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_18595_ _19476_/CLK _18595_/D vssd1 vssd1 vccd1 vccd1 _18595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18339__A1 _12475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18328__A _18328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17232__A _18289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17546_ _17721_/C _17614_/B vssd1 vssd1 vccd1 vccd1 _17917_/A sky130_fd_sc_hd__or2_1
X_14758_ _18934_/Q _14376_/X _14764_/S vssd1 vssd1 vccd1 vccd1 _14759_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10634__A1 _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13709_ _15273_/A vssd1 vssd1 vccd1 vccd1 _14650_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17477_ _17474_/X _17476_/X _17486_/S vssd1 vssd1 vccd1 vccd1 _17477_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12376__A _12376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14689_ _18899_/Q _14382_/X _14691_/S vssd1 vssd1 vccd1 vccd1 _14690_/A sky130_fd_sc_hd__mux2_1
X_19216_ _19313_/CLK _19216_/D vssd1 vssd1 vccd1 vccd1 _19216_/Q sky130_fd_sc_hd__dfxtp_1
X_16428_ _16428_/A vssd1 vssd1 vccd1 vccd1 _16437_/S sky130_fd_sc_hd__buf_4
XFILLER_20_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19147_ _19406_/CLK _19147_/D vssd1 vssd1 vccd1 vccd1 _19147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16359_ _19543_/Q _16358_/X _16365_/S vssd1 vssd1 vccd1 vccd1 _16360_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09685__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19078_ _19302_/CLK _19078_/D vssd1 vssd1 vccd1 vccd1 _19078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18029_ _12391_/Y _18007_/X _18027_/X _18028_/X vssd1 vssd1 vccd1 vccd1 _18029_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_133_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09802_ _09699_/A _09801_/X _09712_/X vssd1 vssd1 vccd1 vccd1 _09802_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09733_ _09722_/A _09729_/X _09732_/X vssd1 vssd1 vccd1 vccd1 _09733_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09664_ _10396_/A vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09595_ _09777_/A _09595_/B vssd1 vssd1 vccd1 vccd1 _09595_/X sky130_fd_sc_hd__or2_1
XANTENNA__14766__A _14823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15361__S _15367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16192__S _16200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14705__S _14713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ _09842_/A _10369_/X _10426_/A vssd1 vssd1 vccd1 vccd1 _10370_/X sky130_fd_sc_hd__a21o_1
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13327__A0 _19911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12040_ _12097_/A _12645_/B _12039_/X vssd1 vssd1 vccd1 vccd1 _17853_/A sky130_fd_sc_hd__a21o_1
XFILLER_85_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11353__A2 _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10561__B1 _10296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13991_ _13991_/A vssd1 vssd1 vccd1 vccd1 _18630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _19904_/Q _12854_/X _15757_/S vssd1 vssd1 vccd1 vccd1 _15730_/X sky130_fd_sc_hd__mux2_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _18321_/A _11135_/X _12942_/S vssd1 vssd1 vccd1 vccd1 _12942_/X sky130_fd_sc_hd__mux2_2
XFILLER_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17241__A1 _15839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10864__A1 _11383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15661_ _09341_/X _13572_/X _15719_/S vssd1 vssd1 vccd1 vccd1 _15661_/X sky130_fd_sc_hd__mux2_2
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _15680_/A _18449_/Q vssd1 vssd1 vccd1 vccd1 _12873_/Y sky130_fd_sc_hd__nand2_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _17419_/A vssd1 vssd1 vccd1 vccd1 _17465_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14612_ _14612_/A vssd1 vssd1 vccd1 vccd1 _14612_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17052__A _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _11824_/A _12207_/C vssd1 vssd1 vccd1 vccd1 _11825_/A sky130_fd_sc_hd__nor2_1
X_18380_ _18380_/A _18380_/B vssd1 vssd1 vccd1 vccd1 _20029_/D sky130_fd_sc_hd__nor2_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _14574_/X _19290_/Q _15600_/S vssd1 vssd1 vccd1 vccd1 _15593_/A sky130_fd_sc_hd__mux2_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17331_/A _17331_/B vssd1 vssd1 vccd1 vccd1 _17331_/X sky130_fd_sc_hd__or2_1
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14543_ _14543_/A vssd1 vssd1 vccd1 vccd1 _18849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11812__B _17431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11755_ _18316_/A _12937_/C _11754_/X _11704_/X vssd1 vssd1 vccd1 vccd1 _11755_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12196__A _12429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_82_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10706_ _11452_/A _10701_/Y _10703_/Y _11383_/A vssd1 vssd1 vccd1 vccd1 _10706_/X
+ sky130_fd_sc_hd__o211a_1
X_17262_ _17262_/A vssd1 vssd1 vccd1 vccd1 _19855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14474_ _16875_/A vssd1 vssd1 vccd1 vccd1 _18404_/A sky130_fd_sc_hd__clkbuf_4
X_11686_ _17381_/C _11686_/B vssd1 vssd1 vccd1 vccd1 _11901_/D sky130_fd_sc_hd__nand2_1
XFILLER_146_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19001_ _19576_/CLK _19001_/D vssd1 vssd1 vccd1 vccd1 _19001_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13566__A0 _11950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16213_ _16213_/A vssd1 vssd1 vccd1 vccd1 _16213_/X sky130_fd_sc_hd__clkbuf_2
X_13425_ _13425_/A vssd1 vssd1 vccd1 vccd1 _18492_/D sky130_fd_sc_hd__clkbuf_1
X_10637_ _10637_/A vssd1 vssd1 vccd1 vccd1 _11452_/A sky130_fd_sc_hd__clkbuf_2
X_17193_ _17191_/Y _17182_/X _17192_/X _17185_/X vssd1 vssd1 vccd1 vccd1 _19831_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10475__S0 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16144_ _16144_/A vssd1 vssd1 vccd1 vccd1 _19487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10568_ _19371_/Q _18985_/Q _19435_/Q _18554_/Q _10382_/A _09815_/A vssd1 vssd1 vccd1
+ vccd1 _10569_/B sky130_fd_sc_hd__mux4_1
X_13356_ _13336_/X _13352_/Y _13355_/Y vssd1 vssd1 vccd1 vccd1 _15260_/A sky130_fd_sc_hd__a21oi_4
XFILLER_115_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12643__B _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12307_ _12283_/A _12283_/B _12279_/A vssd1 vssd1 vccd1 vccd1 _12308_/B sky130_fd_sc_hd__a21bo_1
X_16075_ _16132_/S vssd1 vssd1 vccd1 vccd1 _16084_/S sky130_fd_sc_hd__buf_2
X_10499_ _19115_/Q _18881_/Q _19563_/Q _19211_/Q _10392_/S _10397_/X vssd1 vssd1 vccd1
+ vccd1 _10500_/B sky130_fd_sc_hd__mux4_1
X_13287_ _19625_/Q _12911_/X _13286_/X vssd1 vssd1 vccd1 vccd1 _13287_/X sky130_fd_sc_hd__o21a_1
XFILLER_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15026_ _15026_/A vssd1 vssd1 vccd1 vccd1 _19049_/D sky130_fd_sc_hd__clkbuf_1
X_19903_ _19952_/CLK _19903_/D vssd1 vssd1 vccd1 vccd1 _19903_/Q sky130_fd_sc_hd__dfxtp_4
X_12238_ _19594_/Q vssd1 vssd1 vccd1 vccd1 _16474_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18968__D _18968_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12541__A1 _11745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19834_ _19836_/CLK _19834_/D vssd1 vssd1 vccd1 vccd1 _19834_/Q sky130_fd_sc_hd__dfxtp_1
X_12169_ _12169_/A _17444_/A vssd1 vssd1 vccd1 vccd1 _12170_/B sky130_fd_sc_hd__or2_1
XFILLER_122_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17480__A1 _17853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19765_ _19768_/CLK _19765_/D vssd1 vssd1 vccd1 vccd1 _19765_/Q sky130_fd_sc_hd__dfxtp_1
X_16977_ _19750_/Q _16978_/C _16976_/Y vssd1 vssd1 vccd1 vccd1 _19750_/D sky130_fd_sc_hd__o21a_1
XFILLER_83_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput5 io_dbus_rdata[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
X_18716_ _19563_/CLK _18716_/D vssd1 vssd1 vccd1 vccd1 _18716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15928_ _15928_/A vssd1 vssd1 vccd1 vccd1 _19391_/D sky130_fd_sc_hd__clkbuf_1
X_19696_ _19726_/CLK _19696_/D vssd1 vssd1 vccd1 vccd1 _19696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12844__A2 _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18647_ _19464_/CLK _18647_/D vssd1 vssd1 vccd1 vccd1 _18647_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10855__A1 _10052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15859_ _15916_/S vssd1 vssd1 vccd1 vccd1 _15868_/S sky130_fd_sc_hd__buf_2
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09380_ _09398_/A vssd1 vssd1 vccd1 vccd1 _09394_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12057__B1 _12056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18578_ _19200_/CLK _18578_/D vssd1 vssd1 vccd1 vccd1 _18578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10607__A1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12818__B _12818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17529_ _17542_/A _11898_/X _17802_/C vssd1 vssd1 vccd1 vccd1 _17929_/A sky130_fd_sc_hd__o21ai_2
XFILLER_60_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11583__A2 _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10769__S1 _10037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14260__S _14268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09716_ _10063_/A vssd1 vssd1 vccd1 vccd1 _09717_/A sky130_fd_sc_hd__buf_2
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09647_ _09647_/A vssd1 vssd1 vccd1 vccd1 _10589_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__16187__S _16189_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15785__A1 _15784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09578_ _10307_/A vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_104_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ _11540_/A vssd1 vssd1 vccd1 vccd1 _11540_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11471_ _09807_/Y _11536_/A _11536_/B _11425_/Y _11470_/Y vssd1 vssd1 vccd1 vccd1
+ _11471_/X sky130_fd_sc_hd__a311o_1
XFILLER_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10422_ _10476_/A _10422_/B vssd1 vssd1 vccd1 vccd1 _10422_/X sky130_fd_sc_hd__or2_1
X_13210_ _16864_/A _13202_/X _13203_/X _19684_/Q _13209_/X vssd1 vssd1 vccd1 vccd1
+ _13210_/X sky130_fd_sc_hd__a221o_1
XFILLER_100_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11023__B2 _19899_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14190_ _13803_/X _18715_/Q _14196_/S vssd1 vssd1 vccd1 vccd1 _14191_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10353_ _10490_/A _10352_/X _09695_/A vssd1 vssd1 vccd1 vccd1 _10353_/Y sky130_fd_sc_hd__o21ai_1
X_13141_ _17146_/A _19824_/Q _17146_/B _13140_/X vssd1 vssd1 vccd1 vccd1 _13141_/X
+ sky130_fd_sc_hd__a31o_2
XANTENNA__12771__B2 _18454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13072_ _19929_/Q vssd1 vssd1 vccd1 vccd1 _16219_/B sky130_fd_sc_hd__buf_2
X_10284_ _19473_/Q _19311_/Q _18720_/Q _18490_/Q _09926_/S _09858_/A vssd1 vssd1 vccd1
+ vccd1 _10284_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input56_A io_ibus_inst[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15774__B _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16900_ _16924_/C _19730_/Q _19729_/Q _16900_/D vssd1 vssd1 vccd1 vccd1 _16909_/D
+ sky130_fd_sc_hd__and4_1
X_12023_ _12023_/A _12023_/B vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__xor2_2
XFILLER_151_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_opt_2_0_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_17880_ _17884_/A _17884_/B _18009_/A vssd1 vssd1 vccd1 vccd1 _17881_/B sky130_fd_sc_hd__mux2_1
XANTENNA__14170__S _14174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16831_ _19711_/Q _19710_/Q vssd1 vssd1 vccd1 vccd1 _16863_/D sky130_fd_sc_hd__and2_1
XFILLER_66_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19550_ _19794_/CLK _19550_/D vssd1 vssd1 vccd1 vccd1 _19550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16762_ _19691_/Q _16763_/C _19692_/Q vssd1 vssd1 vccd1 vccd1 _16764_/B sky130_fd_sc_hd__a21oi_1
XFILLER_47_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13974_ _13985_/A vssd1 vssd1 vccd1 vccd1 _13983_/S sky130_fd_sc_hd__buf_2
XFILLER_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18501_ _19745_/CLK _18501_/D vssd1 vssd1 vccd1 vccd1 _18501_/Q sky130_fd_sc_hd__dfxtp_1
X_15713_ _19901_/Q _15708_/X _15712_/Y vssd1 vssd1 vccd1 vccd1 _15713_/X sky130_fd_sc_hd__a21o_1
X_19481_ _19481_/CLK _19481_/D vssd1 vssd1 vccd1 vccd1 _19481_/Q sky130_fd_sc_hd__dfxtp_1
X_12925_ _12829_/X _15799_/A _12855_/B vssd1 vssd1 vccd1 vccd1 _12925_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16693_ _19672_/Q _16691_/B _16692_/Y vssd1 vssd1 vccd1 vccd1 _19672_/D sky130_fd_sc_hd__o21a_1
XFILLER_62_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18432_ _18435_/A _18432_/B vssd1 vssd1 vccd1 vccd1 _20051_/D sky130_fd_sc_hd__nor2_1
X_15644_ _14653_/X _19314_/Q _15644_/S vssd1 vssd1 vccd1 vccd1 _15645_/A sky130_fd_sc_hd__mux2_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _12856_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12856_/X sky130_fd_sc_hd__or2_1
XANTENNA__15776__A1 _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12638__B _12638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _18380_/A _18363_/B vssd1 vssd1 vccd1 vccd1 _20024_/D sky130_fd_sc_hd__nor2_1
X_11807_ _11807_/A _17662_/A vssd1 vssd1 vccd1 vccd1 _11812_/A sky130_fd_sc_hd__xor2_1
X_15575_ _19283_/Q _15279_/X _15583_/S vssd1 vssd1 vccd1 vccd1 _15576_/A sky130_fd_sc_hd__mux2_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _18455_/Q _12787_/B vssd1 vssd1 vccd1 vccd1 _12787_/X sky130_fd_sc_hd__or2_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17314_ _17314_/A vssd1 vssd1 vccd1 vccd1 _19879_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14572_/S vssd1 vssd1 vccd1 vccd1 _14535_/S sky130_fd_sc_hd__buf_4
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10696__S0 _10625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18294_ _20029_/Q _18291_/X _18293_/Y _18289_/X vssd1 vssd1 vccd1 vccd1 _19997_/D
+ sky130_fd_sc_hd__o211a_1
X_11738_ _17414_/A _12672_/A vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__nand2_2
XFILLER_147_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17245_ _19849_/Q _13595_/A _17245_/S vssd1 vssd1 vccd1 vccd1 _17246_/A sky130_fd_sc_hd__mux2_1
X_14457_ _18821_/Q _14456_/X _14466_/S vssd1 vssd1 vccd1 vccd1 _14458_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09947__B _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12654__A _12657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11669_ _12444_/A _11749_/B _12562_/S _11668_/X vssd1 vssd1 vccd1 vccd1 _16444_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12211__A0 _12204_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13408_ _19915_/Q _13407_/X _13483_/A vssd1 vssd1 vccd1 vccd1 _13408_/X sky130_fd_sc_hd__mux2_1
X_17176_ _17176_/A _17180_/B vssd1 vssd1 vccd1 vccd1 _17176_/X sky130_fd_sc_hd__or2_1
X_14388_ _14592_/A vssd1 vssd1 vccd1 vccd1 _14388_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16489__C1 _12908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16127_ _16127_/A vssd1 vssd1 vccd1 vccd1 _19480_/D sky130_fd_sc_hd__clkbuf_1
X_13339_ _19793_/Q vssd1 vssd1 vccd1 vccd1 _17095_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10773__B1 _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18341__A _18341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16058_ _13540_/X _19450_/Q _16060_/S vssd1 vssd1 vccd1 vccd1 _16059_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12514__A1 _19541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15009_ _19042_/Q _14398_/X _15011_/S vssd1 vssd1 vccd1 vccd1 _15010_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10902__A _11147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17453__A1 _17973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19817_ _19817_/CLK _19817_/D vssd1 vssd1 vccd1 vccd1 _19817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16796__A _16818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15904__S _15912_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10113__S _10751_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19748_ _19756_/CLK _19748_/D vssd1 vssd1 vccd1 vccd1 _19748_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12817__A2 _12814_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ _11429_/S vssd1 vssd1 vccd1 vccd1 _11428_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__09902__S _09902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19679_ _19682_/CLK _19679_/D vssd1 vssd1 vccd1 vccd1 _19679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09432_ _12320_/A vssd1 vssd1 vccd1 vccd1 _18324_/A sky130_fd_sc_hd__clkinv_2
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09363_ _09374_/A vssd1 vssd1 vccd1 vccd1 _12689_/B sky130_fd_sc_hd__buf_2
XFILLER_40_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09294_ _20039_/Q _14074_/B vssd1 vssd1 vccd1 vccd1 _09294_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__10068__B _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14255__S _14257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12564__A _19846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16036__A _16047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11005__A1 _10084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11100__S1 _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10084__A _10084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput150 _12269_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[17] sky130_fd_sc_hd__buf_2
Xoutput161 _12519_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[27] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_30_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15086__S _15094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 _16461_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[8] sky130_fd_sc_hd__buf_2
XFILLER_0_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10819__A1 _09475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10971_ _11342_/A vssd1 vssd1 vccd1 vccd1 _11221_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12710_ _19809_/Q _12684_/C _12696_/X _17199_/A _12709_/X vssd1 vssd1 vccd1 vccd1
+ _12710_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11492__A1 _09612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13690_ _18525_/Q _13689_/X _13694_/S vssd1 vssd1 vccd1 vccd1 _13691_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11492__B2 _19923_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _20044_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12641_ _12641_/A vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__buf_8
XFILLER_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11244__A1 _10875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15360_ _15360_/A vssd1 vssd1 vccd1 vccd1 _19187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12572_ _18111_/A _12572_/B vssd1 vssd1 vccd1 vccd1 _12576_/A sky130_fd_sc_hd__xor2_1
XANTENNA__15769__B _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14311_ _18768_/Q _13634_/X _14319_/S vssd1 vssd1 vccd1 vccd1 _14312_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11795__A2 _11767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11523_ _11523_/A vssd1 vssd1 vccd1 vccd1 _18302_/A sky130_fd_sc_hd__buf_2
XFILLER_168_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15291_ _15291_/A vssd1 vssd1 vccd1 vccd1 _19158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17030_ _19766_/Q _17033_/C _17021_/X vssd1 vssd1 vccd1 vccd1 _17030_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14242_ _13774_/X _18738_/Q _14246_/S vssd1 vssd1 vccd1 vccd1 _14243_/A sky130_fd_sc_hd__mux2_1
X_11454_ _18600_/Q _18861_/Q _18760_/Q _19095_/Q _10658_/X _10014_/X vssd1 vssd1 vccd1
+ vccd1 _11454_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17984__B _17985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _10407_/A _10404_/X _09696_/A vssd1 vssd1 vccd1 vccd1 _10405_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_137_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11385_ _11385_/A vssd1 vssd1 vccd1 vccd1 _11385_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16380__S _16382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14173_ _14173_/A vssd1 vssd1 vccd1 vccd1 _18707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16486__A2 _16449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13124_ _13371_/A _19899_/Q vssd1 vssd1 vccd1 vccd1 _13124_/X sky130_fd_sc_hd__or2_1
X_10336_ _10393_/A _10330_/Y _10335_/Y _10500_/A vssd1 vssd1 vccd1 vccd1 _10336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18981_ _19431_/CLK _18981_/D vssd1 vssd1 vccd1 vccd1 _18981_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output162_A _12547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _10439_/S vssd1 vssd1 vccd1 vccd1 _10268_/S sky130_fd_sc_hd__clkbuf_4
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _13036_/X _13051_/X _13054_/Y input23/X _12988_/X vssd1 vssd1 vccd1 vccd1
+ _15206_/A sky130_fd_sc_hd__a32o_4
X_17932_ _17627_/X _17513_/A _17632_/X vssd1 vssd1 vccd1 vccd1 _17932_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_140_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10507__B1 _09756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17435__A1 _12574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ _12027_/A _12027_/C vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__xor2_1
XANTENNA__11537__B _12667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17863_ _17866_/A _17866_/B vssd1 vssd1 vccd1 vccd1 _17863_/Y sky130_fd_sc_hd__nand2_1
X_10198_ _10161_/A _10197_/X _10256_/A vssd1 vssd1 vccd1 vccd1 _10198_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19602_ _19836_/CLK _19602_/D vssd1 vssd1 vccd1 vccd1 _19602_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16814_ _16814_/A _16814_/B vssd1 vssd1 vccd1 vccd1 _19706_/D sky130_fd_sc_hd__nor2_1
X_17794_ _17794_/A vssd1 vssd1 vccd1 vccd1 _17794_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16745_ _16747_/B _16747_/C _16744_/Y vssd1 vssd1 vccd1 vccd1 _19685_/D sky130_fd_sc_hd__o21a_1
XFILLER_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19533_ _19956_/CLK _19533_/D vssd1 vssd1 vccd1 vccd1 _19533_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13957_ _18615_/Q _13664_/X _13961_/S vssd1 vssd1 vccd1 vccd1 _13958_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12649__A _12649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19464_ _19464_/CLK _19464_/D vssd1 vssd1 vccd1 vccd1 _19464_/Q sky130_fd_sc_hd__dfxtp_1
X_12908_ _18281_/B vssd1 vssd1 vccd1 vccd1 _12908_/X sky130_fd_sc_hd__buf_6
X_16676_ _16680_/A _16680_/C _16667_/X vssd1 vssd1 vccd1 vccd1 _16676_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13888_ _13888_/A vssd1 vssd1 vccd1 vccd1 _18584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15627_ _14628_/X _19306_/Q _15633_/S vssd1 vssd1 vccd1 vccd1 _15628_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18415_ input51/X vssd1 vssd1 vccd1 vccd1 _18415_/Y sky130_fd_sc_hd__inv_2
X_12839_ _13204_/A vssd1 vssd1 vccd1 vccd1 _12839_/X sky130_fd_sc_hd__clkbuf_2
X_19395_ _19395_/CLK _19395_/D vssd1 vssd1 vccd1 vccd1 _19395_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18336__A _18336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18346_ _17338_/A _12883_/X _18345_/Y _18341_/X vssd1 vssd1 vccd1 vccd1 _20018_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17240__A _17240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15558_ _15558_/A vssd1 vssd1 vccd1 vccd1 _19275_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14509_ _13758_/X _18834_/Q _14513_/S vssd1 vssd1 vccd1 vccd1 _14510_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16174__A1 _14631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18277_ _19991_/Q _12825_/X _18276_/X _17243_/X vssd1 vssd1 vccd1 vccd1 _19991_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15489_ _19245_/Q _15260_/X _15489_/S vssd1 vssd1 vccd1 vccd1 _15490_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17228_ _17228_/A vssd1 vssd1 vccd1 vccd1 _17228_/Y sky130_fd_sc_hd__inv_2
Xinput30 io_dbus_rdata[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_6
XFILLER_174_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput41 io_ibus_inst[16] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
Xinput52 io_ibus_inst[26] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_8
XFILLER_128_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput63 io_ibus_inst[7] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17159_ _19820_/Q _17153_/X _17158_/X vssd1 vssd1 vccd1 vccd1 _19820_/D sky130_fd_sc_hd__a21o_1
XFILLER_155_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09693__A _09693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10841__S0 _11429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09981_ _09981_/A vssd1 vssd1 vccd1 vccd1 _11305_/S sky130_fd_sc_hd__buf_4
XFILLER_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14488__B2 _14487_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ _12857_/A _16208_/S vssd1 vssd1 vccd1 vccd1 _17247_/C sky130_fd_sc_hd__nand2_1
XFILLER_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10079__A _10606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11226__A1 _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ _19889_/Q vssd1 vssd1 vccd1 vccd1 _13173_/B sky130_fd_sc_hd__buf_4
XFILLER_21_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12974__A1 _18460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09277_ _09420_/A _11622_/A _09277_/C _09277_/D vssd1 vssd1 vccd1 vccd1 _09278_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14713__S _14713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11170_ _11170_/A vssd1 vssd1 vccd1 vccd1 _11183_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_7_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ _10790_/A _10120_/X _10043_/A vssd1 vssd1 vccd1 vccd1 _10121_/X sky130_fd_sc_hd__o21a_1
XFILLER_164_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10052_ _10790_/A vssd1 vssd1 vccd1 vccd1 _10052_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12765__D_N _12764_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13853__A _14148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14860_ _14860_/A vssd1 vssd1 vccd1 vccd1 _18975_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12683__A_N _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13811_ _13811_/A vssd1 vssd1 vccd1 vccd1 _18557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14791_ _18949_/Q _14424_/X _14797_/S vssd1 vssd1 vccd1 vccd1 _14792_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input19_A io_dbus_rdata[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16530_ _16540_/D vssd1 vssd1 vccd1 vccd1 _16538_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13742_ _15298_/A vssd1 vssd1 vccd1 vccd1 _14675_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_151_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19737_/CLK sky130_fd_sc_hd__clkbuf_16
X_10954_ _19491_/Q _18903_/Q _18940_/Q _18514_/Q _09530_/A _11236_/A vssd1 vssd1 vccd1
+ vccd1 _10955_/B sky130_fd_sc_hd__mux4_1
XFILLER_17_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16461_ _18404_/A _16461_/B vssd1 vssd1 vccd1 vccd1 _16462_/A sky130_fd_sc_hd__or2_1
X_13673_ _18521_/Q _13672_/X _13673_/S vssd1 vssd1 vccd1 vccd1 _13674_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10885_ _11491_/A _10885_/B _10885_/C vssd1 vssd1 vccd1 vccd1 _10885_/X sky130_fd_sc_hd__or3_2
X_18200_ _18268_/S vssd1 vssd1 vccd1 vccd1 _18209_/S sky130_fd_sc_hd__clkbuf_2
X_15412_ _15412_/A vssd1 vssd1 vccd1 vccd1 _19210_/D sky130_fd_sc_hd__clkbuf_1
X_19180_ _19407_/CLK _19180_/D vssd1 vssd1 vccd1 vccd1 _19180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12624_ _19545_/Q _12120_/X _16303_/A vssd1 vssd1 vccd1 vccd1 _12624_/Y sky130_fd_sc_hd__o21ai_1
X_16392_ _16392_/A vssd1 vssd1 vccd1 vccd1 _19554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18131_ _18131_/A vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_166_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19930_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12965__A1 _18454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15343_ _19180_/Q _15257_/X _15345_/S vssd1 vssd1 vccd1 vccd1 _15344_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12555_ _12555_/A vssd1 vssd1 vccd1 vccd1 _12555_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16156__A1 _14605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11506_ _11510_/A _11506_/B vssd1 vssd1 vccd1 vccd1 _11506_/Y sky130_fd_sc_hd__nor2_1
X_18062_ _18054_/X _17767_/Y _18061_/X _17953_/X vssd1 vssd1 vccd1 vccd1 _18062_/X
+ sky130_fd_sc_hd__o211a_1
X_15274_ _19153_/Q _15273_/X _15277_/S vssd1 vssd1 vccd1 vccd1 _15275_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ _19604_/Q vssd1 vssd1 vccd1 vccd1 _12487_/A sky130_fd_sc_hd__inv_2
XFILLER_144_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17013_ _19761_/Q _17016_/C _17013_/C vssd1 vssd1 vccd1 vccd1 _17014_/C sky130_fd_sc_hd__and3_1
X_14225_ _14281_/A vssd1 vssd1 vccd1 vccd1 _14294_/S sky130_fd_sc_hd__buf_4
X_11437_ _19385_/Q _18999_/Q _19449_/Q _18568_/Q _10625_/X _10691_/X vssd1 vssd1 vccd1
+ vccd1 _11438_/B sky130_fd_sc_hd__mux4_1
XANTENNA__11076__S0 _11000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output87_A _12436_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14156_ _14156_/A vssd1 vssd1 vccd1 vccd1 _18699_/D sky130_fd_sc_hd__clkbuf_1
X_11368_ _10732_/A _11367_/X _09976_/X vssd1 vssd1 vccd1 vccd1 _11368_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12651__B _12651_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13107_ _13095_/Y _13106_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10319_ _10378_/A _10318_/X _09826_/A vssd1 vssd1 vccd1 vccd1 _10319_/X sky130_fd_sc_hd__o21a_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ _19129_/CLK _18964_/D vssd1 vssd1 vccd1 vccd1 _18964_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _18671_/Q _13630_/X _14087_/S vssd1 vssd1 vccd1 vccd1 _14088_/A sky130_fd_sc_hd__mux2_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _19894_/Q vssd1 vssd1 vccd1 vccd1 _11299_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_104_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19418_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13038_/A vssd1 vssd1 vccd1 vccd1 _13299_/C sky130_fd_sc_hd__buf_2
X_17915_ _17985_/A _17918_/B _17539_/A _17914_/Y vssd1 vssd1 vccd1 vccd1 _17915_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18895_ _19285_/CLK _18895_/D vssd1 vssd1 vccd1 vccd1 _18895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15454__S _15456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18081__A1 _17543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17846_ _17702_/A _17655_/Y _17845_/Y _17931_/S vssd1 vssd1 vccd1 vccd1 _17846_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09992__S1 _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14989_ _15517_/B _15445_/B vssd1 vssd1 vccd1 vccd1 _15046_/A sky130_fd_sc_hd__nor2_4
XFILLER_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17777_ _17521_/X _17764_/X _17775_/X _17776_/X vssd1 vssd1 vccd1 vccd1 _17777_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_119_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19551_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11456__A1 _10052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19516_ _19831_/CLK _19516_/D vssd1 vssd1 vccd1 vccd1 _19516_/Q sky130_fd_sc_hd__dfxtp_1
X_16728_ _16728_/A _16728_/B _16728_/C vssd1 vssd1 vccd1 vccd1 _19680_/D sky130_fd_sc_hd__nor3_1
XFILLER_23_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19447_ _19511_/CLK _19447_/D vssd1 vssd1 vccd1 vccd1 _19447_/Q sky130_fd_sc_hd__dfxtp_1
X_16659_ _16661_/A _16661_/C _16624_/X vssd1 vssd1 vccd1 vccd1 _16659_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09200_ _09272_/C _09269_/B _09275_/D _11627_/C vssd1 vssd1 vccd1 vccd1 _09201_/A
+ sky130_fd_sc_hd__or4_1
XANTENNA__11208__A1 _11202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19378_ _19569_/CLK _19378_/D vssd1 vssd1 vccd1 vccd1 _19378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11303__S1 _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18329_ _18341_/A vssd1 vssd1 vccd1 vccd1 _18329_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12708__A1 _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15629__S _15633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11067__S0 _10999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14533__S _14535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09964_ _09979_/A vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09895_ _09750_/X _09880_/X _09893_/X _09757_/X _09894_/Y vssd1 vssd1 vccd1 vccd1
+ _12663_/B sky130_fd_sc_hd__o32a_4
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10042__S1 _11496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11695__A1 _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11905__B _17421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__A2 _11969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17583__A0 _17488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_83_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19464_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10670_ _09748_/A _10657_/X _10668_/X _09755_/A _10669_/Y vssd1 vssd1 vccd1 vccd1
+ _12650_/A sky130_fd_sc_hd__o32a_4
XFILLER_13_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09329_ _09329_/A _11789_/B vssd1 vssd1 vccd1 vccd1 _11690_/B sky130_fd_sc_hd__or2_1
XFILLER_139_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12340_ _12340_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _12340_/X sky130_fd_sc_hd__xor2_1
XANTENNA__17886__A1 _17533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_98_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19366_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_154_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15539__S _15539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12271_ _12188_/X _12655_/B _12270_/Y vssd1 vssd1 vccd1 vccd1 _17977_/B sky130_fd_sc_hd__a21o_2
X_14010_ _14010_/A vssd1 vssd1 vccd1 vccd1 _18637_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13372__A1 _13370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11222_ _18670_/Q _19165_/Q _11222_/S vssd1 vssd1 vccd1 vccd1 _11223_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19914_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10725__A3 _10723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11153_ _11153_/A _11153_/B vssd1 vssd1 vccd1 vccd1 _11153_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10104_ _10847_/S vssd1 vssd1 vccd1 vccd1 _11449_/S sky130_fd_sc_hd__buf_4
X_15961_ _15961_/A vssd1 vssd1 vccd1 vccd1 _19406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11084_ _19167_/Q vssd1 vssd1 vccd1 vccd1 _11084_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15782__B _15782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14679__A _18299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14912_ _14912_/A vssd1 vssd1 vccd1 vccd1 _18999_/D sky130_fd_sc_hd__clkbuf_1
X_10035_ _10751_/S vssd1 vssd1 vccd1 vccd1 _10640_/S sky130_fd_sc_hd__clkbuf_4
X_17700_ _17810_/S _17702_/B _18109_/S vssd1 vssd1 vccd1 vccd1 _17700_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18063__A1 _12463_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15892_ _15903_/A vssd1 vssd1 vccd1 vccd1 _15901_/S sky130_fd_sc_hd__buf_2
X_18680_ _19268_/CLK _18680_/D vssd1 vssd1 vccd1 vccd1 _18680_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_36_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19470_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14843_ _18359_/A _18407_/B vssd1 vssd1 vccd1 vccd1 _18969_/D sky130_fd_sc_hd__nor2_4
X_17631_ _17629_/X _17604_/B _17741_/S vssd1 vssd1 vccd1 vccd1 _17906_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output125_A _12662_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17562_ _17422_/X _17411_/X _17565_/S vssd1 vssd1 vccd1 vccd1 _17562_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14774_ _14774_/A vssd1 vssd1 vccd1 vccd1 _18941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11986_ _11986_/A _11986_/B vssd1 vssd1 vccd1 vccd1 _11987_/A sky130_fd_sc_hd__and2_4
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19301_ _19301_/CLK _19301_/D vssd1 vssd1 vccd1 vccd1 _19301_/Q sky130_fd_sc_hd__dfxtp_1
X_16513_ _16550_/A _16518_/C vssd1 vssd1 vccd1 vccd1 _16513_/Y sky130_fd_sc_hd__nor2_1
X_13725_ _13725_/A vssd1 vssd1 vccd1 vccd1 _18533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ _18674_/Q _19169_/Q _10937_/S vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__mux2_1
X_17493_ _17493_/A vssd1 vssd1 vccd1 vccd1 _17493_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_clkbuf_leaf_152_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11831__A _16268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15303__A _15371_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16444_ _18341_/A _19578_/Q _16444_/C vssd1 vssd1 vccd1 vccd1 _16445_/A sky130_fd_sc_hd__and3_1
X_19232_ _19490_/CLK _19232_/D vssd1 vssd1 vccd1 vccd1 _19232_/Q sky130_fd_sc_hd__dfxtp_1
X_13656_ _13744_/S vssd1 vssd1 vccd1 vccd1 _13673_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10868_ _10869_/A _12644_/A vssd1 vssd1 vccd1 vccd1 _11578_/A sky130_fd_sc_hd__or2_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19163_ _19258_/CLK _19163_/D vssd1 vssd1 vccd1 vccd1 _19163_/Q sky130_fd_sc_hd__dfxtp_1
X_12607_ _11601_/A _11730_/A _12610_/C _12601_/A vssd1 vssd1 vccd1 vccd1 _12607_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16375_ _16375_/A vssd1 vssd1 vccd1 vccd1 _19546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13587_ _13587_/A vssd1 vssd1 vccd1 vccd1 _13587_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _10775_/Y _10065_/X _09998_/X _10798_/X vssd1 vssd1 vccd1 vccd1 _12645_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18114_ _17626_/X _17595_/X _18113_/X _17619_/A vssd1 vssd1 vccd1 vccd1 _18114_/X
+ sky130_fd_sc_hd__a211o_1
X_15326_ _19172_/Q _15231_/X _15334_/S vssd1 vssd1 vccd1 vccd1 _15327_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11071__C1 _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19094_ _19574_/CLK _19094_/D vssd1 vssd1 vccd1 vccd1 _19094_/Q sky130_fd_sc_hd__dfxtp_1
X_12538_ _12538_/A _12538_/B vssd1 vssd1 vccd1 vccd1 _12538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18045_ _18043_/Y _18044_/X _18078_/S vssd1 vssd1 vccd1 vccd1 _18045_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15257_ _15257_/A vssd1 vssd1 vccd1 vccd1 _15257_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12662__A _12663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12469_ _17223_/A _12470_/C _19842_/Q vssd1 vssd1 vccd1 vccd1 _12469_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_172_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14208_ _14208_/A vssd1 vssd1 vccd1 vccd1 _18723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15188_ _15188_/A vssd1 vssd1 vccd1 vccd1 _19125_/D sky130_fd_sc_hd__clkbuf_1
X_14139_ _14139_/A vssd1 vssd1 vccd1 vccd1 _18694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19996_ _20052_/CLK _19996_/D vssd1 vssd1 vccd1 vccd1 _19996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18947_ _19498_/CLK _18947_/D vssd1 vssd1 vccd1 vccd1 _18947_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_77_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14589__A _14589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09680_ _09680_/A vssd1 vssd1 vccd1 vccd1 _11464_/A sky130_fd_sc_hd__buf_4
X_18878_ _19302_/CLK _18878_/D vssd1 vssd1 vccd1 vccd1 _18878_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10910__A _10910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17829_ _17832_/A _17832_/B vssd1 vssd1 vccd1 vccd1 _17829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15912__S _15912_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12626__B1 _19848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12837__A _12837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17317__A0 _13603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15359__S _15367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09881__A _10216_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09947_ _09947_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _10143_/A sky130_fd_sc_hd__nor2_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15094__S _15094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11916__A _19519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09878_ _10283_/A _09877_/X _09711_/A vssd1 vssd1 vccd1 vccd1 _09878_/X sky130_fd_sc_hd__o21a_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10876__C1 _10875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _09354_/B _11839_/X _13604_/A vssd1 vssd1 vccd1 vccd1 _11840_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13290__A0 _19908_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11771_ _12628_/A vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__buf_4
XANTENNA__10966__S _11026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17556__B1 _09341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16219__A _16219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _19954_/Q vssd1 vssd1 vccd1 vccd1 _16361_/A sky130_fd_sc_hd__clkbuf_4
X_10722_ _10764_/A _10721_/X _10655_/X vssd1 vssd1 vccd1 vccd1 _10722_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _16678_/A vssd1 vssd1 vccd1 vccd1 _17123_/A sky130_fd_sc_hd__buf_4
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13441_ _19667_/Q vssd1 vssd1 vccd1 vccd1 _16680_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10653_ _10700_/S vssd1 vssd1 vccd1 vccd1 _10653_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10267__A _10439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16160_ _16160_/A vssd1 vssd1 vccd1 vccd1 _19494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17859__A1 _12056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13372_ _19913_/Q _13370_/X _13483_/A vssd1 vssd1 vccd1 vccd1 _13372_/X sky130_fd_sc_hd__mux2_1
X_10584_ _19467_/Q _19305_/Q _18714_/Q _18484_/Q _10533_/S _09665_/A vssd1 vssd1 vccd1
+ vccd1 _10584_/X sky130_fd_sc_hd__mux4_1
X_15111_ _15111_/A vssd1 vssd1 vccd1 vccd1 _19087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12323_ _17989_/B _12301_/B _12252_/A vssd1 vssd1 vccd1 vccd1 _12324_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__13578__A _13578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16091_ _13239_/X _19464_/Q _16095_/S vssd1 vssd1 vccd1 vccd1 _16092_/A sky130_fd_sc_hd__mux2_1
X_15042_ _19057_/Q _14446_/X _15044_/S vssd1 vssd1 vccd1 vccd1 _15043_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13345__B2 _19533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ _17964_/B _12254_/B vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__xnor2_4
XFILLER_135_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17484__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ _19454_/Q _19292_/Q _18701_/Q _18471_/Q _10937_/S _09954_/A vssd1 vssd1 vccd1
+ vccd1 _11205_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19850_ _19881_/CLK _19850_/D vssd1 vssd1 vccd1 vccd1 _19850_/Q sky130_fd_sc_hd__dfxtp_1
X_12185_ _17192_/A _12217_/C vssd1 vssd1 vccd1 vccd1 _12185_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18801_ _19042_/CLK _18801_/D vssd1 vssd1 vccd1 vccd1 _18801_/Q sky130_fd_sc_hd__dfxtp_1
X_11136_ _19360_/Q _18974_/Q _19424_/Q _18543_/Q _11035_/X _11168_/A vssd1 vssd1 vccd1
+ vccd1 _11137_/B sky130_fd_sc_hd__mux4_1
XFILLER_110_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19781_ _19783_/CLK _19781_/D vssd1 vssd1 vccd1 vccd1 _19781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16993_ _16993_/A _16993_/B _16993_/C vssd1 vssd1 vccd1 vccd1 _19755_/D sky130_fd_sc_hd__nor3_1
XANTENNA__11108__B1 _09752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18732_ _19734_/CLK _18732_/D vssd1 vssd1 vccd1 vccd1 _18732_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11203__S0 _11306_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10730__A _10730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15944_ _15944_/A vssd1 vssd1 vccd1 vccd1 _19398_/D sky130_fd_sc_hd__clkbuf_1
X_11067_ _18576_/Q _18837_/Q _18736_/Q _19071_/Q _10999_/A _10082_/A vssd1 vssd1 vccd1
+ vccd1 _11068_/B sky130_fd_sc_hd__mux4_1
XFILLER_23_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17244__C1 _17243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10018_ _10018_/A vssd1 vssd1 vccd1 vccd1 _10040_/A sky130_fd_sc_hd__clkbuf_4
X_15875_ _13239_/X _19368_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15876_/A sky130_fd_sc_hd__mux2_1
X_18663_ _19512_/CLK _18663_/D vssd1 vssd1 vccd1 vccd1 _18663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14826_ input40/X vssd1 vssd1 vccd1 vccd1 _14826_/Y sky130_fd_sc_hd__clkinv_4
X_17614_ _17721_/C _17614_/B vssd1 vssd1 vccd1 vccd1 _17791_/A sky130_fd_sc_hd__nor2_2
XFILLER_92_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18594_ _19313_/CLK _18594_/D vssd1 vssd1 vccd1 vccd1 _18594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17545_ _17721_/A _17545_/B vssd1 vssd1 vccd1 vccd1 _17614_/B sky130_fd_sc_hd__nand2_1
X_14757_ _14757_/A vssd1 vssd1 vccd1 vccd1 _18933_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12657__A _12657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11969_ _11969_/A vssd1 vssd1 vccd1 vccd1 _17772_/B sky130_fd_sc_hd__buf_2
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13708_ _13708_/A vssd1 vssd1 vccd1 vccd1 _18529_/D sky130_fd_sc_hd__clkbuf_1
X_17476_ _12407_/A _17820_/B _17506_/S vssd1 vssd1 vccd1 vccd1 _17476_/X sky130_fd_sc_hd__mux2_1
X_14688_ _14688_/A vssd1 vssd1 vccd1 vccd1 _18898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19215_ _19570_/CLK _19215_/D vssd1 vssd1 vccd1 vccd1 _19215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16427_ _16427_/A vssd1 vssd1 vccd1 vccd1 _19570_/D sky130_fd_sc_hd__clkbuf_1
X_13639_ _14596_/A vssd1 vssd1 vccd1 vccd1 _13639_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13584__A1 _12421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19146_ _19405_/CLK _19146_/D vssd1 vssd1 vccd1 vccd1 _19146_/Q sky130_fd_sc_hd__dfxtp_1
X_16358_ _15833_/X _16357_/Y _16364_/S vssd1 vssd1 vccd1 vccd1 _16358_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15309_ _15309_/A vssd1 vssd1 vccd1 vccd1 _19164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19077_ _19431_/CLK _19077_/D vssd1 vssd1 vccd1 vccd1 _19077_/Q sky130_fd_sc_hd__dfxtp_1
X_16289_ _19941_/Q _16290_/B vssd1 vssd1 vccd1 vccd1 _16301_/C sky130_fd_sc_hd__or2_1
XFILLER_145_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18028_ _18028_/A vssd1 vssd1 vccd1 vccd1 _18028_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11347__B1 _11324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16799__A _16818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11442__S0 _11372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14811__S _14819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09801_ _18663_/Q _19254_/Q _19416_/Q _18631_/Q _09724_/S _09730_/X vssd1 vssd1 vccd1
+ vccd1 _09801_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19979_ _19986_/CLK _19979_/D vssd1 vssd1 vccd1 vccd1 _19979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14836__B2 _14835_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ _09699_/A _09731_/X _09712_/X vssd1 vssd1 vccd1 vccd1 _09732_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09663_ _10703_/A vssd1 vssd1 vccd1 vccd1 _10396_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09594_ _18666_/Q _19257_/Q _19419_/Q _18634_/Q _09568_/X _09762_/A vssd1 vssd1 vccd1
+ vccd1 _09595_/B sky130_fd_sc_hd__mux4_1
XFILLER_83_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13024__B1 _13343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09779__B1 _09580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13398__A _13418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13327__A1 _12787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_100_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11433__S0 _10081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10561__A1 _10294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14827__B2 _14826_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18018__A1 _19914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15118__A _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13990_ _18630_/Q _13727_/X _13994_/S vssd1 vssd1 vccd1 vccd1 _13991_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12941_ _12941_/A vssd1 vssd1 vccd1 vccd1 _18440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _15660_/A vssd1 vssd1 vccd1 vccd1 _19321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _18449_/Q _12872_/B vssd1 vssd1 vccd1 vccd1 _12872_/X sky130_fd_sc_hd__or2_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14611_/A vssd1 vssd1 vccd1 vccd1 _18874_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _19581_/Q _11868_/C vssd1 vssd1 vccd1 vccd1 _11823_/X sky130_fd_sc_hd__xor2_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15591_ _15659_/S vssd1 vssd1 vccd1 vccd1 _15600_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14168__S _14174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17392_/A vssd1 vssd1 vccd1 vccd1 _18118_/A sky130_fd_sc_hd__buf_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14542_ _13806_/X _18849_/Q _14546_/S vssd1 vssd1 vccd1 vccd1 _14543_/A sky130_fd_sc_hd__mux2_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11754_ _12378_/A _17327_/B _11895_/C vssd1 vssd1 vccd1 vccd1 _11754_/X sky130_fd_sc_hd__and3_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_25_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _11510_/A vssd1 vssd1 vccd1 vccd1 _11383_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__17479__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17261_ _15688_/X _19855_/Q _17269_/S vssd1 vssd1 vccd1 vccd1 _17262_/A sky130_fd_sc_hd__mux2_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14473_/A vssd1 vssd1 vccd1 vccd1 _18826_/D sky130_fd_sc_hd__clkbuf_1
X_11685_ _12602_/A _12600_/A _12595_/C _17325_/B vssd1 vssd1 vccd1 vccd1 _11686_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_41_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19000_ _19482_/CLK _19000_/D vssd1 vssd1 vccd1 vccd1 _19000_/Q sky130_fd_sc_hd__dfxtp_1
X_16212_ _16212_/A vssd1 vssd1 vccd1 vccd1 _19516_/D sky130_fd_sc_hd__clkbuf_1
X_13424_ _18492_/Q _13423_/X _13434_/S vssd1 vssd1 vccd1 vccd1 _13425_/A sky130_fd_sc_hd__mux2_1
X_10636_ _09614_/A _10623_/X _10635_/X _09621_/A _19907_/Q vssd1 vssd1 vccd1 vccd1
+ _10672_/A sky130_fd_sc_hd__a32o_4
XFILLER_139_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17192_ _17192_/A _17195_/B vssd1 vssd1 vccd1 vccd1 _17192_/X sky130_fd_sc_hd__or2_1
XFILLER_128_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16143_ _19487_/Q _14586_/A _16145_/S vssd1 vssd1 vccd1 vccd1 _16144_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13355_ input11/X _13353_/X _13354_/X vssd1 vssd1 vccd1 vccd1 _13355_/Y sky130_fd_sc_hd__a21oi_2
X_10567_ _10314_/A _10558_/X _10562_/X _10566_/X _10519_/A vssd1 vssd1 vccd1 vccd1
+ _10567_/X sky130_fd_sc_hd__a311o_2
XFILLER_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12306_ _12306_/A _12306_/B vssd1 vssd1 vccd1 vccd1 _12308_/A sky130_fd_sc_hd__and2_1
XFILLER_154_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16074_ _16074_/A vssd1 vssd1 vccd1 vccd1 _19456_/D sky130_fd_sc_hd__clkbuf_1
X_13286_ _19753_/Q _12912_/X _13285_/X _12917_/X vssd1 vssd1 vccd1 vccd1 _13286_/X
+ sky130_fd_sc_hd__a211o_1
X_10498_ _09667_/A _10495_/Y _10497_/Y _10486_/A vssd1 vssd1 vccd1 vccd1 _10498_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15025_ _19049_/Q _14420_/X _15033_/S vssd1 vssd1 vccd1 vccd1 _15026_/A sky130_fd_sc_hd__mux2_1
X_19902_ _19986_/CLK _19902_/D vssd1 vssd1 vccd1 vccd1 _19902_/Q sky130_fd_sc_hd__dfxtp_4
X_12237_ _19591_/Q hold18/A _12237_/C _12237_/D vssd1 vssd1 vccd1 vccd1 _12240_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_151_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19833_ _19836_/CLK _19833_/D vssd1 vssd1 vccd1 vccd1 _19833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12168_ _12169_/A _17444_/A vssd1 vssd1 vccd1 vccd1 _12170_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11119_ _18767_/Q _19038_/Q _19262_/Q _19006_/Q _11004_/S _11061_/A vssd1 vssd1 vccd1
+ vccd1 _11119_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19764_ _19768_/CLK _19764_/D vssd1 vssd1 vccd1 vccd1 _19764_/Q sky130_fd_sc_hd__dfxtp_1
X_16976_ _17007_/A _16984_/D vssd1 vssd1 vccd1 vccd1 _16976_/Y sky130_fd_sc_hd__nor2_1
X_12099_ _18349_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12319_/B sky130_fd_sc_hd__nand2_2
XFILLER_77_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18715_ _19561_/CLK _18715_/D vssd1 vssd1 vccd1 vccd1 _18715_/Q sky130_fd_sc_hd__dfxtp_1
Xinput6 io_dbus_rdata[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15927_ _19391_/Q _15209_/X _15929_/S vssd1 vssd1 vccd1 vccd1 _15928_/A sky130_fd_sc_hd__mux2_1
X_19695_ _19726_/CLK _19695_/D vssd1 vssd1 vccd1 vccd1 _19695_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17243__A _18289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13771__A _14596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18646_ _18777_/CLK _18646_/D vssd1 vssd1 vccd1 vccd1 _18646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15858_ _15858_/A vssd1 vssd1 vccd1 vccd1 _19360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14809_ _14809_/A vssd1 vssd1 vccd1 vccd1 _18957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18577_ _19200_/CLK _18577_/D vssd1 vssd1 vccd1 vccd1 _18577_/Q sky130_fd_sc_hd__dfxtp_1
X_15789_ _18459_/Q _13407_/X _15788_/Y _15700_/X vssd1 vssd1 vccd1 vccd1 _15789_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17528_ _17719_/A vssd1 vssd1 vccd1 vccd1 _17530_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17459_ _17459_/A vssd1 vssd1 vccd1 vccd1 _17832_/B sky130_fd_sc_hd__buf_2
XANTENNA__14806__S _14808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09696__A _09696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19129_ _19129_/CLK _19129_/D vssd1 vssd1 vccd1 vccd1 _19129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13011__A _14074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17418__A _17418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16259__A0 _19524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09715_ _10994_/A vssd1 vssd1 vccd1 vccd1 _10063_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12296__A1 _12127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14777__A _14823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13681__A _14628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17153__A _17229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09646_ _10849_/S vssd1 vssd1 vccd1 vccd1 _09647_/A sky130_fd_sc_hd__buf_8
XFILLER_56_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09577_ _09577_/A vssd1 vssd1 vccd1 vccd1 _10307_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18184__A0 _19950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10154__S0 _09508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14716__S _14724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13548__B2 _19848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11470_ _11470_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _11470_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10421_ _18589_/Q _18850_/Q _18749_/Q _19084_/Q _10466_/S _10312_/A vssd1 vssd1 vccd1
+ vccd1 _10422_/B sky130_fd_sc_hd__mux4_1
XFILLER_137_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10231__B1 _09696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13140_ _19811_/Q _12798_/Y _13138_/X _13139_/X vssd1 vssd1 vccd1 vccd1 _13140_/X
+ sky130_fd_sc_hd__a211o_1
X_10352_ _19504_/Q _18916_/Q _18953_/Q _18527_/Q _10325_/X _10326_/X vssd1 vssd1 vccd1
+ vccd1 _10352_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _13071_/A vssd1 vssd1 vccd1 vccd1 _18472_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17964__A_N _17960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ _10283_/A _10283_/B vssd1 vssd1 vccd1 vccd1 _10283_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12022_ _12002_/A _12002_/B _12052_/A vssd1 vssd1 vccd1 vccd1 _12023_/B sky130_fd_sc_hd__a21o_1
XFILLER_2_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input49_A io_ibus_inst[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16830_ _19710_/Q _16863_/C _16829_/Y vssd1 vssd1 vccd1 vccd1 _19710_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13973_ _13973_/A vssd1 vssd1 vccd1 vccd1 _18622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16761_ _19691_/Q _16763_/C _16760_/Y vssd1 vssd1 vccd1 vccd1 _19691_/D sky130_fd_sc_hd__o21a_1
XANTENNA__16378__S _16382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13591__A _13591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18500_ _19577_/CLK _18500_/D vssd1 vssd1 vccd1 vccd1 _18500_/Q sky130_fd_sc_hd__dfxtp_1
X_15712_ _16364_/S _17175_/A vssd1 vssd1 vccd1 vccd1 _15712_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12924_ _18461_/Q _12903_/A _12923_/X vssd1 vssd1 vccd1 vccd1 _15799_/A sky130_fd_sc_hd__a21oi_4
X_19480_ _19480_/CLK _19480_/D vssd1 vssd1 vccd1 vccd1 _19480_/Q sky130_fd_sc_hd__dfxtp_1
X_16692_ _16731_/A _16692_/B vssd1 vssd1 vccd1 vccd1 _16692_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18431_ _18347_/A _17138_/B _14486_/X _18430_/Y vssd1 vssd1 vccd1 vccd1 _18432_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_46_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15643_ _15643_/A vssd1 vssd1 vccd1 vccd1 _19313_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12855_ _12855_/A _12855_/B vssd1 vssd1 vccd1 vccd1 _12856_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11806_ _11849_/D vssd1 vssd1 vccd1 vccd1 _17662_/A sky130_fd_sc_hd__clkbuf_2
X_15574_ _15574_/A vssd1 vssd1 vccd1 vccd1 _15583_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18362_ _18279_/A _12795_/X _14831_/X _18361_/Y vssd1 vssd1 vccd1 vccd1 _18363_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_109_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12786_/A _12786_/B _12785_/Y vssd1 vssd1 vccd1 vccd1 _12787_/B sky130_fd_sc_hd__or3b_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _15833_/X _19879_/Q _17313_/S vssd1 vssd1 vccd1 vccd1 _17314_/A sky130_fd_sc_hd__mux2_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14525_/A vssd1 vssd1 vccd1 vccd1 _18841_/D sky130_fd_sc_hd__clkbuf_1
X_11737_ _19957_/Q _11324_/X _11809_/A vssd1 vssd1 vccd1 vccd1 _12672_/A sky130_fd_sc_hd__mux2_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14626__S _14638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10696__S1 _10691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18293_ _18293_/A _18326_/B vssd1 vssd1 vccd1 vccd1 _18293_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12935__A _12935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14456_ _14660_/A vssd1 vssd1 vccd1 vccd1 _14456_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17244_ _13603_/B _17197_/A _17242_/X _17243_/X vssd1 vssd1 vccd1 vccd1 _19848_/D
+ sky130_fd_sc_hd__o211a_1
X_11668_ _11797_/A vssd1 vssd1 vccd1 vccd1 _11668_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12654__B _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13407_ _16670_/B _13116_/X _13117_/X _17104_/B _13406_/X vssd1 vssd1 vccd1 vccd1
+ _13407_/X sky130_fd_sc_hd__a221o_4
X_10619_ _18585_/Q _18846_/Q _18745_/Q _19080_/Q _10617_/X _10682_/A vssd1 vssd1 vccd1
+ vccd1 _10620_/B sky130_fd_sc_hd__mux4_1
X_17175_ _17175_/A vssd1 vssd1 vccd1 vccd1 _17175_/Y sky130_fd_sc_hd__inv_2
X_14387_ _14387_/A vssd1 vssd1 vccd1 vccd1 _18799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11599_ _11603_/A _17331_/B vssd1 vssd1 vccd1 vccd1 _11599_/X sky130_fd_sc_hd__or2_1
XFILLER_143_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10222__B1 _09696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16126_ _13506_/X _19480_/Q _16128_/S vssd1 vssd1 vccd1 vccd1 _16127_/A sky130_fd_sc_hd__mux2_1
X_13338_ _19661_/Q vssd1 vssd1 vccd1 vccd1 _16661_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10773__A1 _09748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10773__B2 _10772_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16057_ _16057_/A vssd1 vssd1 vccd1 vccd1 _19449_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17238__A _19846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14361__S _14363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ _19656_/Q _12727_/X _12729_/X _19788_/Q _13268_/X vssd1 vssd1 vccd1 vccd1
+ _13269_/X sky130_fd_sc_hd__a221o_1
XANTENNA__12670__A _12670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ _15008_/A vssd1 vssd1 vccd1 vccd1 _19041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19816_ _19857_/CLK _19816_/D vssd1 vssd1 vccd1 vccd1 _19816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19747_ _19756_/CLK _19747_/D vssd1 vssd1 vccd1 vccd1 _19747_/Q sky130_fd_sc_hd__dfxtp_1
X_16959_ _19746_/Q _16959_/B _16959_/C vssd1 vssd1 vccd1 vccd1 _16967_/C sky130_fd_sc_hd__and3_1
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09500_ _10824_/S vssd1 vssd1 vccd1 vccd1 _11429_/S sky130_fd_sc_hd__buf_4
XANTENNA__10828__A2 _19555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19678_ _19682_/CLK _19678_/D vssd1 vssd1 vccd1 vccd1 _19678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09431_ _20041_/Q vssd1 vssd1 vccd1 vccd1 _12320_/A sky130_fd_sc_hd__clkbuf_2
X_18629_ _19510_/CLK _18629_/D vssd1 vssd1 vccd1 vccd1 _18629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09362_ _20018_/Q _20017_/Q _20020_/Q _20019_/Q vssd1 vssd1 vccd1 vccd1 _09374_/A
+ sky130_fd_sc_hd__or4bb_2
XFILLER_80_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09293_ _19999_/Q vssd1 vssd1 vccd1 vccd1 _14074_/B sky130_fd_sc_hd__buf_4
XFILLER_166_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12450__B2 _12449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15367__S _15367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13676__A _14624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14271__S _14279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17148__A _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 _12644_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[9] sky130_fd_sc_hd__buf_2
Xoutput151 _12297_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[18] sky130_fd_sc_hd__buf_2
XFILLER_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput162 _12547_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[28] sky130_fd_sc_hd__buf_2
XFILLER_88_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput173 _12038_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[9] sky130_fd_sc_hd__buf_2
XANTENNA__11713__A0 _19958_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11908__B _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16198__S _16200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13615__S _13631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__A _11924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ _11096_/A vssd1 vssd1 vccd1 vccd1 _11342_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ _11046_/A vssd1 vssd1 vccd1 vccd1 _10116_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _11600_/A _11704_/A _12670_/A vssd1 vssd1 vccd1 vccd1 _12641_/A sky130_fd_sc_hd__a21oi_2
XFILLER_43_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ _17542_/A _18098_/B _12551_/B vssd1 vssd1 vccd1 vccd1 _12572_/B sky130_fd_sc_hd__a21o_1
XFILLER_169_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14310_ _14367_/S vssd1 vssd1 vccd1 vccd1 _14319_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_169_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11522_ _11471_/X _11535_/A _11521_/Y vssd1 vssd1 vccd1 vccd1 _11534_/B sky130_fd_sc_hd__a21o_4
X_15290_ _19158_/Q _15289_/X hold9/A vssd1 vssd1 vccd1 vccd1 _15291_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14241_ _14241_/A vssd1 vssd1 vccd1 vccd1 _18737_/D sky130_fd_sc_hd__clkbuf_1
X_11453_ _11452_/A _11450_/Y _11452_/Y _10757_/A vssd1 vssd1 vccd1 vccd1 _11453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14493__A1_N _18328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ _19503_/Q _18915_/Q _18952_/Q _18526_/Q _09651_/A _10440_/A vssd1 vssd1 vccd1
+ vccd1 _10404_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14172_ _13777_/X _18707_/Q _14174_/S vssd1 vssd1 vccd1 vccd1 _14173_/A sky130_fd_sc_hd__mux2_1
X_11384_ _18680_/Q _19175_/Q _11384_/S vssd1 vssd1 vccd1 vccd1 _11385_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10755__A1 _10703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13123_ _19712_/Q _12719_/X _12723_/X _19680_/Q _13122_/X vssd1 vssd1 vccd1 vccd1
+ _15693_/C sky130_fd_sc_hd__a221o_2
X_10335_ _10335_/A _10335_/B vssd1 vssd1 vccd1 vccd1 _10335_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14181__S _14185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18980_ _19366_/CLK _18980_/D vssd1 vssd1 vccd1 vccd1 _18980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _13054_/A _16206_/A vssd1 vssd1 vccd1 vccd1 _13054_/Y sky130_fd_sc_hd__nand2_1
X_17931_ _17929_/Y _17930_/X _17931_/S vssd1 vssd1 vccd1 vccd1 _17931_/X sky130_fd_sc_hd__mux2_1
X_10266_ _10266_/A vssd1 vssd1 vccd1 vccd1 _10439_/S sky130_fd_sc_hd__buf_4
XFILLER_87_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10507__A1 _09749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output155_A _12375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12005_ _11818_/X _11819_/X _12003_/A vssd1 vssd1 vccd1 vccd1 _12005_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17862_ _17666_/S _17716_/X _17632_/X vssd1 vssd1 vccd1 vccd1 _17862_/Y sky130_fd_sc_hd__o21bai_2
X_10197_ _18689_/Q _19184_/Q _10197_/S vssd1 vssd1 vccd1 vccd1 _10197_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16643__B1 _16624_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19601_ _19601_/CLK _19601_/D vssd1 vssd1 vccd1 vccd1 _19601_/Q sky130_fd_sc_hd__dfxtp_1
X_16813_ _16812_/A _16812_/B _18365_/A vssd1 vssd1 vccd1 vccd1 _16814_/B sky130_fd_sc_hd__a21o_1
XFILLER_93_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17793_ _17791_/X _17786_/Y _17792_/Y vssd1 vssd1 vccd1 vccd1 _17793_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19532_ _19988_/CLK _19532_/D vssd1 vssd1 vccd1 vccd1 _19532_/Q sky130_fd_sc_hd__dfxtp_2
X_16744_ _16747_/B _16747_/C _16723_/X vssd1 vssd1 vccd1 vccd1 _16744_/Y sky130_fd_sc_hd__a21oi_1
X_13956_ _13956_/A vssd1 vssd1 vccd1 vccd1 _18614_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10366__S0 _09505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12649__B _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19463_ _19557_/CLK _19463_/D vssd1 vssd1 vccd1 vccd1 _19463_/Q sky130_fd_sc_hd__dfxtp_1
X_12907_ _12893_/A _17122_/A _12880_/X _12883_/X _12906_/X vssd1 vssd1 vccd1 vccd1
+ _19770_/D sky130_fd_sc_hd__o32a_1
X_13887_ _13793_/X _18584_/Q _13889_/S vssd1 vssd1 vccd1 vccd1 _13888_/A sky130_fd_sc_hd__mux2_1
X_16675_ _19666_/Q _16672_/B _16674_/Y vssd1 vssd1 vccd1 vccd1 _19666_/D sky130_fd_sc_hd__o21a_1
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15740__S _15747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18414_ _18414_/A vssd1 vssd1 vccd1 vccd1 _18414_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15626_ _15626_/A vssd1 vssd1 vccd1 vccd1 _19305_/D sky130_fd_sc_hd__clkbuf_1
X_12838_ _12911_/A vssd1 vssd1 vccd1 vccd1 _13204_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19394_ _19394_/CLK _19394_/D vssd1 vssd1 vccd1 vccd1 _19394_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10118__S0 _10753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18345_ _18345_/A _18345_/B vssd1 vssd1 vccd1 vccd1 _18345_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15557_ _19275_/Q _15254_/X _15561_/S vssd1 vssd1 vccd1 vccd1 _15558_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12769_ _12853_/A vssd1 vssd1 vccd1 vccd1 _12903_/A sky130_fd_sc_hd__buf_2
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12665__A _12669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13260__S _13278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14508_ _14508_/A vssd1 vssd1 vccd1 vccd1 _18833_/D sky130_fd_sc_hd__clkbuf_1
X_15488_ _15488_/A vssd1 vssd1 vccd1 vccd1 _19244_/D sky130_fd_sc_hd__clkbuf_1
X_18276_ _18276_/A _18345_/B vssd1 vssd1 vccd1 vccd1 _18276_/X sky130_fd_sc_hd__or2_1
Xinput20 io_dbus_rdata[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_4
X_17227_ _17225_/Y _17212_/X _17226_/X _17215_/X vssd1 vssd1 vccd1 vccd1 _19842_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14439_ _14439_/A vssd1 vssd1 vccd1 vccd1 _18815_/D sky130_fd_sc_hd__clkbuf_1
Xinput31 io_dbus_rdata[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_2
XANTENNA__14880__A _14902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18352__A _18352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput42 io_ibus_inst[17] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 io_ibus_inst[27] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_2
Xinput64 io_ibus_inst[8] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17158_ _13595_/A _17164_/B _17123_/A vssd1 vssd1 vccd1 vccd1 _17158_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16109_ _13376_/X _19472_/Q _16117_/S vssd1 vssd1 vccd1 vccd1 _16110_/A sky130_fd_sc_hd__mux2_1
X_09980_ _11378_/A vssd1 vssd1 vccd1 vccd1 _10732_/A sky130_fd_sc_hd__clkbuf_2
X_17089_ _17089_/A _17089_/B _17089_/C vssd1 vssd1 vccd1 vccd1 _19791_/D sky130_fd_sc_hd__nor3_1
XFILLER_89_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10841__S1 _09985_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10913__A _11035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_147_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13160__A2 _13157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15216__A _15299_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__S0 _10337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09414_ _13748_/B vssd1 vssd1 vccd1 vccd1 _16208_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__17431__A _17431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ _19894_/Q vssd1 vssd1 vccd1 vccd1 _09345_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__14266__S _14268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17150__B _17229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16047__A _16047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10434__B1 _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09276_ _09307_/B _09215_/A _09215_/B _11608_/A _09275_/X vssd1 vssd1 vccd1 vccd1
+ _09277_/D sky130_fd_sc_hd__o2111a_1
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11529__A3 _11534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15097__S _15105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10120_ _18790_/Q _19061_/Q _19285_/Q _19029_/Q _10119_/X _10054_/A vssd1 vssd1 vccd1
+ vccd1 _10120_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10051_ _10051_/A vssd1 vssd1 vccd1 vccd1 _10790_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16625__B1 _16624_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13853__B _14501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13439__B1 _19950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13810_ _13809_/X _18557_/Q _13813_/S vssd1 vssd1 vccd1 vccd1 _13811_/A sky130_fd_sc_hd__mux2_1
X_14790_ _14790_/A vssd1 vssd1 vccd1 vccd1 _18948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13741_ _13741_/A vssd1 vssd1 vccd1 vccd1 _18537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10953_ _11250_/A _10953_/B vssd1 vssd1 vccd1 vccd1 _10953_/X sky130_fd_sc_hd__or2_1
XFILLER_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17050__B1 _17021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13672_ _14621_/A vssd1 vssd1 vccd1 vccd1 _13672_/X sky130_fd_sc_hd__clkbuf_2
X_16460_ _11986_/A _11986_/B _16455_/X vssd1 vssd1 vccd1 vccd1 _19585_/D sky130_fd_sc_hd__a21o_1
X_10884_ _11478_/A _10877_/X _10883_/X _09975_/A vssd1 vssd1 vccd1 vccd1 _10885_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15411_ _14628_/X _19210_/Q _15417_/S vssd1 vssd1 vccd1 vccd1 _15412_/A sky130_fd_sc_hd__mux2_1
X_12623_ _12395_/S _12622_/X _11871_/X vssd1 vssd1 vccd1 vccd1 _12623_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16391_ _13178_/X _19554_/Q _16393_/S vssd1 vssd1 vccd1 vccd1 _16392_/A sky130_fd_sc_hd__mux2_1
X_15342_ _15342_/A vssd1 vssd1 vccd1 vccd1 _19179_/D sky130_fd_sc_hd__clkbuf_1
X_18130_ _19926_/Q _19958_/Q _18136_/S vssd1 vssd1 vccd1 vccd1 _18131_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12554_ _12556_/A _18097_/B vssd1 vssd1 vccd1 vccd1 _12555_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10520__S0 _10470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17487__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ _19386_/Q _19000_/Q _19450_/Q _18569_/Q _10119_/X _10112_/A vssd1 vssd1 vccd1
+ vccd1 _11506_/B sky130_fd_sc_hd__mux4_1
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15273_ _15273_/A vssd1 vssd1 vccd1 vccd1 _15273_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18061_ _17781_/X _17764_/X _18060_/X _17940_/X vssd1 vssd1 vccd1 vccd1 _18061_/X
+ sky130_fd_sc_hd__a211o_1
X_12485_ _12520_/A _12485_/B vssd1 vssd1 vccd1 vccd1 _12485_/Y sky130_fd_sc_hd__xnor2_4
X_14224_ _14502_/A _16371_/D vssd1 vssd1 vccd1 vccd1 _14281_/A sky130_fd_sc_hd__or2_4
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17012_ _17016_/C _17013_/C _19761_/Q vssd1 vssd1 vccd1 vccd1 _17014_/B sky130_fd_sc_hd__a21oi_1
XFILLER_171_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11436_ _09476_/A _11427_/X _11431_/X _11435_/X _10623_/A vssd1 vssd1 vccd1 vccd1
+ _11436_/X sky130_fd_sc_hd__a311o_1
XFILLER_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11076__S1 _11065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14155_ _13746_/X _18699_/Q _14163_/S vssd1 vssd1 vccd1 vccd1 _14156_/A sky130_fd_sc_hd__mux2_1
X_11367_ _19465_/Q _19303_/Q _18712_/Q _18482_/Q _10675_/X _10609_/X vssd1 vssd1 vccd1
+ vccd1 _11367_/X sky130_fd_sc_hd__mux4_2
XFILLER_4_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13106_ _19898_/Q _15686_/B _13430_/S vssd1 vssd1 vccd1 vccd1 _13106_/X sky130_fd_sc_hd__mux2_1
X_10318_ _18655_/Q _19246_/Q _19408_/Q _18623_/Q _09505_/A _10312_/X vssd1 vssd1 vccd1
+ vccd1 _10318_/X sky130_fd_sc_hd__mux4_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14086_ _14086_/A vssd1 vssd1 vccd1 vccd1 _18670_/D sky130_fd_sc_hd__clkbuf_1
X_18963_ _19288_/CLK _18963_/D vssd1 vssd1 vccd1 vccd1 _18963_/Q sky130_fd_sc_hd__dfxtp_1
X_11298_ _11291_/Y _11293_/Y _11295_/Y _11297_/Y _10994_/A vssd1 vssd1 vccd1 vccd1
+ _11298_/X sky130_fd_sc_hd__o221a_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _18929_/Q vssd1 vssd1 vccd1 vccd1 _13038_/A sky130_fd_sc_hd__clkbuf_2
X_17914_ _17914_/A _17914_/B vssd1 vssd1 vccd1 vccd1 _17914_/Y sky130_fd_sc_hd__nor2_1
X_10249_ _18592_/Q _18853_/Q _18752_/Q _19087_/Q _09901_/A _09842_/A vssd1 vssd1 vccd1
+ vccd1 _10250_/B sky130_fd_sc_hd__mux4_1
XFILLER_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18894_ _19203_/CLK _18894_/D vssd1 vssd1 vccd1 vccd1 _18894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17845_ _17845_/A _17845_/B vssd1 vssd1 vccd1 vccd1 _17845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17776_ _17953_/A vssd1 vssd1 vccd1 vccd1 _17776_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14988_ _14988_/A vssd1 vssd1 vccd1 vccd1 _19033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19515_ _19577_/CLK _19515_/D vssd1 vssd1 vccd1 vccd1 _19515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16727_ _19680_/Q _16727_/B _16727_/C vssd1 vssd1 vccd1 vccd1 _16728_/C sky130_fd_sc_hd__and3_1
X_13939_ _18607_/Q _13630_/X _13939_/S vssd1 vssd1 vccd1 vccd1 _13940_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15470__S _15478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18347__A _18347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19446_ _19510_/CLK _19446_/D vssd1 vssd1 vccd1 vccd1 _19446_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09969__A _10074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16658_ _19660_/Q _16655_/B _16657_/Y vssd1 vssd1 vccd1 vccd1 _19660_/D sky130_fd_sc_hd__o21a_1
XFILLER_23_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15609_ _14602_/X _19298_/Q _15611_/S vssd1 vssd1 vccd1 vccd1 _15610_/A sky130_fd_sc_hd__mux2_1
X_19377_ _19377_/CLK _19377_/D vssd1 vssd1 vccd1 vccd1 _19377_/Q sky130_fd_sc_hd__dfxtp_1
X_16589_ _19636_/Q _16590_/C _19637_/Q vssd1 vssd1 vccd1 vccd1 _16591_/B sky130_fd_sc_hd__a21oi_1
XFILLER_148_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_73_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18328_ _18328_/A _18333_/B vssd1 vssd1 vccd1 vccd1 _18328_/X sky130_fd_sc_hd__or2_1
X_18259_ _18259_/A vssd1 vssd1 vccd1 vccd1 _19983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11067__S1 _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10643__A _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _20052_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ _19124_/Q _18890_/Q _19572_/Q _19220_/Q _10811_/S _09515_/A vssd1 vssd1 vccd1
+ vccd1 _09963_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10362__B _12657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17426__A _17581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09894_ _19918_/Q vssd1 vssd1 vccd1 vccd1 _09894_/Y sky130_fd_sc_hd__inv_2
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16607__B1 _16577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15380__S _15384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17161__A _17229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09328_ _18279_/A _18276_/A _09328_/C _09328_/D vssd1 vssd1 vccd1 vccd1 _11789_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10502__S0 _10496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ _09271_/C _11786_/A _11787_/A vssd1 vssd1 vccd1 vccd1 _12601_/B sky130_fd_sc_hd__nand3_2
XANTENNA__14724__S _14724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17886__A2 _17877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12270_ _18319_/A _17334_/B _12190_/X vssd1 vssd1 vccd1 vccd1 _12270_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ _11221_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11221_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11152_ _18575_/Q _18836_/Q _18735_/Q _19070_/Q _10968_/S _10024_/A vssd1 vssd1 vccd1
+ vccd1 _11153_/B sky130_fd_sc_hd__mux4_1
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16310__A2 _15770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15555__S _15561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ _09613_/A _10090_/X _10102_/X _09996_/X _19920_/Q vssd1 vssd1 vccd1 vccd1
+ _10137_/A sky130_fd_sc_hd__a32o_4
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15960_ _19406_/Q _15257_/X _15962_/S vssd1 vssd1 vccd1 vccd1 _15961_/A sky130_fd_sc_hd__mux2_1
X_11083_ _18800_/Q _19135_/Q _11083_/S vssd1 vssd1 vccd1 vccd1 _11083_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11135__B2 _19897_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_A io_dbus_rdata[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ _14669_/X _18999_/Q _14911_/S vssd1 vssd1 vccd1 vccd1 _14912_/A sky130_fd_sc_hd__mux2_1
X_10034_ _10040_/A vssd1 vssd1 vccd1 vccd1 _10751_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__13583__B _17152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15891_ _15891_/A vssd1 vssd1 vccd1 vccd1 _19375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17630_ _17662_/A vssd1 vssd1 vccd1 vccd1 _17741_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_84_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14842_ _18321_/A _16315_/A _14825_/X _14841_/Y vssd1 vssd1 vccd1 vccd1 _18407_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15821__A1 _18464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17561_ _17413_/X _17458_/X _17573_/S vssd1 vssd1 vccd1 vccd1 _17561_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11985_ _11978_/X _11979_/X _11984_/Y _12247_/A vssd1 vssd1 vccd1 vccd1 _11986_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_91_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14773_ _18941_/Q _14398_/X _14775_/S vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output118_A _12655_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19300_ _19430_/CLK _19300_/D vssd1 vssd1 vccd1 vccd1 _19300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16512_ _16520_/D vssd1 vssd1 vccd1 vccd1 _16518_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13724_ _18533_/Q _13723_/X _13736_/S vssd1 vssd1 vccd1 vccd1 _13725_/A sky130_fd_sc_hd__mux2_1
X_10936_ _11190_/A vssd1 vssd1 vccd1 vccd1 _11001_/A sky130_fd_sc_hd__clkbuf_2
X_17492_ _17483_/X _17491_/X _17649_/A vssd1 vssd1 vccd1 vccd1 _17493_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19231_ _19489_/CLK _19231_/D vssd1 vssd1 vccd1 vccd1 _19231_/Q sky130_fd_sc_hd__dfxtp_1
X_16443_ _17319_/A vssd1 vssd1 vccd1 vccd1 _18341_/A sky130_fd_sc_hd__buf_2
XFILLER_158_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13655_ _14608_/A vssd1 vssd1 vccd1 vccd1 _13655_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10867_ _09998_/X _10856_/X _10865_/X _10065_/X _10866_/Y vssd1 vssd1 vccd1 vccd1
+ _12644_/A sky130_fd_sc_hd__o32a_4
XFILLER_20_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19162_ _19392_/CLK _19162_/D vssd1 vssd1 vccd1 vccd1 _19162_/Q sky130_fd_sc_hd__dfxtp_1
X_12606_ _12606_/A _18286_/A _18283_/A _12606_/D vssd1 vssd1 vccd1 vccd1 _12610_/C
+ sky130_fd_sc_hd__or4_1
XANTENNA__12938__A2 _09464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _13586_/A vssd1 vssd1 vccd1 vccd1 _18503_/D sky130_fd_sc_hd__clkbuf_1
X_16374_ _13009_/X _19546_/Q _16382_/S vssd1 vssd1 vccd1 vccd1 _16375_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _10783_/X _10788_/X _10797_/X _10063_/X vssd1 vssd1 vccd1 vccd1 _10798_/X
+ sky130_fd_sc_hd__a22o_2
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _17697_/X _18110_/X _18112_/Y _17634_/X vssd1 vssd1 vccd1 vccd1 _18113_/X
+ sky130_fd_sc_hd__o211a_1
X_15325_ _15371_/S vssd1 vssd1 vccd1 vccd1 _15334_/S sky130_fd_sc_hd__buf_2
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12537_ _12537_/A vssd1 vssd1 vccd1 vccd1 _12537_/X sky130_fd_sc_hd__buf_2
XFILLER_145_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19093_ _19317_/CLK _19093_/D vssd1 vssd1 vccd1 vccd1 _19093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13348__C1 _13347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18044_ _18046_/A _18046_/B _18077_/S vssd1 vssd1 vccd1 vccd1 _18044_/X sky130_fd_sc_hd__mux2_1
X_15256_ _15256_/A vssd1 vssd1 vccd1 vccd1 _19147_/D sky130_fd_sc_hd__clkbuf_1
X_12468_ _19539_/Q _12206_/X _12262_/X _12467_/X _12123_/X vssd1 vssd1 vccd1 vccd1
+ _12468_/X sky130_fd_sc_hd__o221a_1
XANTENNA__12662__B _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14207_ _13828_/X _18723_/Q _14207_/S vssd1 vssd1 vccd1 vccd1 _14208_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11419_ _11554_/B vssd1 vssd1 vccd1 vccd1 _11419_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18287__C1 _17243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15187_ _19125_/Q vssd1 vssd1 vccd1 vccd1 _15188_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_153_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12399_ _19839_/Q _12419_/C vssd1 vssd1 vccd1 vccd1 _12399_/X sky130_fd_sc_hd__and2_1
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16837__B1 _16833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14138_ _18694_/Q _13727_/X _14142_/S vssd1 vssd1 vccd1 vccd1 _14139_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19995_ _20027_/CLK _19995_/D vssd1 vssd1 vccd1 vccd1 _19995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13774__A _14599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ _14069_/A vssd1 vssd1 vccd1 vccd1 _18664_/D sky130_fd_sc_hd__clkbuf_1
X_18946_ _19369_/CLK _18946_/D vssd1 vssd1 vccd1 vccd1 _18946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18877_ _19559_/CLK _18877_/D vssd1 vssd1 vccd1 vccd1 _18877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17828_ _17729_/A _17763_/X _17719_/A vssd1 vssd1 vccd1 vccd1 _17828_/X sky130_fd_sc_hd__o21ba_1
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15812__A1 _18463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17759_ _17654_/B _17647_/X _17759_/S vssd1 vssd1 vccd1 vccd1 _17759_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12626__A1 _17240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12837__B _12837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19429_ _19555_/CLK _19429_/D vssd1 vssd1 vccd1 vccd1 _19429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13014__A _14844_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14544__S _14546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__A _12853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_150_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19726_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12562__A0 _12559_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13684__A _15254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17156__A _19819_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09946_ _10144_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_165_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19782_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09877_ _18788_/Q _19059_/Q _19283_/Q _19027_/Q _10173_/S _09887_/A vssd1 vssd1 vccd1
+ vccd1 _09877_/X sky130_fd_sc_hd__mux4_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13623__S _13631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _16487_/A vssd1 vssd1 vccd1 vccd1 _12628_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16219__B _16219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17556__B2 _12946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _19464_/Q _19302_/Q _18711_/Q _18481_/Q _10644_/X _10645_/X vssd1 vssd1 vccd1
+ vccd1 _10721_/X sky130_fd_sc_hd__mux4_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _13460_/B _13439_/Y _11607_/X vssd1 vssd1 vccd1 vccd1 _13440_/Y sky130_fd_sc_hd__o21ai_1
X_10652_ _10652_/A vssd1 vssd1 vccd1 vccd1 _10768_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_103_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19514_/CLK sky130_fd_sc_hd__clkbuf_16
X_13371_ _13371_/A vssd1 vssd1 vccd1 vccd1 _13483_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14454__S _14466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10583_ _10583_/A _10583_/B vssd1 vssd1 vccd1 vccd1 _10583_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15110_ _14644_/X _19087_/Q _15116_/S vssd1 vssd1 vccd1 vccd1 _15111_/A sky130_fd_sc_hd__mux2_1
X_12322_ _12322_/A vssd1 vssd1 vccd1 vccd1 _18001_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16090_ _16090_/A vssd1 vssd1 vccd1 vccd1 _19463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15041_ _15041_/A vssd1 vssd1 vccd1 vccd1 _19056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12253_ _17945_/B _12225_/B _17389_/A vssd1 vssd1 vccd1 vccd1 _12254_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__10283__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_118_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19553_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11204_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11204_/X sky130_fd_sc_hd__or2_1
XFILLER_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12184_ _17192_/A _12217_/C vssd1 vssd1 vccd1 vccd1 _12184_/X sky130_fd_sc_hd__or2_1
X_18800_ _19491_/CLK _18800_/D vssd1 vssd1 vccd1 vccd1 _18800_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17066__A _17066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ _09611_/A _11123_/X _11134_/X _09619_/A _19897_/Q vssd1 vssd1 vccd1 vccd1
+ _11135_/X sky130_fd_sc_hd__a32o_4
XANTENNA_clkbuf_leaf_21_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19780_ _19783_/CLK _19780_/D vssd1 vssd1 vccd1 vccd1 _19780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16992_ _19755_/Q _16994_/C _16992_/C vssd1 vssd1 vccd1 vccd1 _16993_/C sky130_fd_sc_hd__and3_1
XANTENNA__11108__A1 _09745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ _19389_/CLK _18731_/D vssd1 vssd1 vccd1 vccd1 _18731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15943_ _19398_/Q _15231_/X _15951_/S vssd1 vssd1 vccd1 vccd1 _15944_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11066_ _18768_/Q _19039_/Q _19263_/Q _19007_/Q _11000_/S _11065_/X vssd1 vssd1 vccd1
+ vccd1 _11066_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11203__S1 _09511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10017_ _10017_/A vssd1 vssd1 vccd1 vccd1 _10018_/A sky130_fd_sc_hd__clkbuf_4
X_18662_ _19511_/CLK _18662_/D vssd1 vssd1 vccd1 vccd1 _18662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15874_ _15874_/A vssd1 vssd1 vccd1 vccd1 _19367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17613_ _17607_/X _17616_/B _17611_/X _17612_/X vssd1 vssd1 vccd1 vccd1 _17613_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_28_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14825_ _14831_/A vssd1 vssd1 vccd1 vccd1 _14825_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12608__A1 _18302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18593_ _19476_/CLK _18593_/D vssd1 vssd1 vccd1 vccd1 _18593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14629__S _14638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11842__A _19820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15314__A _15371_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17544_ _12673_/A _17748_/S _17541_/X _17543_/X vssd1 vssd1 vccd1 vccd1 _17544_/X
+ sky130_fd_sc_hd__a211o_1
X_14756_ _18933_/Q _14369_/X _14764_/S vssd1 vssd1 vccd1 vccd1 _14757_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11968_ _11968_/A _17412_/A vssd1 vssd1 vccd1 vccd1 _11971_/A sky130_fd_sc_hd__xor2_2
XANTENNA__12657__B _12657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09312__A _20041_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ _18529_/Q _13706_/X _13715_/S vssd1 vssd1 vccd1 vccd1 _13708_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17475_ _17507_/S vssd1 vssd1 vccd1 vccd1 _17506_/S sky130_fd_sc_hd__clkbuf_2
X_10919_ _18830_/Q vssd1 vssd1 vccd1 vccd1 _10920_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10458__A _10459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14687_ _18898_/Q _14379_/X _14691_/S vssd1 vssd1 vccd1 vccd1 _14688_/A sky130_fd_sc_hd__mux2_1
X_11899_ _11961_/A _11899_/B vssd1 vssd1 vccd1 vccd1 _11899_/X sky130_fd_sc_hd__or2_1
X_19214_ _19311_/CLK _19214_/D vssd1 vssd1 vccd1 vccd1 _19214_/Q sky130_fd_sc_hd__dfxtp_1
X_16426_ _13433_/X _19570_/Q _16426_/S vssd1 vssd1 vccd1 vccd1 _16427_/A sky130_fd_sc_hd__mux2_1
X_13638_ _15219_/A vssd1 vssd1 vccd1 vccd1 _14596_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_158_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19145_ _19405_/CLK _19145_/D vssd1 vssd1 vccd1 vccd1 _19145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16357_ _16361_/A _16361_/C vssd1 vssd1 vccd1 vccd1 _16357_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13569_ _18437_/Q _13569_/B vssd1 vssd1 vccd1 vccd1 _13569_/X sky130_fd_sc_hd__or2_1
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15308_ _19164_/Q _15206_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _15309_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19076_ _19430_/CLK _19076_/D vssd1 vssd1 vccd1 vccd1 _19076_/Q sky130_fd_sc_hd__dfxtp_1
X_16288_ _16288_/A vssd1 vssd1 vccd1 vccd1 _19529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17675__S _17675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15730__A0 _19904_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18027_ _17928_/X _17828_/X _18026_/X _17953_/X vssd1 vssd1 vccd1 vccd1 _18027_/X
+ sky130_fd_sc_hd__o211a_1
X_15239_ _19142_/Q _15238_/X _15245_/S vssd1 vssd1 vccd1 vccd1 _15240_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11347__A1 _11302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12544__B1 _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11347__B2 _12631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09982__A _11305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11442__S1 _10813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09800_ _09800_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09800_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_82_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19302_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12612__S _12612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19978_ _19978_/CLK _19978_/D vssd1 vssd1 vccd1 vccd1 _19978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09731_ _18794_/Q _19065_/Q _19289_/Q _19033_/Q _09726_/S _09730_/X vssd1 vssd1 vccd1
+ vccd1 _09731_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18929_ _19954_/CLK _18929_/D vssd1 vssd1 vccd1 vccd1 _18929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15923__S _15929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09662_ _09662_/A vssd1 vssd1 vccd1 vccd1 _10703_/A sky130_fd_sc_hd__buf_6
XANTENNA__13009__A _15197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_97_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19559_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09593_ _09777_/A _09592_/X _09479_/X vssd1 vssd1 vccd1 vccd1 _09593_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09571__S0 _09761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19978_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10368__A _10368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11130__S0 _11129_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19564_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_108_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17710__A1 _19896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11199__A _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11433__S1 _10813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17474__A0 _12385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09929_ _09929_/A vssd1 vssd1 vccd1 vccd1 _09929_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20049_ _20049_/CLK _20049_/D vssd1 vssd1 vccd1 vccd1 _20049_/Q sky130_fd_sc_hd__dfxtp_2
X_12940_ _18440_/Q _12939_/X _17808_/S vssd1 vssd1 vccd1 vccd1 _12941_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10944__S0 _11305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _19654_/Q _12727_/X _12729_/X _19786_/Q _12870_/X vssd1 vssd1 vccd1 vccd1
+ _12872_/B sky130_fd_sc_hd__a221o_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _14608_/X _18874_/Q _14622_/S vssd1 vssd1 vccd1 vccd1 _14611_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11822_ _11976_/B vssd1 vssd1 vccd1 vccd1 _12088_/B sky130_fd_sc_hd__clkbuf_2
X_15590_ _15646_/A vssd1 vssd1 vccd1 vccd1 _15659_/S sky130_fd_sc_hd__buf_4
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17529__A1 _17542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _14541_/A vssd1 vssd1 vccd1 vccd1 _18848_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _20038_/Q vssd1 vssd1 vccd1 vccd1 _18316_/A sky130_fd_sc_hd__buf_4
XFILLER_42_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10704_ _11046_/A vssd1 vssd1 vccd1 vccd1 _11510_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17317_/S vssd1 vssd1 vccd1 vccd1 _17269_/S sky130_fd_sc_hd__buf_2
XFILLER_41_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14472_ _18826_/Q _14471_/X _14472_/S vssd1 vssd1 vccd1 vccd1 _14473_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15788__B _18459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11684_ _11684_/A vssd1 vssd1 vccd1 vccd1 _17325_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16211_ _19516_/Q _16207_/Y _16223_/S vssd1 vssd1 vccd1 vccd1 _16212_/A sky130_fd_sc_hd__mux2_1
X_10635_ _10627_/X _10629_/X _10632_/X _10634_/X _09603_/A vssd1 vssd1 vccd1 vccd1
+ _10635_/X sky130_fd_sc_hd__a221o_1
X_13423_ _15273_/A vssd1 vssd1 vccd1 vccd1 _13423_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17191_ _17191_/A vssd1 vssd1 vccd1 vccd1 _17191_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16142_ _16142_/A vssd1 vssd1 vccd1 vccd1 _19486_/D sky130_fd_sc_hd__clkbuf_1
X_13354_ _13354_/A vssd1 vssd1 vccd1 vccd1 _13354_/X sky130_fd_sc_hd__clkbuf_2
X_10566_ _10571_/A _10563_/X _10565_/X _09577_/A vssd1 vssd1 vccd1 vccd1 _10566_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ _12332_/A _12331_/A vssd1 vssd1 vccd1 vccd1 _12306_/B sky130_fd_sc_hd__or2_1
XFILLER_115_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13285_ _19339_/Q _12802_/A _12704_/A _19529_/Q _13284_/X vssd1 vssd1 vccd1 vccd1
+ _13285_/X sky130_fd_sc_hd__a221o_1
X_16073_ _13089_/X _19456_/Q _16073_/S vssd1 vssd1 vccd1 vccd1 _16074_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10497_ _10497_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10497_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15024_ _15046_/A vssd1 vssd1 vccd1 vccd1 _15033_/S sky130_fd_sc_hd__clkbuf_4
X_12236_ _19584_/Q _19585_/Q _19588_/Q _19589_/Q vssd1 vssd1 vccd1 vccd1 _12237_/D
+ sky130_fd_sc_hd__and4_1
X_19901_ _19971_/CLK _19901_/D vssd1 vssd1 vccd1 vccd1 _19901_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17465__A0 _17866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19832_ _19865_/CLK _19832_/D vssd1 vssd1 vccd1 vccd1 _19832_/Q sky130_fd_sc_hd__dfxtp_1
X_12167_ _19971_/Q _10672_/A _12303_/S vssd1 vssd1 vccd1 vccd1 _17444_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11118_ _11001_/A _11111_/X _11115_/X _11117_/X vssd1 vssd1 vccd1 vccd1 _11118_/X
+ sky130_fd_sc_hd__a211o_1
X_19763_ _19768_/CLK _19763_/D vssd1 vssd1 vccd1 vccd1 _19763_/Q sky130_fd_sc_hd__dfxtp_1
X_16975_ _19750_/Q _19749_/Q _19748_/Q _16975_/D vssd1 vssd1 vccd1 vccd1 _16984_/D
+ sky130_fd_sc_hd__and4_1
X_12098_ _12098_/A vssd1 vssd1 vccd1 vccd1 _12189_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18714_ _19305_/CLK _18714_/D vssd1 vssd1 vccd1 vccd1 _18714_/Q sky130_fd_sc_hd__dfxtp_1
X_15926_ _15926_/A vssd1 vssd1 vccd1 vccd1 _19390_/D sky130_fd_sc_hd__clkbuf_1
X_11049_ _11042_/Y _11044_/Y _11046_/Y _11048_/Y _10063_/A vssd1 vssd1 vccd1 vccd1
+ _11049_/X sky130_fd_sc_hd__o221a_1
X_19694_ _19726_/CLK _19694_/D vssd1 vssd1 vccd1 vccd1 _19694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 io_dbus_rdata[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_4
XFILLER_77_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18645_ _19268_/CLK _18645_/D vssd1 vssd1 vccd1 vccd1 _18645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15857_ _13089_/X _19360_/Q _15857_/S vssd1 vssd1 vccd1 vccd1 _15858_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14359__S _14363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12668__A _12669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14808_ _18957_/Q _14449_/X _14808_/S vssd1 vssd1 vccd1 vccd1 _14809_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18576_ _19293_/CLK _18576_/D vssd1 vssd1 vccd1 vccd1 _18576_/Q sky130_fd_sc_hd__dfxtp_1
X_15788_ _15811_/A _18459_/Q vssd1 vssd1 vccd1 vccd1 _15788_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17527_ _17690_/A _17527_/B vssd1 vssd1 vccd1 vccd1 _17719_/A sky130_fd_sc_hd__nor2_1
X_14739_ _14739_/A vssd1 vssd1 vccd1 vccd1 _18921_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18355__A _18365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17458_ _17820_/B _12407_/A _17460_/S vssd1 vssd1 vccd1 vccd1 _17458_/X sky130_fd_sc_hd__mux2_1
X_16409_ _13309_/X _19562_/Q _16415_/S vssd1 vssd1 vccd1 vccd1 _16410_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14094__S _14098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10916__A _10978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17389_ _17389_/A vssd1 vssd1 vccd1 vccd1 _17721_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19128_ _19203_/CLK _19128_/D vssd1 vssd1 vccd1 vccd1 _19128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19059_ _19287_/CLK _19059_/D vssd1 vssd1 vccd1 vccd1 _19059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10528__C1 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15219__A _15219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15653__S _15655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ _18831_/Q vssd1 vssd1 vccd1 vccd1 _10994_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09697__B1 _09696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10926__S0 _10909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09645_ _11495_/S vssd1 vssd1 vccd1 vccd1 _10849_/S sky130_fd_sc_hd__buf_4
XFILLER_55_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11482__A _11482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09576_ _10621_/A vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__buf_6
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10154__S1 _10148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09887__A _09887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ _18781_/Q _19052_/Q _19276_/Q _19020_/Q _10465_/S _10291_/X vssd1 vssd1 vccd1
+ vccd1 _10420_/X sky130_fd_sc_hd__mux4_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10351_ _10583_/A vssd1 vssd1 vccd1 vccd1 _10490_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ _18472_/Q _13069_/X _13090_/S vssd1 vssd1 vccd1 vccd1 _13071_/A sky130_fd_sc_hd__mux2_1
X_10282_ _18656_/Q _19247_/Q _19409_/Q _18624_/Q _10173_/S _09887_/A vssd1 vssd1 vccd1
+ vccd1 _10283_/B sky130_fd_sc_hd__mux4_1
XFILLER_117_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12021_ _12021_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12023_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16760_ _19691_/Q _16763_/C _16723_/X vssd1 vssd1 vccd1 vccd1 _16760_/Y sky130_fd_sc_hd__a21oi_1
X_13972_ _18622_/Q _13693_/X _13972_/S vssd1 vssd1 vccd1 vccd1 _13973_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10298__A1 _09520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15711_ _13568_/X _15709_/X _15710_/Y _13577_/X _18445_/Q vssd1 vssd1 vccd1 vccd1
+ _17175_/A sky130_fd_sc_hd__a32oi_4
XANTENNA__09783__S0 _09724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13591__B _13591_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ _18461_/Q _12921_/X _12922_/Y _13580_/A vssd1 vssd1 vccd1 vccd1 _12923_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14179__S _14185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16691_ _16728_/A _16691_/B _16691_/C vssd1 vssd1 vccd1 vccd1 _19671_/D sky130_fd_sc_hd__nor3_1
X_18430_ input57/X vssd1 vssd1 vccd1 vccd1 _18430_/Y sky130_fd_sc_hd__inv_2
X_15642_ _14650_/X _19313_/Q _15644_/S vssd1 vssd1 vccd1 vccd1 _15643_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _12735_/X _12851_/X _12852_/Y _12853_/X _18448_/Q vssd1 vssd1 vccd1 vccd1
+ _12854_/X sky130_fd_sc_hd__a32o_4
XFILLER_92_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ input59/X vssd1 vssd1 vccd1 vccd1 _18361_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15799__A _15799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11805_ _12634_/B _11804_/X _11856_/S vssd1 vssd1 vccd1 vccd1 _11849_/D sky130_fd_sc_hd__mux2_1
X_15573_ _15573_/A vssd1 vssd1 vccd1 vccd1 _19282_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output100_A _11972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14907__S _14911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _19628_/Q _13142_/B _12784_/X vssd1 vssd1 vccd1 vccd1 _12785_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _17312_/A vssd1 vssd1 vccd1 vccd1 _19878_/D sky130_fd_sc_hd__clkbuf_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14524_ _13780_/X _18841_/Q _14524_/S vssd1 vssd1 vccd1 vccd1 _14525_/A sky130_fd_sc_hd__mux2_1
X_18292_ _18335_/A vssd1 vssd1 vccd1 vccd1 _18326_/B sky130_fd_sc_hd__buf_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _12097_/A _12631_/B _11735_/Y vssd1 vssd1 vccd1 vccd1 _17414_/A sky130_fd_sc_hd__a21oi_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _18289_/A vssd1 vssd1 vccd1 vccd1 _17243_/X sky130_fd_sc_hd__buf_2
XFILLER_174_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14455_ _14455_/A vssd1 vssd1 vccd1 vccd1 _18820_/D sky130_fd_sc_hd__clkbuf_1
X_11667_ input66/X _12857_/A vssd1 vssd1 vccd1 vccd1 _11797_/A sky130_fd_sc_hd__nand2_1
X_13406_ _16923_/C _13341_/X _13342_/X _19696_/Q _13405_/X vssd1 vssd1 vccd1 vccd1
+ _13406_/X sky130_fd_sc_hd__a221o_1
X_10618_ _10618_/A vssd1 vssd1 vccd1 vccd1 _10682_/A sky130_fd_sc_hd__buf_4
X_17174_ _17141_/A _17167_/X _17173_/X _17171_/X vssd1 vssd1 vccd1 vccd1 _19824_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11598_ _11535_/Y _11537_/X _11538_/X _11534_/B _11597_/X vssd1 vssd1 vccd1 vccd1
+ _11598_/X sky130_fd_sc_hd__a221o_4
XANTENNA__17135__C1 _16480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14386_ _18799_/Q _14385_/X _14386_/S vssd1 vssd1 vccd1 vccd1 _14387_/A sky130_fd_sc_hd__mux2_1
X_16125_ _16125_/A vssd1 vssd1 vccd1 vccd1 _19479_/D sky130_fd_sc_hd__clkbuf_1
X_10549_ _19468_/Q _19306_/Q _18715_/Q _18485_/Q _10266_/A _10592_/A vssd1 vssd1 vccd1
+ vccd1 _10549_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13337_ _13337_/A vssd1 vssd1 vccd1 vccd1 _13337_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14642__S _14654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12951__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16056_ _13523_/X _19449_/Q _16056_/S vssd1 vssd1 vccd1 vccd1 _16057_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13268_ _16920_/B _12989_/X _12990_/X _19688_/Q _13267_/X vssd1 vssd1 vccd1 vccd1
+ _13268_/X sky130_fd_sc_hd__a221o_2
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12670__B _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15007_ _19041_/Q _14395_/X _15011_/S vssd1 vssd1 vccd1 vccd1 _15008_/A sky130_fd_sc_hd__mux2_1
X_12219_ _12215_/X _12216_/Y _12267_/C _12218_/X vssd1 vssd1 vccd1 vccd1 _12219_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_123_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13199_ _19652_/Q vssd1 vssd1 vccd1 vccd1 _16636_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19815_ _19852_/CLK _19815_/D vssd1 vssd1 vccd1 vccd1 _19815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19746_ _19756_/CLK _19746_/D vssd1 vssd1 vccd1 vccd1 _19746_/Q sky130_fd_sc_hd__dfxtp_1
X_16958_ _16958_/A _16958_/B _16964_/A _16958_/D vssd1 vssd1 vccd1 vccd1 _16959_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_110_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15909_ _15909_/A vssd1 vssd1 vccd1 vccd1 _19383_/D sky130_fd_sc_hd__clkbuf_1
X_19677_ _19682_/CLK _19677_/D vssd1 vssd1 vccd1 vccd1 _19677_/Q sky130_fd_sc_hd__dfxtp_1
X_16889_ _16897_/A _16889_/B _16896_/D vssd1 vssd1 vccd1 vccd1 _19727_/D sky130_fd_sc_hd__nor3_1
XFILLER_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09430_ _20042_/Q vssd1 vssd1 vccd1 vccd1 _17339_/A sky130_fd_sc_hd__clkbuf_2
X_18628_ _19569_/CLK _18628_/D vssd1 vssd1 vccd1 vccd1 _18628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13227__B2 _13418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09361_ _09398_/A _09398_/B _20010_/Q _20009_/Q vssd1 vssd1 vccd1 vccd1 _12711_/A
+ sky130_fd_sc_hd__or4b_2
XANTENNA__11238__B1 _10941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18559_ _19311_/CLK _18559_/D vssd1 vssd1 vccd1 vccd1 _18559_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14817__S _14819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__S0 _11035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_143_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15502__A _15502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09292_ _20040_/Q _14074_/A vssd1 vssd1 vccd1 vccd1 _09292_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_61_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09500__A _10824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17429__A _17429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput130 _12668_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[29] sky130_fd_sc_hd__buf_2
XFILLER_133_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput141 _11661_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wr_en sky130_fd_sc_hd__buf_2
XFILLER_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput152 _12318_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[19] sky130_fd_sc_hd__buf_2
Xoutput163 _12567_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[29] sky130_fd_sc_hd__buf_2
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11713__A1 _11302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_68_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14788__A _14810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13692__A _15260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09765__S0 _09763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09628_ _10899_/A vssd1 vssd1 vccd1 vccd1 _11046_/A sky130_fd_sc_hd__buf_2
XFILLER_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09559_ _10296_/A vssd1 vssd1 vccd1 vccd1 _10523_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14727__S _14735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18157__A1 _19970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16508__A _16528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13631__S _13631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11940__A _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ _17538_/A vssd1 vssd1 vccd1 vccd1 _17542_/A sky130_fd_sc_hd__buf_2
XFILLER_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12441__A2 _12436_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11521_ _11538_/B _11584_/B vssd1 vssd1 vccd1 vccd1 _11521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11452_ _11452_/A _11452_/B vssd1 vssd1 vccd1 vccd1 _11452_/Y sky130_fd_sc_hd__nand2_1
X_14240_ _13771_/X _18737_/Q _14246_/S vssd1 vssd1 vccd1 vccd1 _14241_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10403_ _10403_/A _10403_/B vssd1 vssd1 vccd1 vccd1 _10403_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11401__B1 _10000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14171_ _14171_/A vssd1 vssd1 vccd1 vccd1 _18706_/D sky130_fd_sc_hd__clkbuf_1
X_11383_ _11383_/A _11383_/B vssd1 vssd1 vccd1 vccd1 _11383_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17339__A _17339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10334_ _18815_/Q _19150_/Q _10439_/S vssd1 vssd1 vccd1 vccd1 _10335_/B sky130_fd_sc_hd__mux2_1
XFILLER_125_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input61_A io_ibus_inst[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ _19616_/Q _12891_/X _13121_/X vssd1 vssd1 vccd1 vccd1 _13122_/X sky130_fd_sc_hd__o21a_1
XFILLER_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11387__A _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _19927_/Q vssd1 vssd1 vccd1 vccd1 _16206_/A sky130_fd_sc_hd__buf_2
X_17930_ _17800_/X _17803_/X _17930_/S vssd1 vssd1 vccd1 vccd1 _17930_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10291__A _10312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10265_ _10591_/S vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_140_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12004_ _19586_/Q vssd1 vssd1 vccd1 vccd1 _12027_/A sky130_fd_sc_hd__buf_2
XFILLER_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17861_ _17861_/A vssd1 vssd1 vccd1 vccd1 _17861_/X sky130_fd_sc_hd__buf_2
X_10196_ _10196_/A _10196_/B vssd1 vssd1 vccd1 vccd1 _10196_/X sky130_fd_sc_hd__and2_1
XFILLER_79_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15293__S hold9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output148_A _12220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16812_ _16812_/A _16812_/B vssd1 vssd1 vccd1 vccd1 _16814_/A sky130_fd_sc_hd__nor2_1
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19600_ _19987_/CLK _19600_/D vssd1 vssd1 vccd1 vccd1 _19600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17792_ _17792_/A _17792_/B vssd1 vssd1 vccd1 vccd1 _17792_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13457__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19531_ _19956_/CLK _19531_/D vssd1 vssd1 vccd1 vccd1 _19531_/Q sky130_fd_sc_hd__dfxtp_2
X_16743_ _19684_/Q _16738_/C _16742_/Y vssd1 vssd1 vccd1 vccd1 _19684_/D sky130_fd_sc_hd__o21a_1
X_13955_ _18614_/Q _13660_/X _13961_/S vssd1 vssd1 vccd1 vccd1 _13956_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19462_ _19556_/CLK _19462_/D vssd1 vssd1 vccd1 vccd1 _19462_/Q sky130_fd_sc_hd__dfxtp_1
X_12906_ _19772_/Q _14752_/B _12885_/X _12905_/Y vssd1 vssd1 vccd1 vccd1 _12906_/X
+ sky130_fd_sc_hd__o22a_1
X_16674_ _16674_/A _16680_/C vssd1 vssd1 vccd1 vccd1 _16674_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12011__A _17176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13886_ _13886_/A vssd1 vssd1 vccd1 vccd1 _18583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18413_ _18413_/A vssd1 vssd1 vccd1 vccd1 _18413_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15625_ _14624_/X _19305_/Q _15633_/S vssd1 vssd1 vccd1 vccd1 _15626_/A sky130_fd_sc_hd__mux2_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12837_/A _12837_/B vssd1 vssd1 vccd1 vccd1 _12911_/A sky130_fd_sc_hd__or2_1
X_19393_ _19395_/CLK _19393_/D vssd1 vssd1 vccd1 vccd1 _19393_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12946__A _12951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18148__A1 _19966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10118__S1 _10014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18109__S _18109_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13541__S _13558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12968__B1 _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18344_ _16808_/D _18302_/B _18343_/X _18341_/X vssd1 vssd1 vccd1 vccd1 _20017_/D
+ sky130_fd_sc_hd__o211a_1
X_15556_ _15556_/A vssd1 vssd1 vccd1 vccd1 _19274_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _15783_/A _18454_/Q vssd1 vssd1 vccd1 vccd1 _12768_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12665__B _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14507_ _13755_/X _18833_/Q _14513_/S vssd1 vssd1 vccd1 vccd1 _14508_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18275_ _18275_/A vssd1 vssd1 vccd1 vccd1 _19990_/D sky130_fd_sc_hd__clkbuf_1
X_11719_ _20047_/Q vssd1 vssd1 vccd1 vccd1 _12475_/A sky130_fd_sc_hd__clkbuf_4
X_15487_ _19244_/Q _15257_/X _15489_/S vssd1 vssd1 vccd1 vccd1 _15488_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12699_ _12699_/A vssd1 vssd1 vccd1 vccd1 _12755_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17226_ _19842_/Q _17226_/B vssd1 vssd1 vccd1 vccd1 _17226_/X sky130_fd_sc_hd__or2_1
Xinput10 io_dbus_rdata[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_4
X_14438_ _18815_/Q _14436_/X _14450_/S vssd1 vssd1 vccd1 vccd1 _14439_/A sky130_fd_sc_hd__mux2_1
Xinput21 io_dbus_rdata[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput32 io_dbus_rdata[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_2
Xinput43 io_ibus_inst[18] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput54 io_ibus_inst[28] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13777__A _14602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17157_ _13591_/B _17153_/X _17156_/X _17142_/X vssd1 vssd1 vccd1 vccd1 _19819_/D
+ sky130_fd_sc_hd__o211a_1
Xinput65 io_ibus_inst[9] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
X_14369_ _14574_/A vssd1 vssd1 vccd1 vccd1 _14369_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16108_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16117_/S sky130_fd_sc_hd__buf_2
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17088_ _17087_/B _17087_/C _19791_/Q vssd1 vssd1 vccd1 vccd1 _17089_/C sky130_fd_sc_hd__a21oi_1
XFILLER_170_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16039_ _13393_/X _19441_/Q _16045_/S vssd1 vssd1 vccd1 vccd1 _16040_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15992__A _16060_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__C1 _09736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14401__A _14605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19729_ _19734_/CLK _19729_/D vssd1 vssd1 vccd1 vccd1 _19729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10357__S1 _10326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09413_ _09336_/Y _12678_/A _11952_/D _09403_/X _09412_/X vssd1 vssd1 vccd1 vccd1
+ _13748_/B sky130_fd_sc_hd__o2111a_4
XFILLER_80_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15232__A _15299_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09344_ _19894_/Q _09341_/X _09220_/X _09343_/Y vssd1 vssd1 vccd1 vccd1 _11839_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10434__A1 _09615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09230__A _11601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10434__B2 _19911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09275_ _09425_/B _09275_/B _09275_/C _09275_/D vssd1 vssd1 vccd1 vccd1 _09275_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15378__S _15384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14282__S _14290_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16063__A _16119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11934__B2 _17421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10050_ _11395_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _10050_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09986__S0 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10348__S1 _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13740_ _18537_/Q _13739_/X _13744_/S vssd1 vssd1 vccd1 vccd1 _13741_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10952_ _19363_/Q _18977_/Q _19427_/Q _18546_/Q _09530_/A _09512_/A vssd1 vssd1 vccd1
+ vccd1 _10953_/B sky130_fd_sc_hd__mux4_1
XFILLER_113_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16928__A2 _16955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13671_ _15244_/A vssd1 vssd1 vccd1 vccd1 _14621_/A sky130_fd_sc_hd__buf_2
XANTENNA__14457__S _14466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12766__A _13578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ _11250_/A _10883_/B vssd1 vssd1 vccd1 vccd1 _10883_/X sky130_fd_sc_hd__or2_1
XFILLER_44_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15410_ _15410_/A vssd1 vssd1 vccd1 vccd1 _19209_/D sky130_fd_sc_hd__clkbuf_1
X_12622_ _19609_/Q _12622_/B vssd1 vssd1 vccd1 vccd1 _12622_/X sky130_fd_sc_hd__xor2_1
X_16390_ _16390_/A vssd1 vssd1 vccd1 vccd1 _19553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15341_ _19179_/Q _15254_/X _15345_/S vssd1 vssd1 vccd1 vccd1 _15342_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12553_ _12553_/A vssd1 vssd1 vccd1 vccd1 _18097_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_157_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18060_ _17612_/X _18057_/X _18059_/Y _17705_/A vssd1 vssd1 vccd1 vccd1 _18060_/X
+ sky130_fd_sc_hd__o211a_1
X_11504_ _10043_/X _11497_/X _11499_/Y _11503_/Y _09737_/A vssd1 vssd1 vccd1 vccd1
+ _11504_/X sky130_fd_sc_hd__o311a_1
XFILLER_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15272_ _15272_/A vssd1 vssd1 vccd1 vccd1 _19152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12484_ _12521_/A _12521_/B _12521_/C _12483_/Y vssd1 vssd1 vccd1 vccd1 _12485_/B
+ sky130_fd_sc_hd__a31o_2
X_17011_ _17016_/C _17013_/C _17010_/Y vssd1 vssd1 vccd1 vccd1 _19760_/D sky130_fd_sc_hd__o21a_1
X_14223_ _14223_/A vssd1 vssd1 vccd1 vccd1 _18730_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14192__S _14196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11435_ _10632_/A _11432_/X _11434_/X _10621_/X vssd1 vssd1 vccd1 vccd1 _11435_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11925__B2 _12475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10284__S0 _09926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11366_ _11440_/A _11366_/B vssd1 vssd1 vccd1 vccd1 _11366_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14154_ _14222_/S vssd1 vssd1 vccd1 vccd1 _14163_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_99_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10317_ _10380_/A _10317_/B vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__or2_1
X_13105_ _19647_/Q _12752_/X _12753_/X _19779_/Q _13104_/X vssd1 vssd1 vccd1 vccd1
+ _15686_/B sky130_fd_sc_hd__a221o_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18962_ _19063_/CLK _18962_/D vssd1 vssd1 vccd1 vccd1 _18962_/Q sky130_fd_sc_hd__dfxtp_1
X_11297_ _11170_/A _11296_/X _10980_/A vssd1 vssd1 vccd1 vccd1 _11297_/Y sky130_fd_sc_hd__o21ai_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14920__S _14928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14085_ _18670_/Q _13626_/X _14087_/S vssd1 vssd1 vccd1 vccd1 _14086_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10248_ _18784_/Q _19055_/Q _19279_/Q _19023_/Q _09904_/S _10151_/A vssd1 vssd1 vccd1
+ vccd1 _10248_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _13174_/A vssd1 vssd1 vccd1 vccd1 _13036_/X sky130_fd_sc_hd__clkbuf_2
X_17913_ _17918_/B _17914_/B vssd1 vssd1 vccd1 vccd1 _17917_/B sky130_fd_sc_hd__and2b_1
X_18893_ _19481_/CLK _18893_/D vssd1 vssd1 vccd1 vccd1 _18893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12350__B2 _12349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17844_ _17966_/B vssd1 vssd1 vccd1 vccd1 _17844_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10179_ _18594_/Q _18855_/Q _18754_/Q _19089_/Q _09653_/A _09929_/X vssd1 vssd1 vccd1
+ vccd1 _10179_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17775_ _17765_/X _17767_/Y _17774_/X _17619_/A vssd1 vssd1 vccd1 vccd1 _17775_/X
+ sky130_fd_sc_hd__a211o_1
X_14987_ _19033_/Q _14471_/X _14987_/S vssd1 vssd1 vccd1 vccd1 _14988_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17977__A_N _17973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16726_ _16727_/B _16727_/C _19680_/Q vssd1 vssd1 vccd1 vccd1 _16728_/B sky130_fd_sc_hd__a21oi_1
X_19514_ _19514_/CLK _19514_/D vssd1 vssd1 vccd1 vccd1 _19514_/Q sky130_fd_sc_hd__dfxtp_1
X_13938_ _13938_/A vssd1 vssd1 vccd1 vccd1 _18606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19445_ _19571_/CLK _19445_/D vssd1 vssd1 vccd1 vccd1 _19445_/Q sky130_fd_sc_hd__dfxtp_1
X_16657_ _16674_/A _16661_/C vssd1 vssd1 vccd1 vccd1 _16657_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13869_ _13926_/S vssd1 vssd1 vccd1 vccd1 _13878_/S sky130_fd_sc_hd__buf_2
XANTENNA__14367__S _14367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15608_ _15608_/A vssd1 vssd1 vccd1 vccd1 _19297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19376_ _19566_/CLK _19376_/D vssd1 vssd1 vccd1 vccd1 _19376_/Q sky130_fd_sc_hd__dfxtp_1
X_16588_ _19636_/Q _16590_/C _16587_/Y vssd1 vssd1 vccd1 vccd1 _19636_/D sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_16_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18327_ _17339_/A _18291_/X _18326_/Y _18317_/X vssd1 vssd1 vccd1 vccd1 _20010_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15539_ _19267_/Q _15228_/X _15539_/S vssd1 vssd1 vccd1 vccd1 _15540_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14891__A _14902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__A _10196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18363__A _18380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _19983_/Q _19604_/Q _18264_/S vssd1 vssd1 vccd1 vccd1 _18259_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ _17209_/A vssd1 vssd1 vccd1 vccd1 _17209_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18189_ _18189_/A vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__clkbuf_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ _09957_/X _09958_/X _11475_/A vssd1 vssd1 vccd1 vccd1 _09962_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16611__A _16629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ _09883_/Y _09886_/Y _09889_/Y _09892_/Y _09719_/X vssd1 vssd1 vccd1 vccd1
+ _09893_/X sky130_fd_sc_hd__o221a_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09742__C1 _09741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14277__S _14279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09327_ _13578_/A vssd1 vssd1 vccd1 vccd1 _09339_/A sky130_fd_sc_hd__inv_2
XANTENNA__17588__S _17601_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09258_ _09275_/B vssd1 vssd1 vccd1 vccd1 _09426_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09189_ _20024_/Q _20023_/Q _20022_/Q _20021_/Q vssd1 vssd1 vccd1 vccd1 _09196_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_135_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11220_ _19101_/Q _18867_/Q _19549_/Q _19197_/Q _11083_/S _11164_/X vssd1 vssd1 vccd1
+ vccd1 _11221_/B sky130_fd_sc_hd__mux4_1
XFILLER_88_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11649__B _12670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11151_ _11342_/A _11145_/X _11148_/X _11150_/Y vssd1 vssd1 vccd1 vccd1 _11151_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14740__S _14746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10102_ _09979_/X _10094_/X _10096_/X _10101_/X _09602_/A vssd1 vssd1 vccd1 vccd1
+ _10102_/X sky130_fd_sc_hd__a311o_2
XFILLER_122_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _09610_/A _11071_/X _11081_/X _09618_/A _19898_/Q vssd1 vssd1 vccd1 vccd1
+ _11082_/X sky130_fd_sc_hd__a32o_4
XFILLER_68_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11135__A2 _11123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14910_ _14910_/A vssd1 vssd1 vccd1 vccd1 _18998_/D sky130_fd_sc_hd__clkbuf_1
X_10033_ _10792_/A vssd1 vssd1 vccd1 vccd1 _10757_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__14679__C _18295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11665__A _19323_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15890_ _13357_/X _19375_/Q _15890_/S vssd1 vssd1 vccd1 vccd1 _15891_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input24_A io_dbus_rdata[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ input44/X vssd1 vssd1 vccd1 vccd1 _14841_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13880__A _13926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15821__A2 _13483_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17560_ _17560_/A vssd1 vssd1 vccd1 vccd1 _17560_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14772_ _14772_/A vssd1 vssd1 vccd1 vccd1 _18940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11984_ _12034_/C _11984_/B vssd1 vssd1 vccd1 vccd1 _11984_/Y sky130_fd_sc_hd__nor2_1
X_16511_ _19611_/Q _19610_/Q _19673_/Q _16511_/D vssd1 vssd1 vccd1 vccd1 _16520_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__18220__A0 _19966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13723_ _14660_/A vssd1 vssd1 vccd1 vccd1 _13723_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17491_ _17486_/X _17490_/X _17601_/S vssd1 vssd1 vccd1 vccd1 _17491_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10935_ _11355_/A _12643_/A vssd1 vssd1 vccd1 vccd1 _11579_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12496__A _18340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19230_ _19392_/CLK _19230_/D vssd1 vssd1 vccd1 vccd1 _19230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16442_ _16442_/A vssd1 vssd1 vccd1 vccd1 _19577_/D sky130_fd_sc_hd__clkbuf_1
X_13654_ _15231_/A vssd1 vssd1 vccd1 vccd1 _14608_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10866_ _19902_/Q vssd1 vssd1 vccd1 vccd1 _10866_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19161_ _19906_/CLK _19161_/D vssd1 vssd1 vccd1 vccd1 _19161_/Q sky130_fd_sc_hd__dfxtp_1
X_12605_ _17323_/A _18286_/A _18283_/A _12606_/D vssd1 vssd1 vccd1 vccd1 _12605_/X
+ sky130_fd_sc_hd__or4_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _16441_/S vssd1 vssd1 vccd1 vccd1 _16382_/S sky130_fd_sc_hd__clkbuf_4
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14915__S _14915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13585_ _13584_/X _18503_/Q _13598_/S vssd1 vssd1 vccd1 vccd1 _13586_/A sky130_fd_sc_hd__mux2_1
X_10797_ _09693_/A _10790_/Y _10792_/Y _10794_/Y _10796_/Y vssd1 vssd1 vccd1 vccd1
+ _10797_/X sky130_fd_sc_hd__o32a_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _18121_/B _18108_/Y _18111_/Y vssd1 vssd1 vccd1 vccd1 _18112_/Y sky130_fd_sc_hd__a21oi_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11071__A1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15324_ _15324_/A vssd1 vssd1 vccd1 vccd1 _19171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19092_ _19092_/CLK _19092_/D vssd1 vssd1 vccd1 vccd1 _19092_/Q sky130_fd_sc_hd__dfxtp_1
X_12536_ _12536_/A vssd1 vssd1 vccd1 vccd1 _12538_/B sky130_fd_sc_hd__inv_8
XFILLER_40_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18043_ _18046_/A _18046_/B vssd1 vssd1 vccd1 vccd1 _18043_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15255_ _19147_/Q _15254_/X _15261_/S vssd1 vssd1 vccd1 vccd1 _15256_/A sky130_fd_sc_hd__mux2_1
X_12467_ _12463_/Y _12466_/Y _12562_/S vssd1 vssd1 vccd1 vccd1 _12467_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output92_A _12559_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ _14206_/A vssd1 vssd1 vccd1 vccd1 _18722_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10257__S0 _09904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11418_ _11418_/A _12659_/B vssd1 vssd1 vccd1 vccd1 _11554_/B sky130_fd_sc_hd__nand2_1
X_15186_ _15186_/A vssd1 vssd1 vccd1 vccd1 _19124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12398_ _19839_/Q _12419_/C vssd1 vssd1 vccd1 vccd1 _12398_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12571__A1 _17542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ _14137_/A vssd1 vssd1 vccd1 vccd1 _18693_/D sky130_fd_sc_hd__clkbuf_1
X_11349_ _11302_/Y _11582_/D _11348_/Y vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__a21o_1
X_19994_ _20027_/CLK _19994_/D vssd1 vssd1 vccd1 vccd1 _19994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18945_ _19557_/CLK _18945_/D vssd1 vssd1 vccd1 vccd1 _18945_/Q sky130_fd_sc_hd__dfxtp_1
X_14068_ _18664_/Q _13735_/X _14068_/S vssd1 vssd1 vccd1 vccd1 _14069_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13520__A0 _19922_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ _13558_/S vssd1 vssd1 vccd1 vccd1 _13090_/S sky130_fd_sc_hd__buf_2
XFILLER_100_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18876_ _19302_/CLK _18876_/D vssd1 vssd1 vccd1 vccd1 _18876_/Q sky130_fd_sc_hd__dfxtp_1
X_17827_ _17827_/A vssd1 vssd1 vccd1 vccd1 _17971_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13790__A _14615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15481__S _15489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15812__A2 _13467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17758_ _18019_/A vssd1 vssd1 vccd1 vccd1 _17758_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16709_ _16728_/A _16709_/B _16709_/C vssd1 vssd1 vccd1 vccd1 _19674_/D sky130_fd_sc_hd__nor3_1
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17689_ _17684_/X _17687_/X _17930_/S vssd1 vssd1 vccd1 vccd1 _17689_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19428_ _19552_/CLK _19428_/D vssd1 vssd1 vccd1 vccd1 _19428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09211__C _11601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19359_ _19455_/CLK _19359_/D vssd1 vssd1 vccd1 vccd1 _19359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10248__S0 _09904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_144_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14560__S _14568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09945_ _09750_/A _09934_/X _09943_/X _09757_/A _09944_/Y vssd1 vssd1 vccd1 vccd1
+ _12662_/B sky130_fd_sc_hd__o32a_4
X_09876_ _09924_/S vssd1 vssd1 vccd1 vccd1 _10173_/S sky130_fd_sc_hd__buf_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10420__S0 _10465_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10876__B2 _11014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__C1 _10621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11932__B _11969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10720_ _10768_/A _10720_/B vssd1 vssd1 vccd1 vccd1 _10720_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_191_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _11448_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _10651_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14735__S _14735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11053__A1 _10961_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10487__S0 _10390_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ _18650_/Q _19241_/Q _19403_/Q _18618_/Q _10494_/S _10332_/A vssd1 vssd1 vccd1
+ vccd1 _10583_/B sky130_fd_sc_hd__mux4_1
XFILLER_22_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13370_ _19662_/Q _12887_/X _12889_/X _19794_/Q _13369_/X vssd1 vssd1 vccd1 vccd1
+ _13370_/X sky130_fd_sc_hd__a221o_4
XFILLER_167_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10261__C1 _09605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12321_ _12376_/A _12657_/B _12377_/A _12320_/X vssd1 vssd1 vccd1 vccd1 _12322_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15040_ _19056_/Q _14443_/X _15044_/S vssd1 vssd1 vccd1 vccd1 _15041_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12252_ _12252_/A vssd1 vssd1 vccd1 vccd1 _17389_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11203_ _19486_/Q _18898_/Q _18935_/Q _18509_/Q _11306_/S _09511_/A vssd1 vssd1 vccd1
+ vccd1 _11204_/B sky130_fd_sc_hd__mux4_1
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12183_ _19831_/Q vssd1 vssd1 vccd1 vccd1 _17192_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11134_ _10875_/X _11125_/X _11127_/X _11133_/X _09600_/A vssd1 vssd1 vccd1 vccd1
+ _11134_/X sky130_fd_sc_hd__a311o_2
X_16991_ _16994_/C _16992_/C _19755_/Q vssd1 vssd1 vccd1 vccd1 _16993_/B sky130_fd_sc_hd__a21oi_1
XFILLER_150_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15942_ _15988_/S vssd1 vssd1 vccd1 vccd1 _15951_/S sky130_fd_sc_hd__clkbuf_4
X_18730_ _19482_/CLK _18730_/D vssd1 vssd1 vccd1 vccd1 _18730_/Q sky130_fd_sc_hd__dfxtp_1
X_11065_ _11065_/A vssd1 vssd1 vccd1 vccd1 _11065_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11513__C1 _10063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17244__A1 _13603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ _10977_/A vssd1 vssd1 vccd1 vccd1 _10017_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18661_ _19510_/CLK _18661_/D vssd1 vssd1 vccd1 vccd1 _18661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15873_ _13230_/X _19367_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15874_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16452__C1 _18412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17612_ _17785_/A vssd1 vssd1 vccd1 vccd1 _17612_/X sky130_fd_sc_hd__clkbuf_2
X_14824_ _14824_/A vssd1 vssd1 vccd1 vccd1 _18964_/D sky130_fd_sc_hd__clkbuf_1
X_18592_ _19311_/CLK _18592_/D vssd1 vssd1 vccd1 vccd1 _18592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17543_ _17785_/A vssd1 vssd1 vccd1 vccd1 _17543_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14755_ _14823_/S vssd1 vssd1 vccd1 vccd1 _14764_/S sky130_fd_sc_hd__buf_2
XFILLER_44_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11967_ _19964_/Q _10961_/X _12077_/S vssd1 vssd1 vccd1 vccd1 _17412_/A sky130_fd_sc_hd__mux2_4
XANTENNA__10714__S1 _10665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ _14647_/A vssd1 vssd1 vccd1 vccd1 _13706_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17474_ _12385_/A _17832_/B _17504_/S vssd1 vssd1 vccd1 vccd1 _17474_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_1_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _20049_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09312__B _14501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10918_ _18771_/Q _19042_/Q _19266_/Q _19010_/Q _10914_/X _10969_/A vssd1 vssd1 vccd1
+ vccd1 _10918_/X sky130_fd_sc_hd__mux4_1
X_14686_ _14686_/A vssd1 vssd1 vccd1 vccd1 _18897_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10458__B _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11898_ _11712_/C _11849_/D _17739_/S _11898_/D vssd1 vssd1 vccd1 vccd1 _11898_/X
+ sky130_fd_sc_hd__and4bb_2
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19213_ _19311_/CLK _19213_/D vssd1 vssd1 vccd1 vccd1 _19213_/Q sky130_fd_sc_hd__dfxtp_1
X_16425_ _16425_/A vssd1 vssd1 vccd1 vccd1 _19569_/D sky130_fd_sc_hd__clkbuf_1
X_13637_ _13637_/A vssd1 vssd1 vccd1 vccd1 _18512_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14645__S _14654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10849_ _18804_/Q _19139_/Q _10849_/S vssd1 vssd1 vccd1 vccd1 _10850_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12954__A _12976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19144_ _19272_/CLK _19144_/D vssd1 vssd1 vccd1 vccd1 _19144_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11044__A1 _11216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16356_ _19542_/Q _16300_/A _16354_/Y _16355_/X vssd1 vssd1 vccd1 vccd1 _19542_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13568_ _13580_/A vssd1 vssd1 vccd1 vccd1 _13568_/X sky130_fd_sc_hd__buf_2
XFILLER_158_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15307_ _15307_/A vssd1 vssd1 vccd1 vccd1 _19163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12519_ _19605_/Q _12363_/X _12514_/X _12518_/X vssd1 vssd1 vccd1 vccd1 _12519_/X
+ sky130_fd_sc_hd__o22a_4
X_19075_ _19203_/CLK _19075_/D vssd1 vssd1 vccd1 vccd1 _19075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16287_ _19529_/Q _16285_/X _16325_/S vssd1 vssd1 vccd1 vccd1 _16288_/A sky130_fd_sc_hd__mux2_1
X_13499_ _19766_/Q _12840_/X _13498_/X _12846_/X vssd1 vssd1 vccd1 vccd1 _13499_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18026_ _17781_/X _17839_/B _18025_/X _17940_/X vssd1 vssd1 vccd1 vccd1 _18026_/X
+ sky130_fd_sc_hd__a211o_1
X_15238_ _15238_/A vssd1 vssd1 vccd1 vccd1 _15238_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15730__A1 _12854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15476__S _15478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15169_ _19116_/Q vssd1 vssd1 vccd1 vccd1 _15170_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_113_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14380__S _14386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10650__S0 _10649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19977_ _19986_/CLK _19977_/D vssd1 vssd1 vccd1 vccd1 _19977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09730_ _10176_/A vssd1 vssd1 vccd1 vccd1 _09730_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18928_ _20000_/CLK _18928_/D vssd1 vssd1 vccd1 vccd1 _18928_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11504__C1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10402__S0 _10268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09661_ _10105_/A vssd1 vssd1 vccd1 vccd1 _09662_/A sky130_fd_sc_hd__buf_4
X_18859_ _19317_/CLK _18859_/D vssd1 vssd1 vccd1 vccd1 _18859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13724__S _13736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16100__S _16106_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ _19515_/Q _18927_/Q _18964_/Q _18538_/Q _09568_/X _09762_/A vssd1 vssd1 vccd1
+ vccd1 _09592_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09503__A _10560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10649__A _10700_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09571__S1 _09569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14555__S _14557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10469__S0 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11130__S1 _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17710__A2 _17558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14290__S _14290_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17167__A _17197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17474__A1 _17832_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_138_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09928_ _09874_/X _09925_/Y _09927_/Y _10279_/A vssd1 vssd1 vccd1 vccd1 _09928_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20048_ _20048_/CLK _20048_/D vssd1 vssd1 vccd1 vccd1 _20048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09859_ _19123_/Q _18889_/Q _19571_/Q _19219_/Q _10175_/S _09858_/X vssd1 vssd1 vccd1
+ vccd1 _09860_/B sky130_fd_sc_hd__mux4_2
XFILLER_86_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10944__S1 _10943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12870_ _19718_/Q _12775_/X _12777_/X _19686_/Q _12869_/X vssd1 vssd1 vccd1 vccd1
+ _12870_/X sky130_fd_sc_hd__a221o_2
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11821_ _12029_/C vssd1 vssd1 vccd1 vccd1 _11870_/C sky130_fd_sc_hd__clkbuf_2
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _13803_/X _18848_/Q _14546_/S vssd1 vssd1 vccd1 vccd1 _14541_/A sky130_fd_sc_hd__mux2_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11381__A1_N _11369_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _17467_/A _11712_/C _11688_/A vssd1 vssd1 vccd1 vccd1 _11759_/A sky130_fd_sc_hd__o21ai_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10703_/A _10703_/B vssd1 vssd1 vccd1 vccd1 _10703_/Y sky130_fd_sc_hd__nand2_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14675_/A vssd1 vssd1 vccd1 vccd1 _14471_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12774__A _15700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11683_ _12600_/A _11681_/Y _17394_/C vssd1 vssd1 vccd1 vccd1 _17381_/C sky130_fd_sc_hd__o21a_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16299_/A vssd1 vssd1 vccd1 vccd1 _16223_/S sky130_fd_sc_hd__clkbuf_2
X_13422_ _13418_/X _13420_/Y _13421_/Y vssd1 vssd1 vccd1 vccd1 _15273_/A sky130_fd_sc_hd__a21oi_4
XFILLER_174_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10634_ _10574_/A _10633_/X _09577_/A vssd1 vssd1 vccd1 vccd1 _10634_/X sky130_fd_sc_hd__o21a_1
X_17190_ _15738_/X _17182_/X _17189_/X _17185_/X vssd1 vssd1 vccd1 vccd1 _19830_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _19486_/Q _14583_/A _16145_/S vssd1 vssd1 vccd1 vccd1 _16142_/A sky130_fd_sc_hd__mux2_1
X_13353_ _13353_/A vssd1 vssd1 vccd1 vccd1 _13353_/X sky130_fd_sc_hd__clkbuf_2
X_10565_ _10574_/A _10565_/B vssd1 vssd1 vccd1 vccd1 _10565_/X sky130_fd_sc_hd__or2_1
XANTENNA__10294__A _10294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12304_ _12332_/A _12331_/A vssd1 vssd1 vccd1 vccd1 _12306_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16072_ _16072_/A vssd1 vssd1 vccd1 vccd1 _19455_/D sky130_fd_sc_hd__clkbuf_1
X_13284_ _19865_/Q _12842_/A _13343_/A _19832_/Q vssd1 vssd1 vccd1 vccd1 _13284_/X
+ sky130_fd_sc_hd__a22o_1
X_10496_ _18812_/Q _19147_/Q _10496_/S vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__mux2_1
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15023_ _15023_/A vssd1 vssd1 vccd1 vccd1 _19048_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15296__S _15299_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19900_ _19997_/CLK _19900_/D vssd1 vssd1 vccd1 vccd1 _19900_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_108_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12235_ _19586_/Q hold21/A _19590_/Q _19593_/Q vssd1 vssd1 vccd1 vccd1 _12237_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_108_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19831_ _19831_/CLK _19831_/D vssd1 vssd1 vccd1 vccd1 _19831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12166_ _12198_/S vssd1 vssd1 vccd1 vccd1 _12303_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_96_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10741__B _10741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ _11271_/A vssd1 vssd1 vccd1 vccd1 _11117_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19762_ _19762_/CLK _19762_/D vssd1 vssd1 vccd1 vccd1 _19762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16974_ _17073_/A vssd1 vssd1 vccd1 vccd1 _17007_/A sky130_fd_sc_hd__clkbuf_2
X_12097_ _12097_/A vssd1 vssd1 vccd1 vccd1 _12188_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18713_ _19575_/CLK _18713_/D vssd1 vssd1 vccd1 vccd1 _18713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15925_ _19390_/Q _15206_/X _15929_/S vssd1 vssd1 vccd1 vccd1 _15926_/A sky130_fd_sc_hd__mux2_1
X_11048_ _11216_/A _11047_/X _10920_/X vssd1 vssd1 vccd1 vccd1 _11048_/Y sky130_fd_sc_hd__o21ai_1
X_19693_ _19726_/CLK _19693_/D vssd1 vssd1 vccd1 vccd1 _19693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 io_dbus_rdata[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15325__A _15371_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15856_ _15856_/A vssd1 vssd1 vccd1 vccd1 _19359_/D sky130_fd_sc_hd__clkbuf_1
X_18644_ _19204_/CLK _18644_/D vssd1 vssd1 vccd1 vccd1 _18644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12668__B _12668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14807_ _14807_/A vssd1 vssd1 vccd1 vccd1 _18956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15787_ _15787_/A vssd1 vssd1 vccd1 vccd1 _19345_/D sky130_fd_sc_hd__clkbuf_1
X_18575_ _19292_/CLK _18575_/D vssd1 vssd1 vccd1 vccd1 _18575_/Q sky130_fd_sc_hd__dfxtp_1
X_12999_ _19642_/Q _12727_/X _12729_/X _19774_/Q _12998_/X vssd1 vssd1 vccd1 vccd1
+ _13569_/B sky130_fd_sc_hd__a221o_1
XFILLER_33_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17540__A _18118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14738_ _18921_/Q _14452_/X _14746_/S vssd1 vssd1 vccd1 vccd1 _14739_/A sky130_fd_sc_hd__mux2_1
X_17526_ _17603_/A vssd1 vssd1 vccd1 vccd1 _17527_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17457_ _17457_/A vssd1 vssd1 vccd1 vccd1 _17820_/B sky130_fd_sc_hd__clkbuf_2
X_14669_ _14669_/A vssd1 vssd1 vccd1 vccd1 _14669_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16408_ _16408_/A vssd1 vssd1 vccd1 vccd1 _19561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15951__A1 _15244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17388_ _18118_/B _17668_/A vssd1 vssd1 vccd1 vccd1 _17388_/X sky130_fd_sc_hd__or2_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_164_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19789_/CLK sky130_fd_sc_hd__clkbuf_16
X_19127_ _19575_/CLK _19127_/D vssd1 vssd1 vccd1 vccd1 _19127_/Q sky130_fd_sc_hd__dfxtp_1
X_16339_ _16347_/C _16338_/Y _12444_/X vssd1 vssd1 vccd1 vccd1 _16340_/B sky130_fd_sc_hd__a21oi_2
XFILLER_134_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19058_ _19058_/CLK _19058_/D vssd1 vssd1 vccd1 vccd1 _19058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18009_ _18009_/A vssd1 vssd1 vccd1 vccd1 _18088_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_142_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_179_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19876_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17208__A1 _15770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ _09722_/A _09700_/X _09712_/X vssd1 vssd1 vccd1 vccd1 _09713_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_102_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19493_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15235__A _15235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09644_ _10909_/S vssd1 vssd1 vccd1 vccd1 _11495_/S sky130_fd_sc_hd__buf_2
XFILLER_67_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09575_ _09975_/A vssd1 vssd1 vccd1 vccd1 _10621_/A sky130_fd_sc_hd__buf_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12569__A2_N _12669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_117_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19552_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12594__A _12606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17144__B1 _17101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11003__A _11003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10350_ _11464_/A vssd1 vssd1 vccd1 vccd1 _10583_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10281_ _09884_/A _10280_/X _09696_/A vssd1 vssd1 vccd1 vccd1 _10281_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12020_ _12020_/A _17459_/A vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__or2_1
XANTENNA__13181__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13971_ _13971_/A vssd1 vssd1 vccd1 vccd1 _18621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12769__A _12853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13484__A2 _10134_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15710_ _15783_/A _18445_/Q vssd1 vssd1 vccd1 vccd1 _15710_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11673__A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12922_ _15702_/A _18461_/Q vssd1 vssd1 vccd1 vccd1 _12922_/Y sky130_fd_sc_hd__nand2_1
X_16690_ _16689_/B _16689_/C _19671_/Q vssd1 vssd1 vccd1 vccd1 _16691_/C sky130_fd_sc_hd__a21oi_1
XFILLER_20_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15641_ _15641_/A vssd1 vssd1 vccd1 vccd1 _19312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12853_ _12853_/A vssd1 vssd1 vccd1 vccd1 _12853_/X sky130_fd_sc_hd__buf_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _18401_/A vssd1 vssd1 vccd1 vccd1 _18380_/A sky130_fd_sc_hd__buf_2
XFILLER_33_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11804_ _11704_/X _11802_/X _11803_/X _11616_/A vssd1 vssd1 vccd1 vccd1 _11804_/X
+ sky130_fd_sc_hd__o211a_1
X_15572_ _19282_/Q _15276_/X _15572_/S vssd1 vssd1 vccd1 vccd1 _15573_/A sky130_fd_sc_hd__mux2_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _19756_/Q _12692_/X _12783_/X _12714_/X vssd1 vssd1 vccd1 vccd1 _12784_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _15828_/X _19878_/Q _17313_/S vssd1 vssd1 vccd1 vccd1 _17312_/A sky130_fd_sc_hd__mux2_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10455__C1 _09718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14523_/A vssd1 vssd1 vccd1 vccd1 _18840_/D sky130_fd_sc_hd__clkbuf_1
X_18291_ _18345_/B vssd1 vssd1 vccd1 vccd1 _18291_/X sky130_fd_sc_hd__buf_2
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11699_/B _11734_/X _12097_/A vssd1 vssd1 vccd1 vccd1 _11735_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19560_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _19848_/Q _17242_/B vssd1 vssd1 vccd1 vccd1 _17242_/X sky130_fd_sc_hd__or2_1
XANTENNA__12935__C _12937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14454_ _18820_/Q _14452_/X _14466_/S vssd1 vssd1 vccd1 vccd1 _14455_/A sky130_fd_sc_hd__mux2_1
X_11666_ _12286_/A vssd1 vssd1 vccd1 vccd1 _12562_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_174_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13405_ _19632_/Q _13204_/X _13404_/X vssd1 vssd1 vccd1 vccd1 _13405_/X sky130_fd_sc_hd__o21a_1
X_10617_ _11481_/S vssd1 vssd1 vccd1 vccd1 _10617_/X sky130_fd_sc_hd__buf_4
X_17173_ _19824_/Q _17180_/B vssd1 vssd1 vccd1 vccd1 _17173_/X sky130_fd_sc_hd__or2_1
XFILLER_167_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14385_ _14589_/A vssd1 vssd1 vccd1 vccd1 _14385_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11597_ _09807_/A _11538_/A _11545_/X _11595_/X _11596_/Y vssd1 vssd1 vccd1 vccd1
+ _11597_/X sky130_fd_sc_hd__a2111o_1
X_16124_ _13487_/X _19479_/Q _16128_/S vssd1 vssd1 vccd1 vccd1 _16125_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16489__A2 _12494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ _13363_/A _13336_/B _13362_/B vssd1 vssd1 vccd1 vccd1 _13336_/X sky130_fd_sc_hd__or3_1
XFILLER_155_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10548_ _10548_/A _10548_/B vssd1 vssd1 vccd1 vccd1 _10548_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_96_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19268_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10853__S0 _10048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10773__A3 _10771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16055_ _16055_/A vssd1 vssd1 vccd1 vccd1 _19448_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11970__A2 _17772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13267_ _19624_/Q _12911_/X _13266_/X vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__o21a_1
XFILLER_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10479_ _18652_/Q _19243_/Q _19405_/Q _18620_/Q _10417_/S _09841_/A vssd1 vssd1 vccd1
+ vccd1 _10479_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15006_ _15006_/A vssd1 vssd1 vccd1 vccd1 _19040_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09318__A _20044_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ _12218_/A vssd1 vssd1 vccd1 vccd1 _12218_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13198_ _13255_/A vssd1 vssd1 vccd1 vccd1 _13363_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19814_ _20044_/CLK _19814_/D vssd1 vssd1 vccd1 vccd1 _19814_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_96_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12149_ _19591_/Q vssd1 vssd1 vccd1 vccd1 _12152_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19745_ _19745_/CLK _19745_/D vssd1 vssd1 vccd1 vccd1 _19745_/Q sky130_fd_sc_hd__dfxtp_1
X_16957_ _19745_/Q _16957_/B _16957_/C vssd1 vssd1 vccd1 vccd1 _16958_/D sky130_fd_sc_hd__and3_1
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15908_ _13487_/X _19383_/Q _15912_/S vssd1 vssd1 vccd1 vccd1 _15909_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_34_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19308_/CLK sky130_fd_sc_hd__clkbuf_16
X_19676_ _19682_/CLK _19676_/D vssd1 vssd1 vccd1 vccd1 _19676_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16949__B1 _16860_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16888_ _19727_/Q _19726_/Q _19725_/Q _16888_/D vssd1 vssd1 vccd1 vccd1 _16896_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18627_ _19412_/CLK _18627_/D vssd1 vssd1 vccd1 vccd1 _18627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15839_ _15818_/X _18467_/Q _15819_/Y _15838_/X vssd1 vssd1 vccd1 vccd1 _15839_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_18_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11238__A1 _11001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _20011_/Q vssd1 vssd1 vccd1 vccd1 _09398_/B sky130_fd_sc_hd__clkbuf_1
X_18558_ _19565_/CLK _18558_/D vssd1 vssd1 vccd1 vccd1 _18558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10446__C1 _09740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__S1 _10006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17509_ _17505_/X _17508_/X _17677_/S vssd1 vssd1 vccd1 vccd1 _17510_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_49_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19058_/CLK sky130_fd_sc_hd__clkbuf_16
X_09291_ _20000_/Q vssd1 vssd1 vccd1 vccd1 _14074_/A sky130_fd_sc_hd__buf_4
XFILLER_162_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18489_ _19566_/CLK _18489_/D vssd1 vssd1 vccd1 vccd1 _18489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13303__A _13353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15929__S _15929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10749__B1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput120 _12632_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[1] sky130_fd_sc_hd__buf_2
Xoutput131 _12633_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[2] sky130_fd_sc_hd__buf_2
Xoutput142 _11671_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_82_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput153 _16447_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[1] sky130_fd_sc_hd__buf_2
XANTENNA__09228__A _11601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput164 _11799_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_82_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10921__B1 _10920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09765__S1 _09526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09627_ _11291_/A vssd1 vssd1 vccd1 vccd1 _10899_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09558_ _10630_/A vssd1 vssd1 vccd1 vccd1 _10296_/A sky130_fd_sc_hd__buf_4
XFILLER_43_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12977__A1 _18462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09489_ _10521_/A vssd1 vssd1 vccd1 vccd1 _10428_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11520_ _11520_/A _12669_/B vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__or2_1
XFILLER_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11451_ _18824_/Q _19159_/Q _11451_/S vssd1 vssd1 vccd1 vccd1 _11452_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11088__S0 _10017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _19375_/Q _18989_/Q _19439_/Q _18558_/Q _10268_/S _10335_/A vssd1 vssd1 vccd1
+ vccd1 _10403_/B sky130_fd_sc_hd__mux4_1
XANTENNA__11401__A1 _11383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10835__S0 _10735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14170_ _13774_/X _18706_/Q _14174_/S vssd1 vssd1 vccd1 vccd1 _14171_/A sky130_fd_sc_hd__mux2_1
X_11382_ _19111_/Q _18877_/Q _19559_/Q _19207_/Q _10053_/X _10054_/X vssd1 vssd1 vccd1
+ vccd1 _11383_/B sky130_fd_sc_hd__mux4_2
XANTENNA__17339__B _18324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ _19744_/Q _12692_/X _13120_/X _12714_/X vssd1 vssd1 vccd1 vccd1 _13121_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_3_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10333_ _10333_/A vssd1 vssd1 vccd1 vccd1 _10335_/A sky130_fd_sc_hd__buf_2
XFILLER_140_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input54_A io_ibus_inst[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _13066_/A vssd1 vssd1 vccd1 vccd1 _13054_/A sky130_fd_sc_hd__buf_2
X_10264_ _10264_/A _10264_/B vssd1 vssd1 vccd1 vccd1 _10264_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12003_ _12003_/A vssd1 vssd1 vccd1 vccd1 _12003_/Y sky130_fd_sc_hd__inv_6
XFILLER_78_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10195_ _18817_/Q _19152_/Q _10195_/S vssd1 vssd1 vccd1 vccd1 _10196_/B sky130_fd_sc_hd__mux2_1
X_17860_ _10775_/Y _12980_/X _17859_/X vssd1 vssd1 vccd1 vccd1 _19903_/D sky130_fd_sc_hd__a21oi_1
XFILLER_121_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16811_ _16811_/A _16816_/D vssd1 vssd1 vccd1 vccd1 _16812_/B sky130_fd_sc_hd__nand2_4
XFILLER_121_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17840__B2 _12024_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17791_ _17791_/A vssd1 vssd1 vccd1 vccd1 _17791_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19530_ _19988_/CLK _19530_/D vssd1 vssd1 vccd1 vccd1 _19530_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10511__S _10560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13954_ _13954_/A vssd1 vssd1 vccd1 vccd1 _18613_/D sky130_fd_sc_hd__clkbuf_1
X_16742_ _16775_/A _16747_/C vssd1 vssd1 vccd1 vccd1 _16742_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12905_ _12829_/X _17220_/A _14752_/B vssd1 vssd1 vccd1 vccd1 _12905_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_47_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16673_ _16673_/A vssd1 vssd1 vccd1 vccd1 _16680_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_19461_ _19555_/CLK _19461_/D vssd1 vssd1 vccd1 vccd1 _19461_/Q sky130_fd_sc_hd__dfxtp_1
X_13885_ _13790_/X _18583_/Q _13889_/S vssd1 vssd1 vccd1 vccd1 _13886_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18412_ _18412_/A _18412_/B vssd1 vssd1 vccd1 vccd1 _20045_/D sky130_fd_sc_hd__nor2_1
XANTENNA__12417__A0 _12414_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15624_ _15646_/A vssd1 vssd1 vccd1 vccd1 _15633_/S sky130_fd_sc_hd__buf_2
X_12836_ _19621_/Q vssd1 vssd1 vccd1 vccd1 _16547_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _19392_/CLK _19392_/D vssd1 vssd1 vccd1 vccd1 _19392_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09601__A _09601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12968__A1 _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15555_ _19274_/Q _15251_/X _15561_/S vssd1 vssd1 vccd1 vccd1 _15556_/A sky130_fd_sc_hd__mux2_1
X_18343_ _18343_/A _18349_/B vssd1 vssd1 vccd1 vccd1 _18343_/X sky130_fd_sc_hd__or2_1
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _15837_/A vssd1 vssd1 vccd1 vccd1 _15783_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14506_ _14506_/A vssd1 vssd1 vccd1 vccd1 _18832_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18274_ _18352_/A _18274_/B vssd1 vssd1 vccd1 vccd1 _18275_/A sky130_fd_sc_hd__or2_1
X_11718_ _11724_/D vssd1 vssd1 vccd1 vccd1 _17378_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15486_ _15486_/A vssd1 vssd1 vccd1 vccd1 _19243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ _12992_/A vssd1 vssd1 vccd1 vccd1 _12699_/A sky130_fd_sc_hd__buf_2
XFILLER_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14437_ _14453_/A vssd1 vssd1 vccd1 vccd1 _14450_/S sky130_fd_sc_hd__buf_2
X_17225_ _17225_/A vssd1 vssd1 vccd1 vccd1 _17225_/Y sky130_fd_sc_hd__inv_2
Xinput11 io_dbus_rdata[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_4
X_11649_ _11901_/A _12670_/A _11692_/C vssd1 vssd1 vccd1 vccd1 _11650_/D sky130_fd_sc_hd__or3_1
Xinput22 io_dbus_rdata[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12962__A _12976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput33 io_dbus_valid vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_8
XANTENNA__09597__B1 _09580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17156_ _19819_/Q _17164_/B vssd1 vssd1 vccd1 vccd1 _17156_/X sky130_fd_sc_hd__or2_1
Xinput44 io_ibus_inst[19] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
Xinput55 io_ibus_inst[29] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_6
X_14368_ _14368_/A vssd1 vssd1 vccd1 vccd1 _18794_/D sky130_fd_sc_hd__clkbuf_1
Xinput66 io_ibus_valid vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_4
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16107_ _16107_/A vssd1 vssd1 vccd1 vccd1 _19471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13319_ input9/X _13318_/X _13306_/X vssd1 vssd1 vccd1 vccd1 _13319_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17087_ _19791_/Q _17087_/B _17087_/C vssd1 vssd1 vccd1 vccd1 _17089_/B sky130_fd_sc_hd__and3_1
X_14299_ _14367_/S vssd1 vssd1 vccd1 vccd1 _14308_/S sky130_fd_sc_hd__buf_2
X_16038_ _16038_/A vssd1 vssd1 vccd1 vccd1 _19440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_12_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11251__S0 _11057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18084__B2 _12509_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17989_ _17985_/B _17989_/B vssd1 vssd1 vccd1 vccd1 _17990_/D sky130_fd_sc_hd__and2b_1
XFILLER_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19728_ _19734_/CLK _19728_/D vssd1 vssd1 vccd1 vccd1 _19728_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13017__B _18295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19659_ _19792_/CLK _19659_/D vssd1 vssd1 vccd1 vccd1 _19659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13732__S _13736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09412_ _09358_/X _12820_/B _09406_/Y _11952_/B vssd1 vssd1 vccd1 vccd1 _09412_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09343_ _19891_/Q _09342_/Y _19892_/Q vssd1 vssd1 vccd1 vccd1 _09343_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09511__A _09511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13081__B1 _13080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13033__A _15203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09230__B _09238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ _09329_/A _17331_/B _11682_/B vssd1 vssd1 vccd1 vccd1 _11608_/A sky130_fd_sc_hd__or3b_1
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15659__S _15659_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13384__B2 _19535_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10198__A1 _10161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11934__A2 _17418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13179__S _13196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14799__A _14810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13907__S _13911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18075__A1 _19919_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17175__A _17175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11242__S0 _11057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09986__S1 _09985_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10370__A1 _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10951_ _11012_/A _10951_/B _10951_/C vssd1 vssd1 vccd1 vccd1 _10951_/X sky130_fd_sc_hd__or3_2
XANTENNA__14738__S _14746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10122__A1 _10846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16519__A _16528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13670_ _13670_/A vssd1 vssd1 vccd1 vccd1 _18520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10882_ _18579_/Q _18840_/Q _18739_/Q _19074_/Q _11305_/S _11236_/A vssd1 vssd1 vccd1
+ vccd1 _10883_/B sky130_fd_sc_hd__mux4_1
XFILLER_32_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12621_ _12620_/A _12620_/B _12395_/S vssd1 vssd1 vccd1 vccd1 _12621_/X sky130_fd_sc_hd__a21o_1
X_15340_ _15340_/A vssd1 vssd1 vccd1 vccd1 _19178_/D sky130_fd_sc_hd__clkbuf_1
X_12552_ _19986_/Q _11470_/A _12573_/S vssd1 vssd1 vccd1 vccd1 _12553_/A sky130_fd_sc_hd__mux2_4
XFILLER_129_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11503_ _11510_/A _11500_/X _11502_/X vssd1 vssd1 vccd1 vccd1 _11503_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15271_ _19152_/Q _15270_/X _15277_/S vssd1 vssd1 vccd1 vccd1 _15272_/A sky130_fd_sc_hd__mux2_1
X_12483_ _12460_/Y _12458_/A _12458_/B vssd1 vssd1 vccd1 vccd1 _12483_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17010_ _17016_/C _17013_/C _16860_/X vssd1 vssd1 vccd1 vccd1 _17010_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14222_ _13850_/X _18730_/Q _14222_/S vssd1 vssd1 vccd1 vccd1 _14223_/A sky130_fd_sc_hd__mux2_1
X_11434_ _11443_/A _11434_/B vssd1 vssd1 vccd1 vccd1 _11434_/X sky130_fd_sc_hd__or2_1
XFILLER_22_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13597__B _13597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14153_ _14209_/A vssd1 vssd1 vccd1 vccd1 _14222_/S sky130_fd_sc_hd__buf_4
X_11365_ _18648_/Q _19239_/Q _19401_/Q _18616_/Q _10690_/X _10691_/X vssd1 vssd1 vccd1
+ vccd1 _11366_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13127__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13104_ _19711_/Q _12989_/X _12990_/X _16727_/B _13103_/X vssd1 vssd1 vccd1 vccd1
+ _13104_/X sky130_fd_sc_hd__a221o_1
XFILLER_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10316_ _19472_/Q _19310_/Q _18719_/Q _18489_/Q _10302_/X _09817_/A vssd1 vssd1 vccd1
+ vccd1 _10317_/B sky130_fd_sc_hd__mux4_1
XFILLER_140_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18961_ _19512_/CLK _18961_/D vssd1 vssd1 vccd1 vccd1 _18961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14084_ _14084_/A vssd1 vssd1 vccd1 vccd1 _18669_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output160_A _12495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11296_ _18636_/Q _19227_/Q _19389_/Q _18604_/Q _10977_/A _10006_/A vssd1 vssd1 vccd1
+ vccd1 _11296_/X sky130_fd_sc_hd__mux4_2
XFILLER_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13817__S _13829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13035_ _13035_/A vssd1 vssd1 vccd1 vccd1 _18470_/D sky130_fd_sc_hd__clkbuf_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ _17666_/S _17593_/X _17719_/X vssd1 vssd1 vccd1 vccd1 _17912_/Y sky130_fd_sc_hd__o21bai_2
X_10247_ _10196_/A _10244_/X _10246_/X vssd1 vssd1 vccd1 vccd1 _10247_/X sky130_fd_sc_hd__a21o_1
X_18892_ _19574_/CLK _18892_/D vssd1 vssd1 vccd1 vccd1 _18892_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_186_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17843_ _17843_/A vssd1 vssd1 vccd1 vccd1 _19902_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11845__B _19820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10897__C1 _09601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10178_ _18786_/Q _19057_/Q _19281_/Q _19025_/Q _09723_/A _09868_/A vssd1 vssd1 vccd1
+ vccd1 _10178_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17774_ _17612_/X _17770_/X _17773_/Y _17634_/X vssd1 vssd1 vccd1 vccd1 _17774_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14986_ _14986_/A vssd1 vssd1 vccd1 vccd1 _19032_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12102__A2 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19513_ _19575_/CLK _19513_/D vssd1 vssd1 vccd1 vccd1 _19513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16725_ _16727_/B _16727_/C _16724_/Y vssd1 vssd1 vccd1 vccd1 _19679_/D sky130_fd_sc_hd__o21a_1
X_13937_ _18606_/Q _13626_/X _13939_/S vssd1 vssd1 vccd1 vccd1 _13938_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14648__S _14654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19444_ _19508_/CLK _19444_/D vssd1 vssd1 vccd1 vccd1 _19444_/Q sky130_fd_sc_hd__dfxtp_1
X_13868_ _13868_/A vssd1 vssd1 vccd1 vccd1 _18575_/D sky130_fd_sc_hd__clkbuf_1
X_16656_ _16656_/A vssd1 vssd1 vccd1 vccd1 _16661_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12819_ _13595_/A _12796_/X _12856_/A vssd1 vssd1 vccd1 vccd1 _12819_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15607_ _14599_/X _19297_/Q _15611_/S vssd1 vssd1 vccd1 vccd1 _15608_/A sky130_fd_sc_hd__mux2_1
X_19375_ _19566_/CLK _19375_/D vssd1 vssd1 vccd1 vccd1 _19375_/Q sky130_fd_sc_hd__dfxtp_1
X_13799_ _14624_/A vssd1 vssd1 vccd1 vccd1 _13799_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16587_ _19636_/Q _16590_/C _16577_/X vssd1 vssd1 vccd1 vccd1 _16587_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18326_ _18326_/A _18326_/B vssd1 vssd1 vccd1 vccd1 _18326_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11613__A1 _11665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _15538_/A vssd1 vssd1 vccd1 vccd1 _19266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15469_ _15515_/S vssd1 vssd1 vccd1 vccd1 _15478_/S sky130_fd_sc_hd__clkbuf_4
X_18257_ _18257_/A vssd1 vssd1 vccd1 vccd1 _19982_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14383__S _14386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13366__B2 _19534_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17208_ _15770_/X _17197_/X _17207_/X _17201_/X vssd1 vssd1 vccd1 vccd1 _19836_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18188_ _16347_/B _19984_/Q _18192_/S vssd1 vssd1 vccd1 vccd1 _18189_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10416__S _10416_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17139_ _19814_/Q _12880_/X _17138_/X _16480_/X vssd1 vssd1 vccd1 vccd1 _19814_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11472__S0 _09532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09961_ _11478_/A vssd1 vssd1 vccd1 vccd1 _11475_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09892_ _10233_/A _09890_/X _09891_/X vssd1 vssd1 vccd1 vccd1 _09892_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09506__A _10245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09326_ _19884_/Q vssd1 vssd1 vccd1 vccd1 _13578_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_167_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13698__A _13719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09257_ _11645_/B _09307_/B vssd1 vssd1 vccd1 vccd1 _11789_/A sky130_fd_sc_hd__nand2_2
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ _17331_/A _09269_/D vssd1 vssd1 vccd1 vccd1 _09188_/Y sky130_fd_sc_hd__nor2_4
XFILLER_146_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11150_ _10024_/A _11149_/X _11170_/A vssd1 vssd1 vccd1 vccd1 _11150_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_162_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10101_ _10630_/A _10098_/X _10100_/X _10621_/A vssd1 vssd1 vccd1 vccd1 _10101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10850__A _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__S0 _11085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ _10875_/X _11073_/X _11075_/X _11080_/X _09600_/A vssd1 vssd1 vccd1 vccd1
+ _11081_/X sky130_fd_sc_hd__a311o_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11135__A3 _11134_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10032_ _10014_/X _10021_/Y _10030_/Y _10648_/A vssd1 vssd1 vccd1 vccd1 _10032_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11665__B _11665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14840_ _18359_/A _18406_/B vssd1 vssd1 vccd1 vccd1 _18968_/D sky130_fd_sc_hd__nor2_4
XANTENNA__17354__A2_N _17342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14771_ _18940_/Q _14395_/X _14775_/S vssd1 vssd1 vccd1 vccd1 _14772_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input17_A io_dbus_rdata[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11983_ _19824_/Q _11982_/X _16213_/A vssd1 vssd1 vccd1 vccd1 _11984_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11681__A _12602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ _15283_/A vssd1 vssd1 vccd1 vccd1 _14660_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16510_ _17101_/A vssd1 vssd1 vccd1 vccd1 _16550_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ _09998_/A _10923_/X _10932_/X _10065_/A _10933_/Y vssd1 vssd1 vccd1 vccd1
+ _12643_/A sky130_fd_sc_hd__o32a_4
X_17490_ _17487_/X _17488_/X _17590_/S vssd1 vssd1 vccd1 vccd1 _17490_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13653_ _13653_/A vssd1 vssd1 vccd1 vccd1 _18516_/D sky130_fd_sc_hd__clkbuf_1
X_16441_ _13557_/X _19577_/Q _16441_/S vssd1 vssd1 vccd1 vccd1 _16442_/A sky130_fd_sc_hd__mux2_1
X_10865_ _10858_/Y _10860_/Y _10862_/Y _10864_/Y _10063_/X vssd1 vssd1 vccd1 vccd1
+ _10865_/X sky130_fd_sc_hd__o221a_1
XFILLER_140_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _12604_/A _12604_/B _18009_/A vssd1 vssd1 vccd1 vccd1 _12609_/C sky130_fd_sc_hd__or3_1
XFILLER_158_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _16428_/A vssd1 vssd1 vccd1 vccd1 _16441_/S sky130_fd_sc_hd__buf_4
X_19160_ _19398_/CLK _19160_/D vssd1 vssd1 vccd1 vccd1 _19160_/Q sky130_fd_sc_hd__dfxtp_1
X_13584_ _12421_/X _11842_/B _13583_/Y vssd1 vssd1 vccd1 vccd1 _13584_/X sky130_fd_sc_hd__a21o_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _10652_/A _10795_/X _09693_/A vssd1 vssd1 vccd1 vccd1 _10796_/Y sky130_fd_sc_hd__o21ai_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15299__S _15299_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18111_ _18111_/A _18111_/B vssd1 vssd1 vccd1 vccd1 _18111_/Y sky130_fd_sc_hd__nor2_1
X_15323_ _19171_/Q _15228_/X _15323_/S vssd1 vssd1 vccd1 vccd1 _15324_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _12535_/A _12535_/B vssd1 vssd1 vccd1 vccd1 _12536_/A sky130_fd_sc_hd__nand2_2
X_19091_ _19571_/CLK _19091_/D vssd1 vssd1 vccd1 vccd1 _19091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15254_ _15254_/A vssd1 vssd1 vccd1 vccd1 _15254_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18042_ _19916_/Q _18019_/X _18041_/X vssd1 vssd1 vccd1 vccd1 _19916_/D sky130_fd_sc_hd__o21a_1
X_12466_ _12466_/A _12511_/C vssd1 vssd1 vccd1 vccd1 _12466_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14205_ _13825_/X _18722_/Q _14207_/S vssd1 vssd1 vccd1 vccd1 _14206_/A sky130_fd_sc_hd__mux2_1
X_11417_ _11560_/A _11563_/A _11560_/C _10460_/A _11416_/Y vssd1 vssd1 vccd1 vccd1
+ _11556_/C sky130_fd_sc_hd__a311o_1
XANTENNA__10257__S1 _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15185_ _19124_/Q vssd1 vssd1 vccd1 vccd1 _15186_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__14931__S _14939_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12017__A _17832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12397_ _12208_/X _12395_/X _12396_/X vssd1 vssd1 vccd1 vccd1 _12397_/X sky130_fd_sc_hd__o21a_1
XANTENNA_output85_A _12391_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14136_ _18693_/Q _13723_/X _14142_/S vssd1 vssd1 vccd1 vccd1 _14137_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ _11348_/A _12633_/B vssd1 vssd1 vccd1 vccd1 _11348_/Y sky130_fd_sc_hd__nor2_1
X_19993_ _20027_/CLK _19993_/D vssd1 vssd1 vccd1 vccd1 _19993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18944_ _19495_/CLK _18944_/D vssd1 vssd1 vccd1 vccd1 _18944_/Q sky130_fd_sc_hd__dfxtp_1
X_14067_ _14067_/A vssd1 vssd1 vccd1 vccd1 _18663_/D sky130_fd_sc_hd__clkbuf_1
X_11279_ _11291_/A _11279_/B vssd1 vssd1 vccd1 vccd1 _11279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13018_ _13454_/A vssd1 vssd1 vccd1 vccd1 _13558_/S sky130_fd_sc_hd__buf_4
XANTENNA__13520__A1 _13519_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18875_ _19301_/CLK _18875_/D vssd1 vssd1 vccd1 vccd1 _18875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17826_ _19901_/Q _17758_/X _17825_/X vssd1 vssd1 vccd1 vccd1 _19901_/D sky130_fd_sc_hd__o21a_1
XFILLER_94_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11509__S1 _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16470__B1 _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13284__B1 _13343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17757_ _19898_/Q _09419_/X _17753_/X _17756_/X vssd1 vssd1 vccd1 vccd1 _19898_/D
+ sky130_fd_sc_hd__o22a_1
X_14969_ _14969_/A vssd1 vssd1 vccd1 vccd1 _19024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15063__A _15131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16708_ _19674_/Q _16708_/B _17123_/B vssd1 vssd1 vccd1 vccd1 _16709_/C sky130_fd_sc_hd__and3_1
XFILLER_23_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17688_ _17688_/A vssd1 vssd1 vccd1 vccd1 _17930_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19427_ _19553_/CLK _19427_/D vssd1 vssd1 vccd1 vccd1 _19427_/Q sky130_fd_sc_hd__dfxtp_1
X_16639_ _16783_/A vssd1 vssd1 vccd1 vccd1 _16674_/A sky130_fd_sc_hd__buf_2
XFILLER_90_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10000__A _10655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19358_ _19666_/CLK _19358_/D vssd1 vssd1 vccd1 vccd1 _19358_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16606__B _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18309_ _20003_/Q _18285_/X _18308_/Y _18303_/X vssd1 vssd1 vccd1 vccd1 _20003_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19289_ _19952_/CLK _19289_/D vssd1 vssd1 vccd1 vccd1 _19289_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10935__A _11355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10248__S1 _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15238__A _15238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ _19917_/Q vssd1 vssd1 vccd1 vccd1 _09944_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09875_ _18596_/Q _18857_/Q _18756_/Q _19091_/Q _09872_/X _09874_/X vssd1 vssd1 vccd1
+ vccd1 _09875_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A io_dbus_rdata[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10420__S1 _10291_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14288__S _14290_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__B1 _13026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17961__B1 _17607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13920__S _13922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_134_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ _18585_/Q _18846_/Q _18745_/Q _19080_/Q _10649_/X _10014_/X vssd1 vssd1 vccd1
+ vccd1 _10651_/B sky130_fd_sc_hd__mux4_1
XFILLER_167_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09877__S0 _10173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09309_ _20042_/Q _14148_/A vssd1 vssd1 vccd1 vccd1 _09309_/X sky130_fd_sc_hd__xor2_1
XFILLER_139_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12250__A1 _18316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__A2 _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _10583_/A _10580_/X _09694_/A vssd1 vssd1 vccd1 vccd1 _10581_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10487__S1 _10333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12320_ _12320_/A _12320_/B vssd1 vssd1 vccd1 vccd1 _12320_/X sky130_fd_sc_hd__or2_2
XFILLER_10_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ _12188_/A _12654_/B _12250_/Y vssd1 vssd1 vccd1 vccd1 _17964_/B sky130_fd_sc_hd__a21o_2
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11202_ _11202_/A _11202_/B vssd1 vssd1 vccd1 vccd1 _11202_/X sky130_fd_sc_hd__or2_1
XFILLER_134_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _12176_/Y _12180_/X _12181_/X vssd1 vssd1 vccd1 vccd1 _12182_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11133_ _11304_/A _11130_/X _11132_/X _11069_/X vssd1 vssd1 vccd1 vccd1 _11133_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16990_ _16994_/C _16992_/C _16989_/Y vssd1 vssd1 vccd1 vccd1 _19754_/D sky130_fd_sc_hd__o21a_1
XFILLER_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11064_ _18966_/Q vssd1 vssd1 vccd1 vccd1 _11065_/A sky130_fd_sc_hd__buf_4
XFILLER_62_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15941_ _15941_/A vssd1 vssd1 vccd1 vccd1 _19397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09801__S0 _09724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_59_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13891__A _13913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _11280_/S vssd1 vssd1 vccd1 vccd1 _10977_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18660_ _19569_/CLK _18660_/D vssd1 vssd1 vccd1 vccd1 _18660_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17244__A2 _17197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15872_ _15872_/A vssd1 vssd1 vccd1 vccd1 _19366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17611_ _17849_/A _17608_/A _18110_/S _17610_/X vssd1 vssd1 vccd1 vccd1 _17611_/X
+ sky130_fd_sc_hd__o211a_1
X_14823_ _18964_/Q _14471_/X _14823_/S vssd1 vssd1 vccd1 vccd1 _14824_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18591_ _19311_/CLK _18591_/D vssd1 vssd1 vccd1 vccd1 _18591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output123_A _12660_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17542_ _17542_/A _17545_/B _17549_/A _17542_/D vssd1 vssd1 vccd1 vccd1 _17785_/A
+ sky130_fd_sc_hd__and4_1
X_14754_ _14810_/A vssd1 vssd1 vccd1 vccd1 _14823_/S sky130_fd_sc_hd__buf_6
X_11966_ _11966_/A vssd1 vssd1 vccd1 vccd1 _12077_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ _15270_/A vssd1 vssd1 vccd1 vccd1 _14647_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10917_ _10917_/A vssd1 vssd1 vccd1 vccd1 _10969_/A sky130_fd_sc_hd__buf_4
X_14685_ _18897_/Q _14376_/X _14691_/S vssd1 vssd1 vccd1 vccd1 _14686_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17473_ _17443_/X _17470_/X _17845_/A vssd1 vssd1 vccd1 vccd1 _17473_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14926__S _14928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11897_ _11961_/A _12633_/B _11756_/Y vssd1 vssd1 vccd1 vccd1 _17739_/S sky130_fd_sc_hd__o21a_1
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19212_ _19564_/CLK _19212_/D vssd1 vssd1 vccd1 vccd1 _19212_/Q sky130_fd_sc_hd__dfxtp_1
X_16424_ _13423_/X _19569_/Q _16426_/S vssd1 vssd1 vccd1 vccd1 _16425_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13636_ _18512_/Q _13634_/X _13652_/S vssd1 vssd1 vccd1 vccd1 _13637_/A sky130_fd_sc_hd__mux2_1
X_10848_ _10848_/A vssd1 vssd1 vccd1 vccd1 _10848_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19143_ _19401_/CLK _19143_/D vssd1 vssd1 vccd1 vccd1 _19143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13567_ _13567_/A vssd1 vssd1 vccd1 vccd1 _18501_/D sky130_fd_sc_hd__clkbuf_1
X_16355_ _12215_/X _15828_/X _16223_/S vssd1 vssd1 vccd1 vccd1 _16355_/X sky130_fd_sc_hd__a21bo_1
XFILLER_157_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10779_ _18805_/Q _19140_/Q _11386_/S vssd1 vssd1 vccd1 vccd1 _10779_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15306_ _19163_/Q _15203_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _15307_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12792__A2 _15764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12518_ _12421_/X _12516_/X _12517_/Y _12131_/X vssd1 vssd1 vccd1 vccd1 _12518_/X
+ sky130_fd_sc_hd__a31o_1
X_16286_ _16369_/S vssd1 vssd1 vccd1 vccd1 _16325_/S sky130_fd_sc_hd__clkbuf_2
X_19074_ _19074_/CLK _19074_/D vssd1 vssd1 vccd1 vccd1 _19074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13498_ _19352_/Q _13245_/X _13099_/X _19542_/Q _13497_/X vssd1 vssd1 vccd1 vccd1
+ _13498_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18025_ _17612_/X _18022_/X _18024_/Y _17705_/A vssd1 vssd1 vccd1 vccd1 _18025_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15757__S _15757_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15237_ _15237_/A vssd1 vssd1 vccd1 vccd1 _19141_/D sky130_fd_sc_hd__clkbuf_1
X_12449_ _18336_/A _12475_/B vssd1 vssd1 vccd1 vccd1 _12449_/X sky130_fd_sc_hd__or2_2
XANTENNA__14661__S _14670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15168_ _15168_/A vssd1 vssd1 vccd1 vccd1 _19115_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14119_ _14119_/A vssd1 vssd1 vccd1 vccd1 _18685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15099_ _14628_/X _19082_/Q _15105_/S vssd1 vssd1 vccd1 vccd1 _15100_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19976_ _19978_/CLK _19976_/D vssd1 vssd1 vccd1 vccd1 _19976_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10650__S1 _10014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18927_ _19129_/CLK _18927_/D vssd1 vssd1 vccd1 vccd1 _18927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18369__A _18380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09660_ _09660_/A vssd1 vssd1 vccd1 vccd1 _10105_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10402__S1 _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18858_ _19092_/CLK _18858_/D vssd1 vssd1 vccd1 vccd1 _18858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17809_ _17809_/A vssd1 vssd1 vccd1 vccd1 _19900_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17640__C1 _17543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09591_ _09773_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09591_/X sky130_fd_sc_hd__or2_1
X_18789_ _19285_/CLK _18789_/D vssd1 vssd1 vccd1 vccd1 _18789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13740__S _13744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09859__S0 _10175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14509__A0 _13758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16352__A _19953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18120__B1 _17543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11496__A _11496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09927_ _09927_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _09927_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_60_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17183__A _17242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09858_ _09858_/A vssd1 vssd1 vccd1 vccd1 _09858_/X sky130_fd_sc_hd__clkbuf_4
X_20047_ _20048_/CLK _20047_/D vssd1 vssd1 vccd1 vccd1 _20047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _09788_/A _09786_/Y _09788_/Y _09800_/A vssd1 vssd1 vccd1 vccd1 _09789_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11818_/X _11819_/X _11816_/A vssd1 vssd1 vccd1 vccd1 _11820_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11751_ _11856_/S _12632_/B _11708_/Y vssd1 vssd1 vccd1 vccd1 _17467_/A sky130_fd_sc_hd__o21ai_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14746__S _14746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _18807_/Q _19142_/Q _10702_/S vssd1 vssd1 vccd1 vccd1 _10703_/B sky130_fd_sc_hd__mux2_1
XFILLER_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14470_ _14470_/A vssd1 vssd1 vccd1 vccd1 _18825_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11682_/A _11682_/B vssd1 vssd1 vccd1 vccd1 _17394_/C sky130_fd_sc_hd__nand2_1
XFILLER_42_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ input16/X _13303_/X _13306_/X vssd1 vssd1 vccd1 vccd1 _13421_/Y sky130_fd_sc_hd__a21oi_1
X_10633_ _19466_/Q _19304_/Q _18713_/Q _18483_/Q _10678_/S _09813_/A vssd1 vssd1 vccd1
+ vccd1 _10633_/X sky130_fd_sc_hd__mux4_1
X_16140_ _16140_/A vssd1 vssd1 vccd1 vccd1 _19485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13352_ _13337_/X _13350_/X _13351_/X vssd1 vssd1 vccd1 vccd1 _13352_/Y sky130_fd_sc_hd__a21oi_1
X_10564_ _18586_/Q _18847_/Q _18746_/Q _19081_/Q _11428_/S _09814_/A vssd1 vssd1 vccd1
+ vccd1 _10565_/B sky130_fd_sc_hd__mux4_1
XFILLER_128_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15577__S _15583_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _19976_/Q _11415_/A _12303_/S vssd1 vssd1 vccd1 vccd1 _12331_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16071_ _13069_/X _19455_/Q _16073_/S vssd1 vssd1 vccd1 vccd1 _16072_/A sky130_fd_sc_hd__mux2_1
X_13283_ _13282_/A _13297_/C _13038_/A vssd1 vssd1 vccd1 vccd1 _13283_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10495_ _10495_/A vssd1 vssd1 vccd1 vccd1 _10495_/Y sky130_fd_sc_hd__inv_2
X_15022_ _19048_/Q _14417_/X _15022_/S vssd1 vssd1 vccd1 vccd1 _15023_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12234_ _12538_/A _12234_/B vssd1 vssd1 vccd1 vccd1 _12234_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19830_ _19865_/CLK _19830_/D vssd1 vssd1 vccd1 vccd1 _19830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12165_ _17918_/B _12165_/B vssd1 vssd1 vccd1 vccd1 _12169_/A sky130_fd_sc_hd__xor2_1
XFILLER_111_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11116_ _11116_/A vssd1 vssd1 vccd1 vccd1 _11271_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19761_ _19762_/CLK _19761_/D vssd1 vssd1 vccd1 vccd1 _19761_/Q sky130_fd_sc_hd__dfxtp_1
X_12096_ _12096_/A vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__clkbuf_1
X_16973_ _16993_/A _16973_/B _16978_/C vssd1 vssd1 vccd1 vccd1 _19749_/D sky130_fd_sc_hd__nor3_1
XFILLER_122_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18712_ _18845_/CLK _18712_/D vssd1 vssd1 vccd1 vccd1 _18712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15924_ _15924_/A vssd1 vssd1 vccd1 vccd1 _19389_/D sky130_fd_sc_hd__clkbuf_1
X_11047_ _18641_/Q _19232_/Q _19394_/Q _18609_/Q _10018_/A _10974_/X vssd1 vssd1 vccd1
+ vccd1 _11047_/X sky130_fd_sc_hd__mux4_1
X_19692_ _19726_/CLK _19692_/D vssd1 vssd1 vccd1 vccd1 _19692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput9 io_dbus_rdata[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_4
XFILLER_37_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09604__A _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18643_ _19493_/CLK _18643_/D vssd1 vssd1 vccd1 vccd1 _18643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15855_ _13069_/X _19359_/Q _15857_/S vssd1 vssd1 vccd1 vccd1 _15856_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14806_ _18956_/Q _14446_/X _14808_/S vssd1 vssd1 vccd1 vccd1 _14807_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18574_ _19391_/CLK _18574_/D vssd1 vssd1 vccd1 vccd1 _18574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15786_ _15785_/X _19345_/Q _15801_/S vssd1 vssd1 vccd1 vccd1 _15787_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12998_ _19706_/Q _12989_/X _12990_/X _19674_/Q _12997_/X vssd1 vssd1 vccd1 vccd1
+ _12998_/X sky130_fd_sc_hd__a221o_1
XFILLER_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17525_ _17525_/A _17802_/C vssd1 vssd1 vccd1 vccd1 _17603_/A sky130_fd_sc_hd__and2_1
X_14737_ _14737_/A vssd1 vssd1 vccd1 vccd1 _14746_/S sky130_fd_sc_hd__buf_4
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11949_ _19823_/Q _11950_/B vssd1 vssd1 vccd1 vccd1 _11951_/A sky130_fd_sc_hd__and2_1
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17925__B1 _12175_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17456_ _17449_/X _17455_/X _17685_/S vssd1 vssd1 vccd1 vccd1 _17456_/X sky130_fd_sc_hd__mux2_1
X_14668_ _14668_/A vssd1 vssd1 vccd1 vccd1 _18892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16407_ _13293_/X _19561_/Q _16415_/S vssd1 vssd1 vccd1 vccd1 _16408_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _18508_/Q _13618_/X _13631_/S vssd1 vssd1 vccd1 vccd1 _13620_/A sky130_fd_sc_hd__mux2_1
X_17387_ _18118_/B _17668_/A vssd1 vssd1 vccd1 vccd1 _17387_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14599_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14599_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19126_ _19574_/CLK _19126_/D vssd1 vssd1 vccd1 vccd1 _19126_/Q sky130_fd_sc_hd__dfxtp_1
X_16338_ _19950_/Q _16338_/B vssd1 vssd1 vccd1 vccd1 _16338_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13796__A _14621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15487__S _15489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19057_ _19507_/CLK _19057_/D vssd1 vssd1 vccd1 vccd1 _19057_/Q sky130_fd_sc_hd__dfxtp_1
X_16269_ _12874_/X _16267_/Y _16318_/S vssd1 vssd1 vccd1 vccd1 _16269_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18008_ _18012_/A _18012_/B vssd1 vssd1 vccd1 vccd1 _18008_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19959_ _19997_/CLK _19959_/D vssd1 vssd1 vccd1 vccd1 _19959_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ _09712_/A vssd1 vssd1 vccd1 vccd1 _09712_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16111__S _16117_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14420__A _14624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ _10968_/S vssd1 vssd1 vccd1 vccd1 _10909_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _09574_/A vssd1 vssd1 vccd1 vccd1 _09975_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14566__S _14568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16347__A _16347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15251__A _15251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09606__C1 _09605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18281__B _18281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ _19505_/Q _18917_/Q _18954_/Q _18528_/Q _10216_/S _09858_/A vssd1 vssd1 vccd1
+ vccd1 _10280_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13181__A2 _13172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10334__S _10439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11192__A1 _09954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _20027_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16021__S _16023_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13970_ _18621_/Q _13689_/X _13972_/S vssd1 vssd1 vccd1 vccd1 _13971_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12141__A0 _19970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _19666_/Q _12887_/A _12889_/A _19798_/Q _12920_/X vssd1 vssd1 vccd1 vccd1
+ _12921_/X sky130_fd_sc_hd__a221o_2
XFILLER_46_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15640_ _14647_/X _19312_/Q _15644_/S vssd1 vssd1 vccd1 vccd1 _15641_/A sky130_fd_sc_hd__mux2_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12852_ _15680_/A _18448_/Q vssd1 vssd1 vccd1 vccd1 _12852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10289__B _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _20031_/Q _11854_/B vssd1 vssd1 vccd1 vccd1 _11803_/X sky130_fd_sc_hd__or2_1
X_15571_ _15571_/A vssd1 vssd1 vccd1 vccd1 _19281_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _19807_/Q _12684_/C _12696_/A _17205_/A _12782_/X vssd1 vssd1 vccd1 vccd1
+ _12783_/X sky130_fd_sc_hd__a221o_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17310_ _17310_/A vssd1 vssd1 vccd1 vccd1 _19877_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _12320_/A _11690_/X _11693_/X _11695_/X vssd1 vssd1 vccd1 vccd1 _11734_/X
+ sky130_fd_sc_hd__a31o_1
X_14522_ _13777_/X _18840_/Q _14524_/S vssd1 vssd1 vccd1 vccd1 _14523_/A sky130_fd_sc_hd__mux2_1
X_18290_ _14501_/B _18285_/X _18288_/X _18289_/X vssd1 vssd1 vccd1 vccd1 _19996_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _15839_/X _17229_/X _17240_/X _17232_/X vssd1 vssd1 vccd1 vccd1 _19847_/D
+ sky130_fd_sc_hd__o211a_1
X_14453_ _14453_/A vssd1 vssd1 vccd1 vccd1 _14466_/S sky130_fd_sc_hd__buf_4
X_11665_ _19323_/D _11665_/B vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10509__S _10509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10616_ _18777_/Q _19048_/Q _19272_/Q _19016_/Q _10614_/X _11371_/A vssd1 vssd1 vccd1
+ vccd1 _10616_/X sky130_fd_sc_hd__mux4_2
X_13404_ _19760_/Q _12892_/X _13403_/X _12896_/X vssd1 vssd1 vccd1 vccd1 _13404_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_174_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17172_ _17166_/Y _17167_/X _17170_/X _17171_/X vssd1 vssd1 vccd1 vccd1 _19823_/D
+ sky130_fd_sc_hd__o211a_1
X_14384_ _14384_/A vssd1 vssd1 vccd1 vccd1 _18798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11596_ _10139_/X _11545_/A _11545_/B vssd1 vssd1 vccd1 vccd1 _11596_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16123_ _16123_/A vssd1 vssd1 vccd1 vccd1 _19478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13335_ _19943_/Q _19944_/Q _13335_/C vssd1 vssd1 vccd1 vccd1 _13362_/B sky130_fd_sc_hd__and3_1
X_10547_ _18651_/Q _19242_/Q _19404_/Q _18619_/Q _10337_/A _09855_/A vssd1 vssd1 vccd1
+ vccd1 _10548_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10853__S1 _10037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15697__A1 _19899_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16054_ _13506_/X _19448_/Q _16056_/S vssd1 vssd1 vccd1 vccd1 _16055_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13266_ _19752_/Q _12991_/X _13265_/X _12995_/X vssd1 vssd1 vccd1 vccd1 _13266_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10478_ _10478_/A _10478_/B vssd1 vssd1 vccd1 vccd1 _10478_/X sky130_fd_sc_hd__or2_1
X_12217_ _19832_/Q _19831_/Q _12217_/C vssd1 vssd1 vccd1 vccd1 _12267_/C sky130_fd_sc_hd__and3_2
X_15005_ _19040_/Q _14392_/X _15011_/S vssd1 vssd1 vccd1 vccd1 _15006_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10244__S _10244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13197_ _13197_/A vssd1 vssd1 vccd1 vccd1 _18478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12380__B1 _12429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19813_ _20044_/CLK _19813_/D vssd1 vssd1 vccd1 vccd1 _19813_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ _12148_/A vssd1 vssd1 vccd1 vccd1 _12148_/Y sky130_fd_sc_hd__inv_6
XFILLER_111_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11255__A2_N _11348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__A _11864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15336__A _15358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19744_ _19745_/CLK _19744_/D vssd1 vssd1 vccd1 vccd1 _19744_/Q sky130_fd_sc_hd__dfxtp_1
X_16956_ _16993_/A _16956_/B _16971_/C vssd1 vssd1 vccd1 vccd1 _19745_/D sky130_fd_sc_hd__nor3_1
X_12079_ _12079_/A vssd1 vssd1 vccd1 vccd1 _12081_/A sky130_fd_sc_hd__inv_2
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15907_ _15907_/A vssd1 vssd1 vccd1 vccd1 _19382_/D sky130_fd_sc_hd__clkbuf_1
X_19675_ _19682_/CLK _19675_/D vssd1 vssd1 vccd1 vccd1 _19675_/Q sky130_fd_sc_hd__dfxtp_1
X_16887_ _16922_/B _16891_/D _19727_/Q vssd1 vssd1 vccd1 vccd1 _16889_/B sky130_fd_sc_hd__a21oi_1
XFILLER_37_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18626_ _19411_/CLK _18626_/D vssd1 vssd1 vccd1 vccd1 _18626_/Q sky130_fd_sc_hd__dfxtp_1
X_15838_ _18467_/Q _13533_/X _15837_/Y _13587_/A vssd1 vssd1 vccd1 vccd1 _15838_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11891__C1 _16487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18557_ _19564_/CLK _18557_/D vssd1 vssd1 vccd1 vccd1 _18557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12695__A _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14386__S _14386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15769_ _15783_/A _18456_/Q vssd1 vssd1 vccd1 vccd1 _15769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17508_ _17506_/X _17507_/X _17508_/S vssd1 vssd1 vccd1 vccd1 _17508_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09290_ _19996_/Q _20036_/Q vssd1 vssd1 vccd1 vccd1 _09290_/X sky130_fd_sc_hd__or2b_1
X_18488_ _19470_/CLK _18488_/D vssd1 vssd1 vccd1 vccd1 _18488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17439_ _17433_/X _17437_/X _17802_/D vssd1 vssd1 vccd1 vccd1 _17439_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10749__A1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__B2 _19904_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19109_ _19557_/CLK _19109_/D vssd1 vssd1 vccd1 vccd1 _19109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16106__S _16106_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10943__A _11260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_opt_2_0_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput110 _12646_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[10] sky130_fd_sc_hd__buf_2
Xoutput121 _12657_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[20] sky130_fd_sc_hd__buf_2
XANTENNA__15945__S _15951_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput132 _12669_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[30] sky130_fd_sc_hd__buf_2
XFILLER_115_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput143 _16465_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[10] sky130_fd_sc_hd__buf_2
Xoutput154 _12348_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[20] sky130_fd_sc_hd__buf_2
Xoutput165 _12590_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[30] sky130_fd_sc_hd__buf_2
XFILLER_130_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09626_ _11096_/A vssd1 vssd1 vccd1 vccd1 _11291_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09557_ _10606_/A vssd1 vssd1 vccd1 vccd1 _10630_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12426__B2 _12425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11713__S _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09488_ _10569_/A vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10329__S _10496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11014__A _11014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11450_ _11450_/A vssd1 vssd1 vccd1 vccd1 _11450_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11088__S1 _10917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10401_ _09891_/A _10389_/Y _10394_/X _10400_/Y _09741_/A vssd1 vssd1 vccd1 vccd1
+ _10401_/X sky130_fd_sc_hd__o311a_1
XANTENNA__11949__A _19823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _11369_/X _11380_/Y hold15/A _09996_/X vssd1 vssd1 vccd1 vccd1 _11406_/A
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__10835__S1 _09970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _19330_/Q _13154_/A _13562_/A _19520_/Q _13119_/X vssd1 vssd1 vccd1 vccd1
+ _13120_/X sky130_fd_sc_hd__a221o_1
X_10332_ _10332_/A vssd1 vssd1 vccd1 vccd1 _10333_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_124_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15855__S _15857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ _13299_/C _13051_/B vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__or2_1
X_10263_ _19119_/Q _18885_/Q _19567_/Q _19215_/Q _10216_/S _09858_/A vssd1 vssd1 vccd1
+ vccd1 _10264_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12002_ _12002_/A _12002_/B vssd1 vssd1 vccd1 vccd1 _12003_/A sky130_fd_sc_hd__xnor2_4
XFILLER_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input47_A io_ibus_inst[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10194_ _11421_/A _12661_/B vssd1 vssd1 vccd1 vccd1 _11539_/A sky130_fd_sc_hd__or2_1
X_16810_ _11952_/C _13748_/B _16807_/X _16809_/X vssd1 vssd1 vccd1 vccd1 _16816_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_120_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17790_ _17786_/Y _17788_/X _18089_/S vssd1 vssd1 vccd1 vccd1 _17790_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16741_ _16749_/D vssd1 vssd1 vccd1 vccd1 _16747_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13953_ _18613_/Q _13655_/X _13961_/S vssd1 vssd1 vccd1 vccd1 _13954_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_163_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19792_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _12735_/X _12901_/X _12902_/Y _12903_/X _18460_/Q vssd1 vssd1 vccd1 vccd1
+ _17220_/A sky130_fd_sc_hd__a32oi_4
XFILLER_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19460_ _19552_/CLK _19460_/D vssd1 vssd1 vccd1 vccd1 _19460_/Q sky130_fd_sc_hd__dfxtp_1
X_16672_ _16672_/A _16672_/B _16672_/C vssd1 vssd1 vccd1 vccd1 _19665_/D sky130_fd_sc_hd__nor3_1
X_13884_ _13884_/A vssd1 vssd1 vccd1 vccd1 _18582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18411_ _18412_/A _18411_/B vssd1 vssd1 vccd1 vccd1 _20044_/D sky130_fd_sc_hd__nor2_1
X_15623_ _15623_/A vssd1 vssd1 vccd1 vccd1 _19304_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _19685_/Q vssd1 vssd1 vccd1 vccd1 _16747_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19391_ _19391_/CLK _19391_/D vssd1 vssd1 vccd1 vccd1 _19391_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _09389_/A _18302_/B _18340_/X _18341_/X vssd1 vssd1 vccd1 vccd1 _20016_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_178_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19879_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15554_ _15554_/A vssd1 vssd1 vccd1 vccd1 _19273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12766_ _13578_/A vssd1 vssd1 vccd1 vccd1 _15837_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _13746_/X _18832_/Q _14513_/S vssd1 vssd1 vccd1 vccd1 _14506_/A sky130_fd_sc_hd__mux2_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _09328_/C _19990_/Q _18273_/S vssd1 vssd1 vccd1 vccd1 _18274_/B sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_182_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11717_/A _11717_/B vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__nand2_2
X_15485_ _19243_/Q _15254_/X _15489_/S vssd1 vssd1 vccd1 vccd1 _15486_/A sky130_fd_sc_hd__mux2_1
X_12697_ _12697_/A vssd1 vssd1 vccd1 vccd1 _12992_/A sky130_fd_sc_hd__buf_2
XFILLER_159_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17224_ _15799_/Y _17212_/X _17223_/X _17215_/X vssd1 vssd1 vccd1 vccd1 _19841_/D
+ sky130_fd_sc_hd__o211a_1
X_14436_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14436_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11648_ _11648_/A _17331_/B _11648_/C vssd1 vssd1 vccd1 vccd1 _11692_/C sky130_fd_sc_hd__nor3_2
Xclkbuf_leaf_101_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19204_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput12 io_dbus_rdata[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_2
Xinput23 io_dbus_rdata[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_8
XFILLER_168_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput34 io_ibus_inst[0] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_6
Xinput45 io_ibus_inst[1] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_4
X_17155_ _17152_/Y _17153_/X _17154_/X _17142_/X vssd1 vssd1 vccd1 vccd1 _19818_/D
+ sky130_fd_sc_hd__o211a_1
X_11579_ _11579_/A _11579_/B vssd1 vssd1 vccd1 vccd1 _11579_/Y sky130_fd_sc_hd__nand2_1
X_14367_ _18794_/Q _13743_/X _14367_/S vssd1 vssd1 vccd1 vccd1 _14368_/A sky130_fd_sc_hd__mux2_1
Xinput56 io_ibus_inst[2] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput67 io_irq_motor_irq vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_4
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16106_ _13357_/X _19471_/Q _16106_/S vssd1 vssd1 vccd1 vccd1 _16107_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10600__B1 _09756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13318_ _13353_/A vssd1 vssd1 vccd1 vccd1 _13318_/X sky130_fd_sc_hd__clkbuf_2
X_14298_ _14354_/A vssd1 vssd1 vccd1 vccd1 _14367_/S sky130_fd_sc_hd__buf_6
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17086_ _17087_/B _17087_/C _17085_/Y vssd1 vssd1 vccd1 vccd1 _19790_/D sky130_fd_sc_hd__o21a_1
XFILLER_170_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16037_ _13376_/X _19440_/Q _16045_/S vssd1 vssd1 vccd1 vccd1 _16038_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_116_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19895_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13249_ _19623_/Q _13204_/X _13248_/X vssd1 vssd1 vccd1 vccd1 _13249_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16450__A _16678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__A1 _10920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09763__S _09763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11251__S1 _10943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10702__S _10702_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17988_ _18000_/A _17988_/B vssd1 vssd1 vccd1 vccd1 _17990_/C sky130_fd_sc_hd__nor2_1
XFILLER_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19727_ _19727_/CLK _19727_/D vssd1 vssd1 vccd1 vccd1 _19727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16939_ _16939_/A _16939_/B _16939_/C vssd1 vssd1 vccd1 vccd1 _16940_/A sky130_fd_sc_hd__and3_1
XFILLER_65_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18377__A _18380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19658_ _19792_/CLK _19658_/D vssd1 vssd1 vccd1 vccd1 _19658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10003__A _10909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09411_ _11774_/A vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__inv_2
XFILLER_52_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18609_ _19490_/CLK _18609_/D vssd1 vssd1 vccd1 vccd1 _18609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19589_ _19966_/CLK _19589_/D vssd1 vssd1 vccd1 vccd1 _19589_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10938__A _11001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ _19893_/Q vssd1 vssd1 vccd1 vccd1 _09342_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15005__S _15011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17347__B2 _15818_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09273_ _18279_/A _18276_/A _09328_/C _09328_/D vssd1 vssd1 vccd1 vccd1 _11682_/B
+ sky130_fd_sc_hd__and4b_2
XFILLER_20_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11700__A2_N _12631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11242__S1 _10943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_80_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19402_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15833__A1 _15818_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17035__B1 _17021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17191__A _17191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ _10955_/A _10946_/X _10948_/X _10949_/X vssd1 vssd1 vccd1 vccd1 _10951_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_95_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19572_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ _09617_/A _09609_/B vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__nor2_2
X_10881_ _11260_/A vssd1 vssd1 vccd1 vccd1 _11236_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12620_ _12620_/A _12620_/B vssd1 vssd1 vccd1 vccd1 _12620_/Y sky130_fd_sc_hd__nand2_4
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12551_ _18098_/B _12551_/B vssd1 vssd1 vccd1 vccd1 _12556_/A sky130_fd_sc_hd__xor2_1
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11502_ _10039_/A _11501_/X _10043_/A vssd1 vssd1 vccd1 vccd1 _11502_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15270_ _15270_/A vssd1 vssd1 vccd1 vccd1 _15270_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12482_ _12482_/A _12482_/B vssd1 vssd1 vccd1 vccd1 _12521_/C sky130_fd_sc_hd__nor2_1
XFILLER_138_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11433_ _18600_/Q _18861_/Q _18760_/Q _19095_/Q _10081_/X _10813_/A vssd1 vssd1 vccd1
+ vccd1 _11434_/B sky130_fd_sc_hd__mux4_1
X_14221_ _14221_/A vssd1 vssd1 vccd1 vccd1 _18729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12583__A0 _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19563_/CLK sky130_fd_sc_hd__clkbuf_16
X_14152_ _15918_/B _16062_/B vssd1 vssd1 vccd1 vccd1 _14209_/A sky130_fd_sc_hd__or2_4
XFILLER_4_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11364_ _10730_/A _11363_/X _09475_/A vssd1 vssd1 vccd1 vccd1 _11364_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10315_ _10378_/A _10313_/X _10314_/X vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__o21a_1
X_13103_ _16527_/B _12861_/X _13102_/X vssd1 vssd1 vccd1 vccd1 _13103_/X sky130_fd_sc_hd__o21a_1
XANTENNA__15585__S _15587_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18960_ _19092_/CLK _18960_/D vssd1 vssd1 vccd1 vccd1 _18960_/Q sky130_fd_sc_hd__dfxtp_1
X_14083_ _18669_/Q _13622_/X _14087_/S vssd1 vssd1 vccd1 vccd1 _14084_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11295_ _11295_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11295_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17911_ _11403_/Y _17861_/X _17910_/X vssd1 vssd1 vccd1 vccd1 _19906_/D sky130_fd_sc_hd__a21oi_1
X_13034_ _18470_/Q _13033_/X _13090_/S vssd1 vssd1 vccd1 vccd1 _13035_/A sky130_fd_sc_hd__mux2_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10246_ _10368_/A _10245_/X _09918_/A vssd1 vssd1 vccd1 vccd1 _10246_/X sky130_fd_sc_hd__a21o_1
X_18891_ _19573_/CLK _18891_/D vssd1 vssd1 vccd1 vccd1 _18891_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10346__C1 _09741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output153_A _16447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_129_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19507_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17274__A0 _12854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17842_ _19902_/Q _17840_/X _18085_/S vssd1 vssd1 vccd1 vccd1 _17843_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10177_ _10176_/A _10174_/Y _10176_/Y _09860_/A vssd1 vssd1 vccd1 vccd1 _10177_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17773_ _17771_/X _17768_/Y _17772_/Y vssd1 vssd1 vccd1 vccd1 _17773_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14985_ _19032_/Q _14468_/X _14987_/S vssd1 vssd1 vccd1 vccd1 _14986_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13833__S _13845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19512_ _19512_/CLK _19512_/D vssd1 vssd1 vccd1 vccd1 _19512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16724_ _16727_/B _16727_/C _16723_/X vssd1 vssd1 vccd1 vccd1 _16724_/Y sky130_fd_sc_hd__a21oi_1
X_13936_ _13936_/A vssd1 vssd1 vccd1 vccd1 _18605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10744__S0 _10614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19443_ _19443_/CLK _19443_/D vssd1 vssd1 vccd1 vccd1 _19443_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09612__A _09612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16655_ _16672_/A _16655_/B _16655_/C vssd1 vssd1 vccd1 vccd1 _19659_/D sky130_fd_sc_hd__nor3_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13867_ _13764_/X _18575_/Q _13867_/S vssd1 vssd1 vccd1 vccd1 _13868_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15606_ _15606_/A vssd1 vssd1 vccd1 vccd1 _19296_/D sky130_fd_sc_hd__clkbuf_1
X_19374_ _19565_/CLK _19374_/D vssd1 vssd1 vccd1 vccd1 _19374_/Q sky130_fd_sc_hd__dfxtp_1
X_12818_ _17247_/B _12818_/B _17149_/A vssd1 vssd1 vccd1 vccd1 _12856_/A sky130_fd_sc_hd__or3_1
XANTENNA__13063__A1 _16206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16586_ _19635_/Q _16584_/B _16585_/Y vssd1 vssd1 vccd1 vccd1 _19635_/D sky130_fd_sc_hd__o21a_1
X_13798_ _13798_/A vssd1 vssd1 vccd1 vccd1 _18553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18325_ _17146_/A _18323_/X _18324_/Y _18317_/X vssd1 vssd1 vccd1 vccd1 _20009_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ _19266_/Q _15225_/X _15539_/S vssd1 vssd1 vccd1 vccd1 _15538_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14664__S _14670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _16939_/A vssd1 vssd1 vccd1 vccd1 _12749_/X sky130_fd_sc_hd__buf_2
XANTENNA__12973__A _17861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18256_ _19982_/Q _19603_/Q _18264_/S vssd1 vssd1 vccd1 vccd1 _18257_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15468_ _15468_/A vssd1 vssd1 vccd1 vccd1 _19235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17207_ _19836_/Q _17210_/B vssd1 vssd1 vccd1 vccd1 _17207_/X sky130_fd_sc_hd__or2_1
X_14419_ _14419_/A vssd1 vssd1 vccd1 vccd1 _18809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18187_ _18187_/A vssd1 vssd1 vccd1 vccd1 _19951_/D sky130_fd_sc_hd__clkbuf_1
X_15399_ _15399_/A vssd1 vssd1 vccd1 vccd1 _19204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17138_ input69/X _17138_/B vssd1 vssd1 vccd1 vccd1 _17138_/X sky130_fd_sc_hd__or2_1
XFILLER_171_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17069_ _17070_/B _17070_/C _17068_/Y vssd1 vssd1 vccd1 vccd1 _19784_/D sky130_fd_sc_hd__o21a_1
X_09960_ _10955_/A vssd1 vssd1 vccd1 vccd1 _11478_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16180__A _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09891_ _09891_/A vssd1 vssd1 vccd1 vccd1 _09891_/X sky130_fd_sc_hd__clkbuf_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17265__A0 _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13309__A _15251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15815__A1 _19919_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17568__A1 _17484_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09522__A _09809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09325_ _09325_/A _09339_/B vssd1 vssd1 vccd1 vccd1 _09325_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12801__B2 _19517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09256_ _11675_/A _11678_/A vssd1 vssd1 vccd1 vccd1 _09307_/B sky130_fd_sc_hd__nor2_2
X_09187_ _09272_/A _09272_/C vssd1 vssd1 vccd1 vccd1 _09269_/D sky130_fd_sc_hd__or2_2
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12565__B1 _12421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18296__A2 _18291_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11463__S1 _10703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10576__C1 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13918__S _13922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10100_ _10817_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10100_/X sky130_fd_sc_hd__or2_1
XFILLER_122_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11080_ _11127_/A _11076_/X _11079_/X _11069_/X vssd1 vssd1 vccd1 vccd1 _11080_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11215__S1 _11164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_130_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17256__A0 _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10031_ _10116_/A vssd1 vssd1 vccd1 vccd1 _10648_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__13219__A _15231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12123__A _12492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14770_ _14770_/A vssd1 vssd1 vccd1 vccd1 _18939_/D sky130_fd_sc_hd__clkbuf_1
X_11982_ _11951_/A _11980_/Y _11957_/A vssd1 vssd1 vccd1 vccd1 _11982_/X sky130_fd_sc_hd__o21a_1
XFILLER_57_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13721_ _13721_/A vssd1 vssd1 vccd1 vccd1 _18532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10933_ _19901_/Q vssd1 vssd1 vccd1 vccd1 _10933_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16440_ _16440_/A vssd1 vssd1 vccd1 vccd1 _19576_/D sky130_fd_sc_hd__clkbuf_1
X_10864_ _11383_/A _10863_/X _09706_/A vssd1 vssd1 vccd1 vccd1 _10864_/Y sky130_fd_sc_hd__o21ai_1
X_13652_ _18516_/Q _13651_/X _13652_/S vssd1 vssd1 vccd1 vccd1 _13653_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _17323_/A _11600_/A _12601_/Y _18308_/A vssd1 vssd1 vccd1 vccd1 _18009_/A
+ sky130_fd_sc_hd__o211a_4
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _16371_/A _16371_/B _16371_/C _16371_/D vssd1 vssd1 vccd1 vccd1 _16428_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _19494_/Q _18906_/Q _18943_/Q _18517_/Q _10700_/S _11496_/A vssd1 vssd1 vccd1
+ vccd1 _10795_/X sky130_fd_sc_hd__mux4_1
X_13583_ _16364_/S _17152_/A vssd1 vssd1 vccd1 vccd1 _13583_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18110_ _18108_/Y _18109_/X _18110_/S vssd1 vssd1 vccd1 vccd1 _18110_/X sky130_fd_sc_hd__mux2_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_55_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15322_ _15322_/A vssd1 vssd1 vccd1 vccd1 _19170_/D sky130_fd_sc_hd__clkbuf_1
X_19090_ _19314_/CLK _19090_/D vssd1 vssd1 vccd1 vccd1 _19090_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12534_/A _12534_/B _12534_/C vssd1 vssd1 vccd1 vccd1 _12535_/B sky130_fd_sc_hd__nand3_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18041_ _12414_/Y _18007_/X _18040_/X _18028_/X vssd1 vssd1 vccd1 vccd1 _18041_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_145_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15253_ _15253_/A vssd1 vssd1 vccd1 vccd1 _19146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12465_ _19603_/Q _12465_/B vssd1 vssd1 vccd1 vccd1 _12511_/C sky130_fd_sc_hd__and2_1
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14204_ _14204_/A vssd1 vssd1 vccd1 vccd1 _18721_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11202__A _11202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ _11558_/B vssd1 vssd1 vccd1 vccd1 _11416_/Y sky130_fd_sc_hd__inv_2
X_15184_ _15184_/A vssd1 vssd1 vccd1 vccd1 _19123_/D sky130_fd_sc_hd__clkbuf_1
X_12396_ _19536_/Q _12120_/X _12314_/A vssd1 vssd1 vccd1 vccd1 _12396_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11454__S1 _10014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10567__C1 _10519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17495__A0 _12432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14135_ _14135_/A vssd1 vssd1 vccd1 vccd1 _18692_/D sky130_fd_sc_hd__clkbuf_1
X_11347_ _11302_/A _11301_/A _11324_/X _12631_/B vssd1 vssd1 vccd1 vccd1 _11582_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19992_ _20027_/CLK _19992_/D vssd1 vssd1 vccd1 vccd1 _19992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16204__S _16204_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14066_ _18663_/Q _13731_/X _14068_/S vssd1 vssd1 vccd1 vccd1 _14067_/A sky130_fd_sc_hd__mux2_1
X_18943_ _19366_/CLK _18943_/D vssd1 vssd1 vccd1 vccd1 _18943_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12859__A1 _16315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _19099_/Q _18865_/Q _19547_/Q _19195_/Q _10977_/A _10006_/A vssd1 vssd1 vccd1
+ vccd1 _11279_/B sky130_fd_sc_hd__mux4_1
XANTENNA_output78_A _12234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11206__S1 _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10229_ _10229_/A _10229_/B vssd1 vssd1 vccd1 vccd1 _10229_/Y sky130_fd_sc_hd__nor2_1
X_13017_ _14151_/B _18295_/A _14917_/D vssd1 vssd1 vccd1 vccd1 _13454_/A sky130_fd_sc_hd__and3b_4
X_18874_ _19430_/CLK _18874_/D vssd1 vssd1 vccd1 vccd1 _18874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17825_ _12003_/Y _17755_/X _17824_/X _17778_/X vssd1 vssd1 vccd1 vccd1 _17825_/X
+ sky130_fd_sc_hd__a211o_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17756_ _11907_/X _17755_/X _09464_/X vssd1 vssd1 vccd1 vccd1 _17756_/X sky130_fd_sc_hd__a21o_1
X_14968_ _19024_/Q _14443_/X _14972_/S vssd1 vssd1 vccd1 vccd1 _14969_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16707_ _16708_/B _17123_/B _19674_/Q vssd1 vssd1 vccd1 vccd1 _16709_/B sky130_fd_sc_hd__a21oi_1
X_13919_ _13919_/A vssd1 vssd1 vccd1 vccd1 _18598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17687_ _17685_/X _17686_/X _17760_/S vssd1 vssd1 vccd1 vccd1 _17687_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14899_ _14899_/A vssd1 vssd1 vccd1 vccd1 _18993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11390__S0 _10048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11083__S _11083_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19426_ _19552_/CLK _19426_/D vssd1 vssd1 vccd1 vccd1 _19426_/Q sky130_fd_sc_hd__dfxtp_1
X_16638_ _16672_/A _16638_/B _16638_/C vssd1 vssd1 vccd1 vccd1 _19653_/D sky130_fd_sc_hd__nor3_1
XFILLER_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13799__A _14624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19357_ _19726_/CLK _19357_/D vssd1 vssd1 vccd1 vccd1 _19357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16569_ _19630_/Q _16572_/C _16533_/X vssd1 vssd1 vccd1 vccd1 _16569_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11142__S0 _11224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11598__B2 _11534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18308_ _18308_/A _18331_/B vssd1 vssd1 vccd1 vccd1 _18308_/Y sky130_fd_sc_hd__nand2_1
X_19288_ _19288_/CLK _19288_/D vssd1 vssd1 vccd1 vccd1 _19288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10935__B _12643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15733__A0 _19905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18239_ _18239_/A vssd1 vssd1 vccd1 vccd1 _19974_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18390__A _18396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12208__A _14477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17486__A0 _17484_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15519__A _15587_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10951__A _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09943_ _09936_/Y _09938_/Y _09940_/Y _09942_/Y _09719_/A vssd1 vssd1 vccd1 vccd1
+ _09943_/X sky130_fd_sc_hd__o221a_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11258__S _11306_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _09887_/A vssd1 vssd1 vccd1 vccd1 _09874_/X sky130_fd_sc_hd__clkbuf_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09951__S _10826_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10956__S0 _10893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12878__A _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15254__A _15254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10089__A1 _10746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11038__B1 _09703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09877__S1 _09887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ _20044_/Q vssd1 vssd1 vccd1 vccd1 _18331_/A sky130_fd_sc_hd__clkinv_2
X_10580_ _19499_/Q _18911_/Q _18948_/Q _18522_/Q _10533_/S _09665_/A vssd1 vssd1 vccd1
+ vccd1 _10580_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_clock clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_139_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09239_ _20052_/Q _20027_/Q _20026_/Q _20025_/Q vssd1 vssd1 vccd1 vccd1 _09266_/B
+ sky130_fd_sc_hd__or4bb_2
XFILLER_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12250_ _18316_/A _12189_/A _12190_/X vssd1 vssd1 vccd1 vccd1 _12250_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11201_ _19358_/Q _18972_/Q _19422_/Q _18541_/Q _11306_/S _09511_/A vssd1 vssd1 vccd1
+ vccd1 _11202_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13648__S _13652_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12181_ _19528_/Q _11915_/A _12032_/A vssd1 vssd1 vccd1 vccd1 _12181_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11132_ _11315_/A _11132_/B vssd1 vssd1 vccd1 vccd1 _11132_/X sky130_fd_sc_hd__or2_1
X_11063_ _11001_/A _11057_/X _11061_/X _11127_/A vssd1 vssd1 vccd1 vccd1 _11063_/X
+ sky130_fd_sc_hd__a211o_1
X_15940_ _19397_/Q _15228_/X _15940_/S vssd1 vssd1 vccd1 vccd1 _15941_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10947__S0 _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09801__S1 _09730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _10014_/A vssd1 vssd1 vccd1 vccd1 _10014_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15871_ _13219_/X _19366_/Q _15879_/S vssd1 vssd1 vccd1 vccd1 _15872_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17610_ _17815_/A _17610_/B vssd1 vssd1 vccd1 vccd1 _17610_/X sky130_fd_sc_hd__or2_1
XANTENNA__16452__A1 _16449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__A _11704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14822_ _14822_/A vssd1 vssd1 vccd1 vccd1 _18963_/D sky130_fd_sc_hd__clkbuf_1
X_18590_ _19565_/CLK _18590_/D vssd1 vssd1 vccd1 vccd1 _18590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17541_ _12673_/A _12673_/B _17607_/A _17849_/A vssd1 vssd1 vccd1 vccd1 _17541_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14753_ _15918_/B _16134_/B vssd1 vssd1 vccd1 vccd1 _14810_/A sky130_fd_sc_hd__nor2_4
XFILLER_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11965_ _17792_/A _11965_/B vssd1 vssd1 vccd1 vccd1 _11968_/A sky130_fd_sc_hd__xor2_2
XANTENNA_output116_A _12653_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13704_ _13704_/A vssd1 vssd1 vccd1 vccd1 _18528_/D sky130_fd_sc_hd__clkbuf_1
X_10916_ _10978_/A vssd1 vssd1 vccd1 vccd1 _10917_/A sky130_fd_sc_hd__buf_2
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17472_ _17688_/A vssd1 vssd1 vccd1 vccd1 _17845_/A sky130_fd_sc_hd__clkbuf_2
X_14684_ _14684_/A vssd1 vssd1 vccd1 vccd1 _18896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11896_ _11961_/A _12637_/B _11962_/A _18336_/A vssd1 vssd1 vccd1 vccd1 _17749_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19211_ _19308_/CLK _19211_/D vssd1 vssd1 vccd1 vccd1 _19211_/Q sky130_fd_sc_hd__dfxtp_1
X_16423_ _16423_/A vssd1 vssd1 vccd1 vccd1 _19568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13635_ _13744_/S vssd1 vssd1 vccd1 vccd1 _13652_/S sky130_fd_sc_hd__buf_2
X_10847_ _18676_/Q _19171_/Q _10847_/S vssd1 vssd1 vccd1 vccd1 _10848_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15103__S _15105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11124__S0 _11004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13412__A _15270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19142_ _19272_/CLK _19142_/D vssd1 vssd1 vccd1 vccd1 _19142_/Q sky130_fd_sc_hd__dfxtp_1
X_16354_ _16361_/C _16353_/Y _16303_/X vssd1 vssd1 vccd1 vccd1 _16354_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ _11950_/B _18501_/Q _13598_/S vssd1 vssd1 vccd1 vccd1 _13567_/A sky130_fd_sc_hd__mux2_1
X_10778_ _10644_/X _10776_/Y _10777_/Y _10010_/X vssd1 vssd1 vccd1 vccd1 _10778_/X
+ sky130_fd_sc_hd__a211o_1
X_15305_ _15305_/A vssd1 vssd1 vccd1 vccd1 _19162_/D sky130_fd_sc_hd__clkbuf_1
X_12517_ _17234_/A _12545_/C vssd1 vssd1 vccd1 vccd1 _12517_/Y sky130_fd_sc_hd__nand2_1
X_19073_ _19200_/CLK _19073_/D vssd1 vssd1 vccd1 vccd1 _19073_/Q sky130_fd_sc_hd__dfxtp_1
X_16285_ _16285_/A _16285_/B vssd1 vssd1 vccd1 vccd1 _16285_/X sky130_fd_sc_hd__or2_1
X_13497_ _19878_/Q _12992_/X _12695_/A _19845_/Q vssd1 vssd1 vccd1 vccd1 _13497_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18024_ _17771_/X _18020_/Y _18023_/Y vssd1 vssd1 vccd1 vccd1 _18024_/Y sky130_fd_sc_hd__a21oi_1
X_15236_ _19141_/Q _15235_/X _15245_/S vssd1 vssd1 vccd1 vccd1 _15237_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ _19602_/Q _11771_/X _12447_/X vssd1 vssd1 vccd1 vccd1 _12448_/X sky130_fd_sc_hd__o21a_4
XFILLER_160_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13558__S _13558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15167_ _19115_/Q vssd1 vssd1 vccd1 vccd1 _15168_/A sky130_fd_sc_hd__clkbuf_1
X_12379_ _12473_/A _12660_/B _12474_/A _12378_/X vssd1 vssd1 vccd1 vccd1 _18023_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14118_ _18685_/Q _13689_/X _14120_/S vssd1 vssd1 vccd1 vccd1 _14119_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15098_ _15098_/A vssd1 vssd1 vccd1 vccd1 _19081_/D sky130_fd_sc_hd__clkbuf_1
X_19975_ _19978_/CLK _19975_/D vssd1 vssd1 vccd1 vccd1 _19975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10960__C1 _09601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14049_ _18655_/Q _13697_/X _14057_/S vssd1 vssd1 vccd1 vccd1 _14050_/A sky130_fd_sc_hd__mux2_1
X_18926_ _19514_/CLK _18926_/D vssd1 vssd1 vccd1 vccd1 _18926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11504__A1 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18857_ _19449_/CLK _18857_/D vssd1 vssd1 vccd1 vccd1 _18857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12698__A _12992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15074__A _15131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09590_ _19387_/Q _19001_/Q _19451_/Q _18570_/Q _09568_/X _09526_/A vssd1 vssd1 vccd1
+ vccd1 _09591_/B sky130_fd_sc_hd__mux4_1
X_17808_ _19900_/Q _17807_/X _17808_/S vssd1 vssd1 vccd1 vccd1 _17809_/A sky130_fd_sc_hd__mux2_1
X_18788_ _19443_/CLK _18788_/D vssd1 vssd1 vccd1 vccd1 _18788_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13257__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17739_ _17591_/X _17581_/X _17739_/S vssd1 vssd1 vccd1 vccd1 _17740_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18196__A1 _19988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__S0 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11107__A _19898_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17943__A1 _12204_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19409_ _19409_/CLK _19409_/D vssd1 vssd1 vccd1 vccd1 _19409_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16109__S _16117_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09859__S1 _09858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14852__S _14856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14153__A _14209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09926_ _18819_/Q _19154_/Q _09926_/S vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__mux2_1
XFILLER_132_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12299__A2 _12656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09795__S0 _09726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20046_ _20048_/CLK _20046_/D vssd1 vssd1 vccd1 vccd1 _20046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09857_ _10393_/A vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09788_/Y sky130_fd_sc_hd__nand2_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18295__A _18295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13931__S _13939_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11750_ _11745_/X _11740_/Y _11749_/X _16444_/C _19579_/Q vssd1 vssd1 vccd1 vccd1
+ _16447_/B sky130_fd_sc_hd__a32o_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17934__A1 _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10701_ _10701_/A vssd1 vssd1 vccd1 vccd1 _10701_/Y sky130_fd_sc_hd__inv_2
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16019__S _16023_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ _12602_/A _12596_/A vssd1 vssd1 vccd1 vccd1 _11681_/Y sky130_fd_sc_hd__nand2_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11451__S _11451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13420_ _13363_/A _13419_/X _13351_/X vssd1 vssd1 vccd1 vccd1 _13420_/Y sky130_fd_sc_hd__a21oi_2
X_10632_ _10632_/A _10632_/B vssd1 vssd1 vccd1 vccd1 _10632_/X sky130_fd_sc_hd__or2_1
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ _18778_/Q _19049_/Q _19273_/Q _19017_/Q _10382_/A _09815_/A vssd1 vssd1 vccd1
+ vccd1 _10563_/X sky130_fd_sc_hd__mux4_1
X_13351_ _13351_/A vssd1 vssd1 vccd1 vccd1 _13351_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14762__S _14764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12302_ _17989_/B _12302_/B vssd1 vssd1 vccd1 vccd1 _12332_/A sky130_fd_sc_hd__xnor2_1
XFILLER_5_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16070_ _16070_/A vssd1 vssd1 vccd1 vccd1 _19454_/D sky130_fd_sc_hd__clkbuf_1
X_10494_ _18684_/Q _19179_/Q _10494_/S vssd1 vssd1 vccd1 vccd1 _10495_/A sky130_fd_sc_hd__mux2_1
X_13282_ _13282_/A _13297_/C vssd1 vssd1 vccd1 vccd1 _13282_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15021_ _15021_/A vssd1 vssd1 vccd1 vccd1 _19047_/D sky130_fd_sc_hd__clkbuf_1
X_12233_ _12233_/A vssd1 vssd1 vccd1 vccd1 _12234_/B sky130_fd_sc_hd__clkinv_8
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10093__S0 _10081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ _17903_/B _12139_/B _12252_/A vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__a21o_1
XFILLER_151_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11115_ _11115_/A _11115_/B vssd1 vssd1 vccd1 vccd1 _11115_/X sky130_fd_sc_hd__and2_1
XFILLER_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19760_ _19762_/CLK _19760_/D vssd1 vssd1 vccd1 vccd1 _19760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16972_ _19749_/Q _19748_/Q _16972_/C vssd1 vssd1 vccd1 vccd1 _16978_/C sky130_fd_sc_hd__and3_1
X_12095_ _12095_/A _12095_/B vssd1 vssd1 vccd1 vccd1 _12096_/A sky130_fd_sc_hd__and2_4
XFILLER_150_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18711_ _19302_/CLK _18711_/D vssd1 vssd1 vccd1 vccd1 _18711_/Q sky130_fd_sc_hd__dfxtp_1
X_15923_ _19389_/Q _15203_/X _15929_/S vssd1 vssd1 vccd1 vccd1 _15924_/A sky130_fd_sc_hd__mux2_1
X_11046_ _11046_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11046_/Y sky130_fd_sc_hd__nor2_1
X_19691_ _19804_/CLK _19691_/D vssd1 vssd1 vccd1 vccd1 _19691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17622__B1 _09419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18642_ _19042_/CLK _18642_/D vssd1 vssd1 vccd1 vccd1 _18642_/Q sky130_fd_sc_hd__dfxtp_1
X_15854_ _15854_/A vssd1 vssd1 vccd1 vccd1 _19358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14805_ _14805_/A vssd1 vssd1 vccd1 vccd1 _18955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18573_ _19389_/CLK _18573_/D vssd1 vssd1 vccd1 vccd1 _18573_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12447__C1 _12494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15785_ _19914_/Q _15784_/X _15800_/S vssd1 vssd1 vccd1 vccd1 _15785_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12997_ _19610_/Q _12861_/X _12996_/X vssd1 vssd1 vccd1 vccd1 _12997_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14937__S _14939_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17524_ _17995_/A vssd1 vssd1 vccd1 vccd1 _17524_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14736_ _14736_/A vssd1 vssd1 vccd1 vccd1 _18920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11948_ _12420_/A vssd1 vssd1 vccd1 vccd1 _16226_/A sky130_fd_sc_hd__buf_2
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _17450_/X _17453_/X _17573_/S vssd1 vssd1 vccd1 vccd1 _17455_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14667_ _14666_/X _18892_/Q _14670_/S vssd1 vssd1 vccd1 vccd1 _14668_/A sky130_fd_sc_hd__mux2_1
X_11879_ _19882_/Q _09345_/X _13604_/A vssd1 vssd1 vccd1 vccd1 _11879_/Y sky130_fd_sc_hd__a21oi_1
X_16406_ _16428_/A vssd1 vssd1 vccd1 vccd1 _16415_/S sky130_fd_sc_hd__buf_2
X_13618_ _14580_/A vssd1 vssd1 vccd1 vccd1 _13618_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17386_ _17545_/B vssd1 vssd1 vccd1 vccd1 _17668_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14598_ _14598_/A vssd1 vssd1 vccd1 vccd1 _18870_/D sky130_fd_sc_hd__clkbuf_1
X_19125_ _19401_/CLK _19125_/D vssd1 vssd1 vccd1 vccd1 _19125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16337_ _19950_/Q _16338_/B vssd1 vssd1 vccd1 vccd1 _16347_/C sky130_fd_sc_hd__or2_2
X_13549_ _19769_/Q _12991_/X _13548_/X _12995_/X vssd1 vssd1 vccd1 vccd1 _13549_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16453__A _18404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19056_ _19411_/CLK _19056_/D vssd1 vssd1 vccd1 vccd1 _19056_/Q sky130_fd_sc_hd__dfxtp_1
X_16268_ _16268_/A vssd1 vssd1 vccd1 vccd1 _16318_/S sky130_fd_sc_hd__buf_2
XFILLER_145_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18007_ _18007_/A vssd1 vssd1 vccd1 vccd1 _18007_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15219_ _15219_/A vssd1 vssd1 vccd1 vccd1 _15219_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16199_ _16199_/A vssd1 vssd1 vccd1 vccd1 _19512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11186__C1 _10994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16900__B _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10006__A _10006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19958_ _20000_/CLK _19958_/D vssd1 vssd1 vccd1 vccd1 _19958_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13478__B2 _19541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_177_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ _09711_/A vssd1 vssd1 vccd1 vccd1 _09712_/A sky130_fd_sc_hd__clkbuf_2
X_18909_ _19497_/CLK _18909_/D vssd1 vssd1 vccd1 vccd1 _18909_/Q sky130_fd_sc_hd__dfxtp_1
X_19889_ _19892_/CLK _19889_/D vssd1 vssd1 vccd1 vccd1 _19889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09642_ _11222_/S vssd1 vssd1 vccd1 vccd1 _10968_/S sky130_fd_sc_hd__buf_4
XFILLER_67_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09573_ _18968_/Q vssd1 vssd1 vccd1 vccd1 _09574_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16347__B _16347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09530__A _09530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14148__A _14148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10075__S0 _10073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13926__S _13926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17194__A _17194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13469__A1 _13054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09909_ _18787_/Q _19058_/Q _19282_/Q _19026_/Q _10244_/S _10148_/A vssd1 vssd1 vccd1
+ vccd1 _09909_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09768__S0 _09761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12141__A1 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ _19730_/Q _13144_/S _12723_/A _19698_/Q _12919_/X vssd1 vssd1 vccd1 vccd1
+ _12920_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20029_ _20032_/CLK _20029_/D vssd1 vssd1 vccd1 vccd1 _20029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _18448_/Q _12851_/B vssd1 vssd1 vccd1 vccd1 _12851_/X sky130_fd_sc_hd__or2_1
XFILLER_62_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13661__S _13673_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _20044_/Q _18319_/A _11853_/S vssd1 vssd1 vccd1 vccd1 _11802_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15570_ _19281_/Q _15273_/X _15572_/S vssd1 vssd1 vccd1 vccd1 _15571_/A sky130_fd_sc_hd__mux2_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _19868_/Q _12755_/A _12758_/A _19532_/Q _12781_/X vssd1 vssd1 vccd1 vccd1
+ _12782_/X sky130_fd_sc_hd__a221o_1
XFILLER_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09440__A _20044_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14521_/A vssd1 vssd1 vccd1 vccd1 _18839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _11733_/A _11733_/B _11733_/C vssd1 vssd1 vccd1 vccd1 _12097_/A sky130_fd_sc_hd__or3_4
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _17240_/A _17240_/B vssd1 vssd1 vccd1 vccd1 _17240_/X sky130_fd_sc_hd__or2_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14452_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11664_ _17338_/B _18328_/A _12207_/C _12207_/D vssd1 vssd1 vccd1 vccd1 _11749_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_30_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13403_ _19346_/Q _12759_/X _12704_/X _19536_/Q _13402_/X vssd1 vssd1 vccd1 vccd1
+ _13403_/X sky130_fd_sc_hd__a221o_1
X_10615_ _10691_/A vssd1 vssd1 vccd1 vccd1 _11371_/A sky130_fd_sc_hd__buf_4
X_17171_ _17185_/A vssd1 vssd1 vccd1 vccd1 _17171_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14383_ _18798_/Q _14382_/X _14386_/S vssd1 vssd1 vccd1 vccd1 _14384_/A sky130_fd_sc_hd__mux2_1
X_11595_ _10146_/A _11546_/X _11547_/X _11548_/Y _11594_/X vssd1 vssd1 vccd1 vccd1
+ _11595_/X sky130_fd_sc_hd__a221o_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16122_ _13471_/X _19478_/Q _16128_/S vssd1 vssd1 vccd1 vccd1 _16123_/A sky130_fd_sc_hd__mux2_1
X_13334_ _16301_/B _13335_/C _19944_/Q vssd1 vssd1 vccd1 vccd1 _13336_/B sky130_fd_sc_hd__a21oi_1
X_10546_ _10583_/A _10545_/X _09695_/A vssd1 vssd1 vccd1 vccd1 _10546_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_3_4_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_157_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16053_ _16053_/A vssd1 vssd1 vccd1 vccd1 _19447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13265_ _19338_/Q _12707_/X _12704_/A _19528_/Q _13264_/X vssd1 vssd1 vccd1 vccd1
+ _13265_/X sky130_fd_sc_hd__a221o_1
XFILLER_157_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10477_ _19501_/Q _18913_/Q _18950_/Q _18524_/Q _10382_/X _10462_/X vssd1 vssd1 vccd1
+ vccd1 _10478_/B sky130_fd_sc_hd__mux4_1
XFILLER_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15004_ _15004_/A vssd1 vssd1 vccd1 vccd1 _19039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12216_ _17192_/A _12217_/C _19832_/Q vssd1 vssd1 vccd1 vccd1 _12216_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09318__C _20042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13196_ _18478_/Q _13195_/X _13196_/S vssd1 vssd1 vccd1 vccd1 _13197_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13836__S _13845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19812_ _20044_/CLK _19812_/D vssd1 vssd1 vccd1 vccd1 _19812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ _12147_/A _12147_/B vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__xnor2_2
XFILLER_151_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09615__A _09615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19743_ _19745_/CLK _19743_/D vssd1 vssd1 vccd1 vccd1 _19743_/Q sky130_fd_sc_hd__dfxtp_1
X_16955_ _16955_/A _16955_/B _16955_/C vssd1 vssd1 vccd1 vccd1 _16971_/C sky130_fd_sc_hd__and3_1
X_12078_ _12080_/A _12080_/B vssd1 vssd1 vccd1 vccd1 _12079_/A sky130_fd_sc_hd__or2_1
XANTENNA__12132__A1 _12127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18399__B2 _18398_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15906_ _13471_/X _19382_/Q _15912_/S vssd1 vssd1 vccd1 vccd1 _15907_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17832__A _17832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ _11327_/S vssd1 vssd1 vccd1 vccd1 _11030_/A sky130_fd_sc_hd__clkbuf_4
X_19674_ _19805_/CLK _19674_/D vssd1 vssd1 vccd1 vccd1 _19674_/Q sky130_fd_sc_hd__dfxtp_1
X_16886_ _16922_/B _16891_/D _16885_/X vssd1 vssd1 vccd1 vccd1 _19726_/D sky130_fd_sc_hd__o21ba_1
XFILLER_38_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18625_ _19411_/CLK _18625_/D vssd1 vssd1 vccd1 vccd1 _18625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15837_ _15837_/A _18467_/Q vssd1 vssd1 vccd1 vccd1 _15837_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14667__S _14670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12976__A _12976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18556_ _19563_/CLK _18556_/D vssd1 vssd1 vccd1 vccd1 _18556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15768_ _18456_/Q _15768_/B vssd1 vssd1 vccd1 vccd1 _15768_/X sky130_fd_sc_hd__or2_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14719_ _14719_/A vssd1 vssd1 vccd1 vccd1 _18912_/D sky130_fd_sc_hd__clkbuf_1
X_17507_ _12553_/A _17642_/B _17507_/S vssd1 vssd1 vccd1 vccd1 _17507_/X sky130_fd_sc_hd__mux2_1
X_18487_ _19470_/CLK _18487_/D vssd1 vssd1 vccd1 vccd1 _18487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15699_ _15699_/A vssd1 vssd1 vccd1 vccd1 _19330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17438_ _17677_/S vssd1 vssd1 vccd1 vccd1 _17802_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17369_ _11673_/A _18301_/A _17358_/X _19890_/Q vssd1 vssd1 vccd1 vccd1 _17370_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11946__A1 _19520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19108_ _19556_/CLK _19108_/D vssd1 vssd1 vccd1 vccd1 _19108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039_ _19487_/CLK _19039_/D vssd1 vssd1 vccd1 vccd1 _19039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput100 _11972_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[7] sky130_fd_sc_hd__buf_2
Xoutput111 _12647_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[11] sky130_fd_sc_hd__buf_2
Xoutput122 _12659_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[21] sky130_fd_sc_hd__buf_2
Xoutput133 _12671_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[31] sky130_fd_sc_hd__buf_2
XFILLER_161_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput144 _12096_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[11] sky130_fd_sc_hd__buf_2
XFILLER_161_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput155 _12375_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[21] sky130_fd_sc_hd__buf_2
XANTENNA__09228__C _09238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput166 _12629_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[31] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_opt_6_0_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16122__S _16128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09625_ _18829_/Q vssd1 vssd1 vccd1 vccd1 _11096_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12886__A _13527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__S0 _11129_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09556_ _11016_/A vssd1 vssd1 vccd1 vccd1 _10606_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09922__S0 _10173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09487_ _10574_/A vssd1 vssd1 vccd1 vccd1 _10569_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15201__S _15213_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10400_ _10407_/A _10395_/X _10399_/X vssd1 vssd1 vccd1 vccd1 _10400_/Y sky130_fd_sc_hd__o21ai_1
X_11380_ _10834_/A _11375_/X _11379_/X _09612_/A vssd1 vssd1 vccd1 vccd1 _11380_/Y
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__11949__B _11950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13139__B1 _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ _10396_/A vssd1 vssd1 vccd1 vccd1 _10332_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16821__A _17073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12126__A _16226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11030__A _11030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10262_ _09616_/A _10252_/X _10261_/X _09623_/A _19914_/Q vssd1 vssd1 vccd1 vccd1
+ _11418_/A sky130_fd_sc_hd__a32o_2
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13050_ _19895_/Q _13588_/B _13371_/A vssd1 vssd1 vccd1 vccd1 _13051_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ _11938_/A _11936_/A _11971_/A _12000_/X vssd1 vssd1 vccd1 vccd1 _12002_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_121_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11965__A _17792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16032__S _16034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ _09750_/X _10182_/X _10191_/X _09757_/X _10192_/Y vssd1 vssd1 vccd1 vccd1
+ _12661_/B sky130_fd_sc_hd__o32a_4
XFILLER_132_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15871__S _15879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16740_ _19684_/Q _19683_/Q _19682_/Q _16740_/D vssd1 vssd1 vccd1 vccd1 _16749_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_59_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13952_ _13998_/S vssd1 vssd1 vccd1 vccd1 _13961_/S sky130_fd_sc_hd__buf_2
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _12903_/A vssd1 vssd1 vccd1 vccd1 _12903_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_74_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16671_ _16670_/B _16670_/C _19665_/Q vssd1 vssd1 vccd1 vccd1 _16672_/C sky130_fd_sc_hd__a21oi_1
XFILLER_47_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13883_ _13787_/X _18582_/Q _13889_/S vssd1 vssd1 vccd1 vccd1 _13884_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16268__A _16268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15622_ _14621_/X _19304_/Q _15622_/S vssd1 vssd1 vccd1 vccd1 _15623_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18410_ _18412_/A _18410_/B vssd1 vssd1 vccd1 vccd1 _20043_/D sky130_fd_sc_hd__nor2_1
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12834_ _19717_/Q vssd1 vssd1 vccd1 vccd1 _16868_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_19390_ _19392_/CLK _19390_/D vssd1 vssd1 vccd1 vccd1 _19390_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _18341_/A vssd1 vssd1 vccd1 vccd1 _18341_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _19273_/Q _15247_/X _15561_/S vssd1 vssd1 vccd1 vccd1 _15554_/A sky130_fd_sc_hd__mux2_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12765_ _18454_/Q _13316_/B _13316_/C _12764_/Y vssd1 vssd1 vccd1 vccd1 _12765_/X
+ sky130_fd_sc_hd__or4b_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14572_/S vssd1 vssd1 vccd1 vccd1 _14513_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_125_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18272_ _18272_/A vssd1 vssd1 vccd1 vccd1 _19989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11764_/A _11764_/B _17610_/B vssd1 vssd1 vccd1 vccd1 _11717_/B sky130_fd_sc_hd__or3_1
X_15484_ _15484_/A vssd1 vssd1 vccd1 vccd1 _19242_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12696_/A vssd1 vssd1 vccd1 vccd1 _12696_/X sky130_fd_sc_hd__buf_2
XFILLER_42_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17223_ _17223_/A _17226_/B vssd1 vssd1 vccd1 vccd1 _17223_/X sky130_fd_sc_hd__or2_1
XFILLER_174_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14435_ _14435_/A vssd1 vssd1 vccd1 vccd1 _18814_/D sky130_fd_sc_hd__clkbuf_1
X_11647_ _11697_/B vssd1 vssd1 vccd1 vccd1 _12670_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 io_dbus_rdata[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_4
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput24 io_dbus_rdata[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_4
XFILLER_174_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17154_ _19818_/Q _17164_/B vssd1 vssd1 vccd1 vccd1 _17154_/X sky130_fd_sc_hd__or2_1
XFILLER_167_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput35 io_ibus_inst[10] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11859__B _17418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14366_ _14366_/A vssd1 vssd1 vccd1 vccd1 _18793_/D sky130_fd_sc_hd__clkbuf_1
Xinput46 io_ibus_inst[20] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
X_11578_ _11578_/A _11578_/B vssd1 vssd1 vccd1 vccd1 _11578_/Y sky130_fd_sc_hd__nand2_1
Xinput57 io_ibus_inst[30] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
X_16105_ _16105_/A vssd1 vssd1 vccd1 vccd1 _19470_/D sky130_fd_sc_hd__clkbuf_1
Xinput68 io_irq_spi_irq vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10600__A1 _09749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13317_ _13534_/S _19910_/Q _13337_/A _13316_/X vssd1 vssd1 vccd1 vccd1 _13317_/X
+ sky130_fd_sc_hd__o211a_1
X_10529_ _09615_/A _10519_/X _10528_/X _09622_/A _19909_/Q vssd1 vssd1 vccd1 vccd1
+ _10555_/A sky130_fd_sc_hd__a32o_4
X_17085_ _17087_/B _17087_/C _17059_/X vssd1 vssd1 vccd1 vccd1 _17085_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14297_ _16134_/A _15517_/B vssd1 vssd1 vccd1 vccd1 _14354_/A sky130_fd_sc_hd__nor2_4
XFILLER_6_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16036_ _16047_/A vssd1 vssd1 vccd1 vccd1 _16045_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13248_ _19751_/Q _12692_/A _13247_/X _12714_/A vssd1 vssd1 vccd1 vccd1 _13248_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15347__A _15358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13179_ _18477_/Q _13178_/X _13196_/S vssd1 vssd1 vccd1 vccd1 _13180_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09345__A _19894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17987_ _18078_/S _17988_/B _17986_/X _17723_/A vssd1 vssd1 vccd1 vccd1 _17990_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13302__B1 _13418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19726_ _19726_/CLK _19726_/D vssd1 vssd1 vccd1 vccd1 _19726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16938_ _16957_/C _16959_/B _16964_/A vssd1 vssd1 vccd1 vccd1 _16939_/C sky130_fd_sc_hd__nand3_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10211__S0 _10195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19657_ _19792_/CLK _19657_/D vssd1 vssd1 vccd1 vccd1 _19657_/Q sky130_fd_sc_hd__dfxtp_1
X_16869_ _16920_/B _16873_/D _19721_/Q vssd1 vssd1 vccd1 vccd1 _16871_/B sky130_fd_sc_hd__a21oi_1
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09410_ _09407_/X _11837_/A _09409_/X _19806_/Q vssd1 vssd1 vccd1 vccd1 _11774_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18608_ _19491_/CLK _18608_/D vssd1 vssd1 vccd1 vccd1 _18608_/Q sky130_fd_sc_hd__dfxtp_1
X_19588_ _19963_/CLK _19588_/D vssd1 vssd1 vccd1 vccd1 _19588_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10419__A1 _09899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ _19893_/Q vssd1 vssd1 vccd1 vccd1 _09341_/X sky130_fd_sc_hd__buf_4
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18539_ _19734_/CLK _18539_/D vssd1 vssd1 vccd1 vccd1 _18539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18393__A _18396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11115__A _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09272_ _09272_/A _09272_/B _09272_/C vssd1 vssd1 vccd1 vccd1 _17331_/B sky130_fd_sc_hd__or3_4
XFILLER_166_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16117__S _16117_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10278__S0 _09926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15956__S _15962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16641__A _16674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15257__A _15257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16491__C1 _12749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15833__A2 _18466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10202__S0 _09902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09608_ _09608_/A _11640_/A vssd1 vssd1 vccd1 vccd1 _09609_/B sky130_fd_sc_hd__nor2_4
XFILLER_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10880_ _10880_/A vssd1 vssd1 vccd1 vccd1 _11260_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ _10195_/S vssd1 vssd1 vccd1 vccd1 _10162_/S sky130_fd_sc_hd__buf_2
XFILLER_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _17538_/A _18090_/A _12527_/B vssd1 vssd1 vccd1 vccd1 _12551_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11501_ _18793_/Q _19064_/Q _19288_/Q _19032_/Q _10040_/A _10041_/A vssd1 vssd1 vccd1
+ vccd1 _11501_/X sky130_fd_sc_hd__mux4_1
X_12481_ _12481_/A _18068_/B vssd1 vssd1 vccd1 vccd1 _12520_/A sky130_fd_sc_hd__xor2_4
X_14220_ _13847_/X _18729_/Q _14222_/S vssd1 vssd1 vccd1 vccd1 _14221_/A sky130_fd_sc_hd__mux2_1
X_11432_ _18792_/Q _19063_/Q _19287_/Q _19031_/Q _10625_/X _10604_/A vssd1 vssd1 vccd1
+ vccd1 _11432_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14151_ _16371_/A _14151_/B _16371_/C vssd1 vssd1 vccd1 vccd1 _16062_/B sky130_fd_sc_hd__or3_1
XFILLER_138_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11363_ _19497_/Q _18909_/Q _18946_/Q _18520_/Q _10675_/X _09957_/X vssd1 vssd1 vccd1
+ vccd1 _11363_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ _16958_/A _12991_/X _13101_/X _12995_/X vssd1 vssd1 vccd1 vccd1 _13102_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10314_ _10314_/A vssd1 vssd1 vccd1 vccd1 _10314_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14082_ _14082_/A vssd1 vssd1 vccd1 vccd1 _18668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11294_ _19453_/Q _19291_/Q _18700_/Q _18470_/Q _11329_/S _11283_/A vssd1 vssd1 vccd1
+ vccd1 _11295_/B sky130_fd_sc_hd__mux4_1
XFILLER_3_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13033_ _15203_/A vssd1 vssd1 vccd1 vccd1 _13033_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17910_ _12148_/A _17966_/B _17905_/X _17909_/Y _11657_/S vssd1 vssd1 vccd1 vccd1
+ _17910_/X sky130_fd_sc_hd__o221a_2
XFILLER_98_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10245_ _18688_/Q _19183_/Q _10245_/S vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18890_ _19572_/CLK _18890_/D vssd1 vssd1 vccd1 vccd1 _18890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10176_ _10176_/A _10176_/B vssd1 vssd1 vccd1 vccd1 _10176_/Y sky130_fd_sc_hd__nand2_1
X_17841_ _18127_/A vssd1 vssd1 vccd1 vccd1 _18085_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_51_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10992__S1 _10974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14984_ _14984_/A vssd1 vssd1 vccd1 vccd1 _19031_/D sky130_fd_sc_hd__clkbuf_1
X_17772_ _17772_/A _17772_/B vssd1 vssd1 vccd1 vccd1 _17772_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18223__A0 _19967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19511_ _19511_/CLK _19511_/D vssd1 vssd1 vccd1 vccd1 _19511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16723_ _16860_/A vssd1 vssd1 vccd1 vccd1 _16723_/X sky130_fd_sc_hd__clkbuf_2
X_13935_ _18605_/Q _13622_/X _13939_/S vssd1 vssd1 vccd1 vccd1 _13936_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19442_ _19508_/CLK _19442_/D vssd1 vssd1 vccd1 vccd1 _19442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16654_ _16653_/B _16653_/C _19659_/Q vssd1 vssd1 vccd1 vccd1 _16655_/C sky130_fd_sc_hd__a21oi_1
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13866_ _13866_/A vssd1 vssd1 vccd1 vccd1 _18574_/D sky130_fd_sc_hd__clkbuf_1
X_15605_ _14596_/X _19296_/Q _15611_/S vssd1 vssd1 vccd1 vccd1 _15606_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12817_ _18440_/Q _12814_/Y _12816_/X vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__o21a_4
X_19373_ _19470_/CLK _19373_/D vssd1 vssd1 vccd1 vccd1 _19373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16585_ _16593_/A _16590_/C vssd1 vssd1 vccd1 vccd1 _16585_/Y sky130_fd_sc_hd__nor2_1
X_13797_ _13796_/X _18553_/Q _13797_/S vssd1 vssd1 vccd1 vccd1 _13798_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13063__A2 _16219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18324_ _18324_/A _18331_/B vssd1 vssd1 vccd1 vccd1 _18324_/Y sky130_fd_sc_hd__nand2_1
X_15536_ _15536_/A vssd1 vssd1 vccd1 vccd1 _19265_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _17319_/A vssd1 vssd1 vccd1 vccd1 _16939_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18255_ _18255_/A vssd1 vssd1 vccd1 vccd1 _18264_/S sky130_fd_sc_hd__clkbuf_2
X_15467_ _19235_/Q _15228_/X _15467_/S vssd1 vssd1 vccd1 vccd1 _15468_/A sky130_fd_sc_hd__mux2_1
X_12679_ _12893_/B _17140_/C _17149_/A vssd1 vssd1 vccd1 vccd1 _17247_/D sky130_fd_sc_hd__or3_2
XANTENNA__10774__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17206_ _15764_/Y _17197_/X _17205_/X _17201_/X vssd1 vssd1 vccd1 vccd1 _19835_/D
+ sky130_fd_sc_hd__o211a_1
X_14418_ _18809_/Q _14417_/X _14418_/S vssd1 vssd1 vccd1 vccd1 _14419_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18186_ _16347_/A _19983_/Q _18192_/S vssd1 vssd1 vccd1 vccd1 _18187_/A sky130_fd_sc_hd__mux2_1
X_15398_ _14608_/X _19204_/Q _15406_/S vssd1 vssd1 vccd1 vccd1 _15399_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17137_ _19813_/Q _12880_/X _17136_/X _16480_/X vssd1 vssd1 vccd1 vccd1 _19813_/D
+ sky130_fd_sc_hd__o211a_1
X_14349_ _14349_/A vssd1 vssd1 vccd1 vccd1 _18785_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17557__A _18127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16461__A _18404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17068_ _17070_/B _17070_/C _17059_/X vssd1 vssd1 vccd1 vccd1 _17068_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_144_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16019_ _13239_/X _19432_/Q _16023_/S vssd1 vssd1 vccd1 vccd1 _16020_/A sky130_fd_sc_hd__mux2_1
X_09890_ _18660_/Q _19251_/Q _19413_/Q _18628_/Q _09872_/X _09858_/X vssd1 vssd1 vccd1
+ vccd1 _09890_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16400__S _16404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10014__A _10014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18214__A0 _19963_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19709_ _19769_/CLK _19709_/D vssd1 vssd1 vccd1 vccd1 _19709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09324_ _19886_/Q _15819_/B vssd1 vssd1 vccd1 vccd1 _09339_/B sky130_fd_sc_hd__or2_1
XANTENNA__10499__S0 _10392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09255_ _09272_/B vssd1 vssd1 vccd1 vccd1 _11678_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09186_ _20033_/Q vssd1 vssd1 vccd1 vccd1 _09272_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__15751__A1 _18452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_162_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19794_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12565__A1 _19846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14590__S _14590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13514__B1 _13205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_177_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19844_/CLK sky130_fd_sc_hd__clkbuf_16
X_10030_ _10030_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10030_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17914__B _17914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14842__A1_N _18321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_3_0_clock clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_100_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19556_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__18205__A0 _19959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ _11951_/A _11980_/Y _19824_/Q _11776_/A vssd1 vssd1 vccd1 vccd1 _12034_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13720_ _18532_/Q _13718_/X _13736_/S vssd1 vssd1 vccd1 vccd1 _13721_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10932_ _10925_/Y _10927_/Y _10929_/Y _10931_/Y _10063_/A vssd1 vssd1 vccd1 vccd1
+ _10932_/X sky130_fd_sc_hd__o221a_1
XFILLER_90_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13651_ _14605_/A vssd1 vssd1 vccd1 vccd1 _13651_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10863_ _19461_/Q _19299_/Q _18708_/Q _18478_/Q _10702_/S _09662_/A vssd1 vssd1 vccd1
+ vccd1 _10863_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_115_clock clkbuf_opt_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19954_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ _12602_/A vssd1 vssd1 vccd1 vccd1 _18308_/A sky130_fd_sc_hd__clkinv_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _16370_/A vssd1 vssd1 vccd1 vccd1 _19545_/D sky130_fd_sc_hd__clkbuf_1
X_13582_ _18438_/Q _13577_/X _13581_/X vssd1 vssd1 vccd1 vccd1 _17152_/A sky130_fd_sc_hd__a21oi_4
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _10794_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _10794_/Y sky130_fd_sc_hd__nor2_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _19170_/Q _15225_/X _15323_/S vssd1 vssd1 vccd1 vccd1 _15322_/A sky130_fd_sc_hd__mux2_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _12534_/A _12534_/B _12534_/C vssd1 vssd1 vccd1 vccd1 _12535_/A sky130_fd_sc_hd__a21o_2
XANTENNA__10803__A1 _10746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18040_ _17928_/X _17812_/X _18039_/X _17953_/X vssd1 vssd1 vccd1 vccd1 _18040_/X
+ sky130_fd_sc_hd__o211a_1
X_15252_ _19146_/Q _15251_/X _15261_/S vssd1 vssd1 vccd1 vccd1 _15253_/A sky130_fd_sc_hd__mux2_1
X_12464_ _19603_/Q _12465_/B vssd1 vssd1 vccd1 vccd1 _12466_/A sky130_fd_sc_hd__nor2_1
XFILLER_173_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14203_ _13822_/X _18721_/Q _14207_/S vssd1 vssd1 vccd1 vccd1 _14204_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15596__S _15600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11415_ _11415_/A _12656_/B vssd1 vssd1 vccd1 vccd1 _11558_/B sky130_fd_sc_hd__nand2_1
X_15183_ _19123_/Q vssd1 vssd1 vccd1 vccd1 _15184_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_138_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12395_ _12391_/Y _12394_/Y _12395_/S vssd1 vssd1 vccd1 vccd1 _12395_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14134_ _18692_/Q _13718_/X _14142_/S vssd1 vssd1 vccd1 vccd1 _14135_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17495__A1 _17792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11346_ _09745_/A _11336_/X _11345_/X _09752_/A _09342_/Y vssd1 vssd1 vccd1 vccd1
+ _12631_/B sky130_fd_sc_hd__o32a_4
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19991_ _20027_/CLK _19991_/D vssd1 vssd1 vccd1 vccd1 _19991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14065_ _14065_/A vssd1 vssd1 vccd1 vccd1 _18662_/D sky130_fd_sc_hd__clkbuf_1
X_18942_ _19204_/CLK _18942_/D vssd1 vssd1 vccd1 vccd1 _18942_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10319__B1 _09826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14005__S _14013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11277_ _09610_/A _11267_/X _11276_/X _09618_/A _19894_/Q vssd1 vssd1 vccd1 vccd1
+ _11302_/A sky130_fd_sc_hd__a32o_4
XANTENNA__12859__A2 _12854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13016_ _14148_/A _14501_/B _14000_/B vssd1 vssd1 vccd1 vccd1 _14917_/D sky130_fd_sc_hd__and3_1
XANTENNA__10414__S0 _10367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ _19378_/Q _18992_/Q _19442_/Q _18561_/Q _09872_/X _09874_/X vssd1 vssd1 vccd1
+ vccd1 _10229_/B sky130_fd_sc_hd__mux4_1
X_18873_ _19203_/CLK _18873_/D vssd1 vssd1 vccd1 vccd1 _18873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17824_ _17521_/X _17811_/X _17823_/X _17776_/X vssd1 vssd1 vccd1 vccd1 _17824_/X
+ sky130_fd_sc_hd__o211a_1
X_10159_ _19121_/Q _18887_/Q _19569_/Q _19217_/Q _09508_/A _10148_/X vssd1 vssd1 vccd1
+ vccd1 _10159_/X sky130_fd_sc_hd__mux4_2
XANTENNA__13269__C1 _13268_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14967_ _14967_/A vssd1 vssd1 vccd1 vccd1 _19023_/D sky130_fd_sc_hd__clkbuf_1
X_17755_ _17755_/A vssd1 vssd1 vccd1 vccd1 _17755_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16706_ _16710_/D vssd1 vssd1 vccd1 vccd1 _17123_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13918_ _13838_/X _18598_/Q _13922_/S vssd1 vssd1 vccd1 vccd1 _13919_/A sky130_fd_sc_hd__mux2_1
X_14898_ _14650_/X _18993_/Q _14900_/S vssd1 vssd1 vccd1 vccd1 _14899_/A sky130_fd_sc_hd__mux2_1
X_17686_ _17568_/X _17582_/X _17686_/S vssd1 vssd1 vccd1 vccd1 _17686_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11390__S1 _10037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19425_ _19551_/CLK _19425_/D vssd1 vssd1 vccd1 vccd1 _19425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16637_ _16636_/B _16636_/C _19653_/Q vssd1 vssd1 vccd1 vccd1 _16638_/C sky130_fd_sc_hd__a21oi_1
X_13849_ _13849_/A vssd1 vssd1 vccd1 vccd1 _18569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17970__A2 _17861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19356_ _19726_/CLK _19356_/D vssd1 vssd1 vccd1 vccd1 _19356_/Q sky130_fd_sc_hd__dfxtp_1
X_16568_ _19629_/Q _16566_/B _16567_/Y vssd1 vssd1 vccd1 vccd1 _19629_/D sky130_fd_sc_hd__o21a_1
X_18307_ _20002_/Q _18285_/X _18306_/Y _18303_/X vssd1 vssd1 vccd1 vccd1 _20002_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11142__S1 _11330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15519_ _15587_/S vssd1 vssd1 vccd1 vccd1 _15528_/S sky130_fd_sc_hd__buf_2
X_19287_ _19287_/CLK _19287_/D vssd1 vssd1 vccd1 vccd1 _19287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16499_ _19655_/Q _19657_/Q _19656_/Q _16640_/A vssd1 vssd1 vccd1 vccd1 _16648_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__15733__A1 _12874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18238_ _19974_/Q _12263_/A _18242_/S vssd1 vssd1 vccd1 vccd1 _18239_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12547__A1 _19606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16191__A _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18169_ _18169_/A vssd1 vssd1 vccd1 vccd1 _19943_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14704__A _14750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__A _10910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_94_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19401_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09942_ _10279_/A _09941_/X _09711_/A vssd1 vssd1 vccd1 vccd1 _09942_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09873_ _10393_/A vssd1 vssd1 vccd1 vccd1 _09887_/A sky130_fd_sc_hd__clkbuf_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10956__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16130__S _16132_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09533__A _10811_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_32_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19306_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15270__A _15270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11038__A1 _11141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09307_ _11523_/A _09307_/B _09467_/B _11682_/B vssd1 vssd1 vccd1 vccd1 _12611_/A
+ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_47_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19377_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09238_ _09238_/A _11730_/C vssd1 vssd1 vccd1 vccd1 _09244_/A sky130_fd_sc_hd__or2_1
XFILLER_166_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17197__A _17197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11200_ _11259_/S vssd1 vssd1 vccd1 vccd1 _11306_/S sky130_fd_sc_hd__buf_4
XFILLER_163_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12180_ _12153_/A _12153_/B _12179_/Y _11977_/A vssd1 vssd1 vccd1 vccd1 _12180_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11449__S _11449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11131_ _18639_/Q _19230_/Q _19392_/Q _18607_/Q _11003_/A _11059_/A vssd1 vssd1 vccd1
+ vccd1 _11132_/B sky130_fd_sc_hd__mux4_1
XFILLER_122_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11062_ _11315_/A vssd1 vssd1 vccd1 vccd1 _11127_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10013_ _10105_/A vssd1 vssd1 vccd1 vccd1 _10014_/A sky130_fd_sc_hd__buf_4
XFILLER_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10947__S1 _09511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15870_ _15916_/S vssd1 vssd1 vccd1 vccd1 _15879_/S sky130_fd_sc_hd__buf_6
XFILLER_48_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12788__B _18455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14821_ _18963_/Q _14468_/X _14823_/S vssd1 vssd1 vccd1 vccd1 _14822_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input22_A io_dbus_rdata[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14752_ _14828_/A _14752_/B vssd1 vssd1 vccd1 vccd1 _18932_/D sky130_fd_sc_hd__nor2_1
X_17540_ _18118_/A vssd1 vssd1 vccd1 vccd1 _17849_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11277__B2 _19894_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ _11990_/A _11926_/A _11990_/C _11928_/A vssd1 vssd1 vccd1 vccd1 _11965_/B
+ sky130_fd_sc_hd__o31a_1
X_13703_ _18528_/Q _13702_/X _13715_/S vssd1 vssd1 vccd1 vccd1 _13704_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10915_ _18828_/Q vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__buf_2
X_17471_ _17662_/A vssd1 vssd1 vccd1 vccd1 _17688_/A sky130_fd_sc_hd__clkbuf_2
X_14683_ _18896_/Q _14369_/X _14691_/S vssd1 vssd1 vccd1 vccd1 _14684_/A sky130_fd_sc_hd__mux2_1
X_11895_ _12320_/B _17327_/B _11895_/C vssd1 vssd1 vccd1 vccd1 _11962_/A sky130_fd_sc_hd__and3_1
XANTENNA_output109_A _12631_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19210_ _19306_/CLK _19210_/D vssd1 vssd1 vccd1 vccd1 _19210_/Q sky130_fd_sc_hd__dfxtp_1
X_16422_ _13412_/X _19568_/Q _16426_/S vssd1 vssd1 vccd1 vccd1 _16423_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13634_ _14592_/A vssd1 vssd1 vccd1 vccd1 _13634_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10846_ _10846_/A _10846_/B vssd1 vssd1 vccd1 vccd1 _10846_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11124__S1 _11065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19141_ _19272_/CLK _19141_/D vssd1 vssd1 vccd1 vccd1 _19141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16353_ _19953_/Q _16353_/B vssd1 vssd1 vccd1 vccd1 _16353_/Y sky130_fd_sc_hd__nand2_1
X_13565_ _13605_/S vssd1 vssd1 vccd1 vccd1 _13598_/S sky130_fd_sc_hd__clkbuf_2
X_10777_ _10777_/A _18677_/Q vssd1 vssd1 vccd1 vccd1 _10777_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10788__B1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15304_ _19162_/Q _15197_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _15305_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12516_ _17234_/A _12545_/C vssd1 vssd1 vccd1 vccd1 _12516_/X sky130_fd_sc_hd__or2_1
X_19072_ _19200_/CLK _19072_/D vssd1 vssd1 vccd1 vccd1 _19072_/Q sky130_fd_sc_hd__dfxtp_1
X_16284_ _16290_/B _16283_/Y _12444_/X vssd1 vssd1 vccd1 vccd1 _16285_/B sky130_fd_sc_hd__a21oi_2
X_13496_ _19734_/Q vssd1 vssd1 vccd1 vccd1 _16925_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13839__S _13845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15235_ _15235_/A vssd1 vssd1 vccd1 vccd1 _15235_/X sky130_fd_sc_hd__clkbuf_2
X_18023_ _18023_/A _18023_/B vssd1 vssd1 vccd1 vccd1 _18023_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12447_ _12441_/X _12442_/X _12446_/X _12494_/A vssd1 vssd1 vccd1 vccd1 _12447_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output90_A _12509_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15166_ _15166_/A vssd1 vssd1 vccd1 vccd1 _19114_/D sky130_fd_sc_hd__clkbuf_1
X_12378_ _12378_/A _12378_/B vssd1 vssd1 vccd1 vccd1 _12378_/X sky130_fd_sc_hd__or2_2
XFILLER_154_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14117_ _14117_/A vssd1 vssd1 vccd1 vccd1 _18684_/D sky130_fd_sc_hd__clkbuf_1
X_11329_ _18795_/Q _19130_/Q _11329_/S vssd1 vssd1 vccd1 vccd1 _11330_/B sky130_fd_sc_hd__mux2_1
X_15097_ _14624_/X _19081_/Q _15105_/S vssd1 vssd1 vccd1 vccd1 _15098_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12044__A _12137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19974_ _19978_/CLK _19974_/D vssd1 vssd1 vccd1 vccd1 _19974_/Q sky130_fd_sc_hd__dfxtp_1
X_18925_ _19063_/CLK _18925_/D vssd1 vssd1 vccd1 vccd1 _18925_/Q sky130_fd_sc_hd__dfxtp_1
X_14048_ _14059_/A vssd1 vssd1 vccd1 vccd1 _14057_/S sky130_fd_sc_hd__buf_2
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18856_ _19570_/CLK _18856_/D vssd1 vssd1 vccd1 vccd1 _18856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17807_ _17624_/X _17797_/X _17806_/X _18007_/A _11972_/Y vssd1 vssd1 vccd1 vccd1
+ _17807_/X sky130_fd_sc_hd__a32o_1
XANTENNA__17640__A1 _17607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18787_ _19412_/CLK _18787_/D vssd1 vssd1 vccd1 vccd1 _18787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15999_ _13069_/X _19423_/Q _16001_/S vssd1 vssd1 vccd1 vccd1 _16000_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17738_ _17736_/X _17737_/X _17810_/S vssd1 vssd1 vccd1 vccd1 _17738_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11363__S1 _09957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17669_ _17754_/A vssd1 vssd1 vccd1 vccd1 _18007_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19408_ _19409_/CLK _19408_/D vssd1 vssd1 vccd1 vccd1 _19408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19339_ _19873_/CLK _19339_/D vssd1 vssd1 vccd1 vccd1 _19339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_173_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10874__S0 _09983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17729__B _17729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10626__S0 _10625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10173__S _10173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09925_ _09925_/A vssd1 vssd1 vccd1 vccd1 _09925_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20045_ _20052_/CLK _20045_/D vssd1 vssd1 vccd1 vccd1 _20045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09856_ _10497_/A vssd1 vssd1 vccd1 vccd1 _10393_/A sky130_fd_sc_hd__clkbuf_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09795__S1 _09730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_98_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _18823_/Q _19158_/Q _09787_/S vssd1 vssd1 vccd1 vccd1 _09788_/B sky130_fd_sc_hd__mux2_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18295__B _18326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15712__B _17175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14609__A _14676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17934__A2 _17937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10700_ _18679_/Q _19174_/Q _10700_/S vssd1 vssd1 vccd1 vccd1 _10701_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15204__S _15213_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11645_/B _11785_/A _11680_/C _11680_/D vssd1 vssd1 vccd1 vccd1 _12596_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _18649_/Q _19240_/Q _19402_/Q _18617_/Q _10678_/S _10604_/A vssd1 vssd1 vccd1
+ vccd1 _10632_/B sky130_fd_sc_hd__mux4_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12129__A _17187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09624__B2 _19924_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11431__A1 _09814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13350_ _19912_/Q _15768_/B _13534_/S vssd1 vssd1 vccd1 vccd1 _13350_/X sky130_fd_sc_hd__mux2_1
X_10562_ _10462_/X _10559_/X _10561_/X vssd1 vssd1 vccd1 vccd1 _10562_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12301_ _17389_/A _12301_/B vssd1 vssd1 vccd1 vccd1 _12302_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ _19940_/Q vssd1 vssd1 vccd1 vccd1 _13282_/A sky130_fd_sc_hd__clkbuf_2
X_10493_ _10486_/Y _10488_/Y _10490_/Y _10492_/Y _09718_/A vssd1 vssd1 vccd1 vccd1
+ _10493_/X sky130_fd_sc_hd__o221a_1
XFILLER_136_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15020_ _19047_/Q _14414_/X _15022_/S vssd1 vssd1 vccd1 vccd1 _15021_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13184__B2 _19523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09438__A _18333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ _12232_/A _12232_/B vssd1 vssd1 vccd1 vccd1 _12233_/A sky130_fd_sc_hd__xnor2_4
XFILLER_142_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12931__A1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ _12188_/A _12650_/A _12162_/Y vssd1 vssd1 vccd1 vccd1 _17918_/B sky130_fd_sc_hd__a21o_2
XANTENNA__10093__S1 _10813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10942__B1 _10941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11114_ _18799_/Q _19134_/Q _11114_/S vssd1 vssd1 vccd1 vccd1 _11115_/B sky130_fd_sc_hd__mux2_1
XANTENNA__17870__A1 _17705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16971_ _19747_/Q _19746_/Q _16971_/C vssd1 vssd1 vccd1 vccd1 _16972_/C sky130_fd_sc_hd__and3_1
X_12094_ _12089_/X _12090_/X _12093_/X vssd1 vssd1 vccd1 vccd1 _12095_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__12799__A _12837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18710_ _19301_/CLK _18710_/D vssd1 vssd1 vccd1 vccd1 _18710_/Q sky130_fd_sc_hd__dfxtp_1
X_15922_ _15922_/A vssd1 vssd1 vccd1 vccd1 _19388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11045_ _19458_/Q _19296_/Q _18705_/Q _18475_/Q _10914_/X _10969_/A vssd1 vssd1 vccd1
+ vccd1 _11046_/B sky130_fd_sc_hd__mux4_1
XFILLER_89_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10811__S _10811_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19690_ _19804_/CLK _19690_/D vssd1 vssd1 vccd1 vccd1 _19690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18641_ _19490_/CLK _18641_/D vssd1 vssd1 vccd1 vccd1 _18641_/Q sky130_fd_sc_hd__dfxtp_1
X_15853_ _13056_/X _19358_/Q _15857_/S vssd1 vssd1 vccd1 vccd1 _15854_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10170__B2 _19916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15903__A _15903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804_ _18955_/Q _14443_/X _14808_/S vssd1 vssd1 vccd1 vccd1 _14805_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10112__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18572_ _19734_/CLK _18572_/D vssd1 vssd1 vccd1 vccd1 _18572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12996_ _19738_/Q _12991_/X _12994_/X _12995_/X vssd1 vssd1 vccd1 vccd1 _12996_/X
+ sky130_fd_sc_hd__a211o_2
X_15784_ _13587_/X _15782_/X _15783_/Y _12770_/X _18458_/Q vssd1 vssd1 vccd1 vccd1
+ _15784_/X sky130_fd_sc_hd__a32o_2
XFILLER_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17523_ _17919_/A vssd1 vssd1 vccd1 vccd1 _17995_/A sky130_fd_sc_hd__clkbuf_2
X_14735_ _18920_/Q _14449_/X _14735_/S vssd1 vssd1 vccd1 vccd1 _14736_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11947_ _11942_/X _11944_/X _11946_/Y vssd1 vssd1 vccd1 vccd1 _11947_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15114__S _15116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13423__A _15273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _14666_/A vssd1 vssd1 vccd1 vccd1 _14666_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17454_ _17508_/S vssd1 vssd1 vccd1 vccd1 _17573_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11878_ _13172_/A _09352_/X _11839_/C vssd1 vssd1 vccd1 vccd1 _11878_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16405_ _16405_/A vssd1 vssd1 vccd1 vccd1 _19560_/D sky130_fd_sc_hd__clkbuf_1
X_13617_ _15203_/A vssd1 vssd1 vccd1 vccd1 _14580_/A sky130_fd_sc_hd__clkbuf_2
X_10829_ _10825_/X _10827_/X _10828_/X _10840_/A _09964_/X vssd1 vssd1 vccd1 vccd1
+ _10834_/B sky130_fd_sc_hd__o221a_1
XANTENNA__13142__B _13142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14953__S _14961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17385_ _17534_/B vssd1 vssd1 vccd1 vccd1 _17545_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14597_ _14596_/X _18870_/Q _14606_/S vssd1 vssd1 vccd1 vccd1 _14598_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12039__A _18347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19124_ _19572_/CLK _19124_/D vssd1 vssd1 vccd1 vccd1 _19124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13548_ _19881_/Q _12842_/X _12863_/X _19848_/Q _13547_/X vssd1 vssd1 vccd1 vccd1
+ _13548_/X sky130_fd_sc_hd__a221o_1
X_16336_ _19538_/Q _16300_/X _16334_/Y _16335_/Y vssd1 vssd1 vccd1 vccd1 _19538_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16453__B _16453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19055_ _19504_/CLK _19055_/D vssd1 vssd1 vccd1 vccd1 _19055_/Q sky130_fd_sc_hd__dfxtp_1
X_16267_ _16273_/B _16267_/B vssd1 vssd1 vccd1 vccd1 _16267_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10782__A _10794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13479_ _19765_/Q _12692_/A _13478_/X _12714_/A vssd1 vssd1 vccd1 vccd1 _13479_/X
+ sky130_fd_sc_hd__a211o_1
X_18006_ _10360_/Y _09464_/X _18005_/X vssd1 vssd1 vccd1 vccd1 _19913_/D sky130_fd_sc_hd__a21oi_1
X_15218_ _15218_/A vssd1 vssd1 vccd1 vccd1 _19135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09348__A _19888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16198_ _19512_/Q _14666_/A _16200_/S vssd1 vssd1 vccd1 vccd1 _16199_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15149_ _19106_/Q vssd1 vssd1 vccd1 vccd1 _15150_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19957_ _20000_/CLK _19957_/D vssd1 vssd1 vccd1 vccd1 _19957_/Q sky130_fd_sc_hd__dfxtp_2
X_09710_ _09891_/A vssd1 vssd1 vccd1 vccd1 _09711_/A sky130_fd_sc_hd__clkbuf_2
X_18908_ _19557_/CLK _18908_/D vssd1 vssd1 vccd1 vccd1 _18908_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15085__A _15131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19888_ _19888_/CLK _19888_/D vssd1 vssd1 vccd1 vccd1 _19888_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12321__A2_N _12657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ _11280_/S vssd1 vssd1 vccd1 vccd1 _11222_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18839_ _19200_/CLK _18839_/D vssd1 vssd1 vccd1 vccd1 _18839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18396__A _18396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09572_ _10166_/A _09572_/B vssd1 vssd1 vccd1 vccd1 _09572_/X sky130_fd_sc_hd__or2_1
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14148__B _15198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11788__A _20028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17475__A _17507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10075__S1 _10609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09908_ _10254_/A _09908_/B vssd1 vssd1 vccd1 vccd1 _09908_/X sky130_fd_sc_hd__or2_1
XFILLER_104_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09768__S1 _09569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09839_ _19477_/Q _19315_/Q _18724_/Q _18494_/Q _10160_/S _09809_/A vssd1 vssd1 vccd1
+ vccd1 _09839_/X sky130_fd_sc_hd__mux4_2
X_20028_ _20032_/CLK _20028_/D vssd1 vssd1 vccd1 vccd1 _20028_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13942__S _13950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ _19653_/Q _12832_/X _12833_/X _19785_/Q _12849_/X vssd1 vssd1 vccd1 vccd1
+ _12851_/B sky130_fd_sc_hd__a221o_2
XFILLER_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _20039_/Q vssd1 vssd1 vccd1 vccd1 _18319_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12781_ _19812_/Q _12677_/A _12802_/A _19342_/Q vssd1 vssd1 vccd1 vccd1 _12781_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _13774_/X _18839_/Q _14524_/S vssd1 vssd1 vccd1 vccd1 _14521_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11732_ _12598_/A _12598_/B vssd1 vssd1 vccd1 vccd1 _11733_/C sky130_fd_sc_hd__nand2_1
XFILLER_54_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14451_/A vssd1 vssd1 vccd1 vccd1 _18819_/D sky130_fd_sc_hd__clkbuf_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11663_ _20028_/Q _11663_/B _11663_/C vssd1 vssd1 vccd1 vccd1 _12207_/D sky130_fd_sc_hd__or3_2
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14773__S _14775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13402_ _19872_/Q _12913_/X _13343_/X _19839_/Q vssd1 vssd1 vccd1 vccd1 _13402_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09867__S _10218_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10614_ _10824_/S vssd1 vssd1 vccd1 vccd1 _10614_/X sky130_fd_sc_hd__clkbuf_4
X_17170_ _19823_/Q _17180_/B vssd1 vssd1 vccd1 vccd1 _17170_/X sky130_fd_sc_hd__or2_1
XFILLER_168_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11404__B2 _11403_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14382_ _14586_/A vssd1 vssd1 vccd1 vccd1 _14382_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11594_ _11549_/X _11550_/Y _11551_/X _11552_/Y _11593_/X vssd1 vssd1 vccd1 vccd1
+ _11594_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16121_ _16121_/A vssd1 vssd1 vccd1 vccd1 _19477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13333_ _13333_/A vssd1 vssd1 vccd1 vccd1 _18487_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10612__C1 _09475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A _20028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10545_ _19500_/Q _18912_/Q _18949_/Q _18523_/Q _10266_/A _10332_/A vssd1 vssd1 vccd1
+ vccd1 _10545_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14074__A _14074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ _13487_/X _19447_/Q _16056_/S vssd1 vssd1 vccd1 vccd1 _16053_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13157__B2 _19522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13264_ _19864_/Q _12842_/A _12695_/A _17192_/A vssd1 vssd1 vccd1 vccd1 _13264_/X
+ sky130_fd_sc_hd__a22o_1
X_10476_ _10476_/A _10476_/B vssd1 vssd1 vccd1 vccd1 _10476_/X sky130_fd_sc_hd__or2_1
XFILLER_142_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15003_ _19039_/Q _14388_/X _15011_/S vssd1 vssd1 vccd1 vccd1 _15004_/A sky130_fd_sc_hd__mux2_1
X_12215_ _12314_/A vssd1 vssd1 vccd1 vccd1 _12215_/X sky130_fd_sc_hd__buf_2
XANTENNA__18096__A1 _19921_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17385__A _17534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12904__B2 _18460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10107__A _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13195_ _15228_/A vssd1 vssd1 vccd1 vccd1 _13195_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09318__D _20041_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19811_ _19857_/CLK _19811_/D vssd1 vssd1 vccd1 vccd1 _19811_/Q sky130_fd_sc_hd__dfxtp_1
X_12146_ _12108_/A _17884_/B _12111_/A _12111_/B vssd1 vssd1 vccd1 vccd1 _12147_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_121_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19742_ _19745_/CLK _19742_/D vssd1 vssd1 vccd1 vccd1 _19742_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11015__S0 _10893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__A _13418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16954_ _16958_/A _16958_/B _16957_/C _19738_/Q vssd1 vssd1 vccd1 vccd1 _16955_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__14013__S _14013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ _12075_/Y _12076_/Y _12077_/S vssd1 vssd1 vccd1 vccd1 _12080_/B sky130_fd_sc_hd__mux2_1
XFILLER_110_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15905_ _15905_/A vssd1 vssd1 vccd1 vccd1 _19381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11028_ _18827_/Q vssd1 vssd1 vccd1 vccd1 _11327_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_38_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17832__B _17832_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19673_ _19877_/CLK _19673_/D vssd1 vssd1 vccd1 vccd1 _19673_/Q sky130_fd_sc_hd__dfxtp_1
X_16885_ _16922_/B _16922_/C _16888_/D _16875_/X vssd1 vssd1 vccd1 vccd1 _16885_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11340__B1 _10988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18624_ _19412_/CLK _18624_/D vssd1 vssd1 vccd1 vccd1 _18624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15836_ _15836_/A vssd1 vssd1 vccd1 vccd1 _19353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11891__B2 _11890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09631__A _10794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18555_ _19563_/CLK _18555_/D vssd1 vssd1 vccd1 vccd1 _18555_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10777__A _10777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ _18464_/Q _12973_/X _10137_/A _12976_/X vssd1 vssd1 vccd1 vccd1 _18464_/D
+ sky130_fd_sc_hd__a22o_1
X_15767_ _15767_/A vssd1 vssd1 vccd1 vccd1 _19342_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17359__B1 _18273_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11372__S _11372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17506_ _12529_/A _17702_/B _17506_/S vssd1 vssd1 vccd1 vccd1 _17506_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14718_ _18912_/Q _14424_/X _14724_/S vssd1 vssd1 vccd1 vccd1 _14719_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18486_ _19563_/CLK _18486_/D vssd1 vssd1 vccd1 vccd1 _18486_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09931__S1 _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15698_ _15697_/X _19330_/Q _15720_/S vssd1 vssd1 vccd1 vccd1 _15699_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17437_ _17434_/X _17435_/X _17565_/S vssd1 vssd1 vccd1 vccd1 _17437_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10851__C1 _10794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14649_ _14649_/A vssd1 vssd1 vccd1 vccd1 _18886_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12992__A _12992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14683__S _14691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16464__A _16875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_46_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17368_ _17368_/A vssd1 vssd1 vccd1 vccd1 _19889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10749__A3 _10748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19107_ _19203_/CLK _19107_/D vssd1 vssd1 vccd1 vccd1 _19107_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13600__B _13600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16319_ _19535_/Q _16318_/X _16325_/S vssd1 vssd1 vccd1 vccd1 _16320_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17299_ _17299_/A vssd1 vssd1 vccd1 vccd1 _19872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13148__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19038_ _19486_/CLK _19038_/D vssd1 vssd1 vccd1 vccd1 _19038_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput101 _12003_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[8] sky130_fd_sc_hd__buf_2
XANTENNA__11159__B1 _11135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput112 _12648_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[12] sky130_fd_sc_hd__buf_2
Xoutput123 _12660_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[22] sky130_fd_sc_hd__buf_2
XANTENNA__15808__A _15808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12931__S _17808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput134 _12635_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[3] sky130_fd_sc_hd__buf_2
XFILLER_114_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput145 _12133_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[12] sky130_fd_sc_hd__buf_2
XANTENNA__10017__A _10017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput156 _12401_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[22] sky130_fd_sc_hd__buf_2
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput167 _16453_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_141_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11006__S0 _09530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13320__A1 _13060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13762__S _13765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09624_ _09589_/X _09606_/X _09616_/X _09623_/X _19924_/Q vssd1 vssd1 vccd1 vccd1
+ _12593_/A sky130_fd_sc_hd__a32oi_4
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16270__A0 _19526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09541__A _09761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__S1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09555_ _11204_/A vssd1 vssd1 vccd1 vccd1 _11016_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09486_ _10840_/A vssd1 vssd1 vccd1 vccd1 _10574_/A sky130_fd_sc_hd__buf_4
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12407__A _12407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13139__A1 _19521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ _10330_/A vssd1 vssd1 vccd1 vccd1 _10330_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13937__S _13939_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ _09820_/X _10254_/X _10256_/X _10260_/X _09605_/A vssd1 vssd1 vccd1 vccd1
+ _10261_/X sky130_fd_sc_hd__a311o_1
XANTENNA__11245__S0 _11129_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12000_ _11938_/A _11936_/B _11971_/A _11999_/X vssd1 vssd1 vccd1 vccd1 _12000_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_79_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17825__A1 _12003_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__A _10063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _19916_/Q vssd1 vssd1 vccd1 vccd1 _10192_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13951_ _13951_/A vssd1 vssd1 vccd1 vccd1 _18612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12902_ _15680_/A _18460_/Q vssd1 vssd1 vccd1 vccd1 _12902_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13882_ _13882_/A vssd1 vssd1 vccd1 vccd1 _18581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16670_ _19665_/Q _16670_/B _16670_/C vssd1 vssd1 vccd1 vccd1 _16672_/B sky130_fd_sc_hd__and3_1
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12796__B input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09451__A _20049_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15621_ _15621_/A vssd1 vssd1 vccd1 vccd1 _19303_/D sky130_fd_sc_hd__clkbuf_1
X_12833_ _13117_/A vssd1 vssd1 vccd1 vccd1 _12833_/X sky130_fd_sc_hd__buf_2
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _18340_/A _18349_/B vssd1 vssd1 vccd1 vccd1 _18340_/X sky130_fd_sc_hd__or2_1
XANTENNA__11086__C1 _09659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15574_/A vssd1 vssd1 vccd1 vccd1 _15561_/S sky130_fd_sc_hd__clkbuf_4
X_12764_ _19627_/Q _13142_/B _12763_/X vssd1 vssd1 vccd1 vccd1 _12764_/Y sky130_fd_sc_hd__o21ai_4
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _14559_/A vssd1 vssd1 vccd1 vccd1 _14572_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__10833__C1 _10621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11715_ _11764_/C vssd1 vssd1 vccd1 vccd1 _17610_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15483_ _19242_/Q _15251_/X _15489_/S vssd1 vssd1 vccd1 vccd1 _15484_/A sky130_fd_sc_hd__mux2_1
X_18271_ _18352_/A _18271_/B vssd1 vssd1 vccd1 vccd1 _18272_/A sky130_fd_sc_hd__or2_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12695_/A vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13701__A _15267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17222_ _17220_/Y _17212_/X _17221_/X _17215_/X vssd1 vssd1 vccd1 vccd1 _19840_/D
+ sky130_fd_sc_hd__o211a_1
X_14434_ _18814_/Q _14433_/X _14434_/S vssd1 vssd1 vccd1 vccd1 _14435_/A sky130_fd_sc_hd__mux2_1
X_11646_ _11678_/A _11680_/C _11646_/C _17337_/A vssd1 vssd1 vccd1 vccd1 _11697_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_156_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 io_dbus_rdata[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_2
Xinput25 io_dbus_rdata[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_4
XFILLER_156_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14365_ _18793_/Q _13739_/X _14367_/S vssd1 vssd1 vccd1 vccd1 _14366_/A sky130_fd_sc_hd__mux2_1
X_17153_ _17229_/A vssd1 vssd1 vccd1 vccd1 _17153_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16316__A1 _19534_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput36 io_ibus_inst[11] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
X_11577_ _11578_/A _11575_/C _11575_/A vssd1 vssd1 vccd1 vccd1 _11577_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16316__B2 _16315_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput47 io_ibus_inst[21] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_4
XFILLER_116_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16104_ _13331_/X _19470_/Q _16106_/S vssd1 vssd1 vccd1 vccd1 _16105_/A sky130_fd_sc_hd__mux2_1
Xinput58 io_ibus_inst[31] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_1
X_13316_ _13316_/A _13316_/B _13316_/C _12764_/Y vssd1 vssd1 vccd1 vccd1 _13316_/X
+ sky130_fd_sc_hd__or4b_2
Xinput69 io_irq_uart_irq vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_4
X_10528_ _10314_/A _10521_/X _10523_/X _10527_/X _09604_/A vssd1 vssd1 vccd1 vccd1
+ _10528_/X sky130_fd_sc_hd__a311o_2
X_17084_ _19789_/Q _17081_/B _17083_/Y vssd1 vssd1 vccd1 vccd1 _19789_/D sky130_fd_sc_hd__o21a_1
XFILLER_115_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14296_ _15061_/A _18297_/A _18295_/A _14844_/D vssd1 vssd1 vccd1 vccd1 _15517_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_109_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16035_ _16035_/A vssd1 vssd1 vccd1 vccd1 _19439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13247_ _19337_/Q _13245_/X _12758_/A _19527_/Q _13246_/X vssd1 vssd1 vccd1 vccd1
+ _13247_/X sky130_fd_sc_hd__a221o_1
X_10459_ _10459_/A _12655_/B vssd1 vssd1 vccd1 vccd1 _10460_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13178_ _15225_/A vssd1 vssd1 vccd1 vccd1 _13178_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12129_ _17187_/A _12157_/C vssd1 vssd1 vccd1 vccd1 _12129_/X sky130_fd_sc_hd__or2_1
XFILLER_112_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17986_ _18033_/A _17989_/B _17539_/A _17985_/Y vssd1 vssd1 vccd1 vccd1 _17986_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_111_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19725_ _19737_/CLK _19725_/D vssd1 vssd1 vccd1 vccd1 _19725_/Q sky130_fd_sc_hd__dfxtp_1
X_16937_ _19741_/Q _19740_/Q vssd1 vssd1 vccd1 vccd1 _16964_/A sky130_fd_sc_hd__and2_1
XFILLER_78_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19656_ _19792_/CLK _19656_/D vssd1 vssd1 vccd1 vccd1 _19656_/Q sky130_fd_sc_hd__dfxtp_1
X_16868_ _19719_/Q _19718_/Q _16868_/C _16868_/D vssd1 vssd1 vccd1 vccd1 _16873_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__16252__A0 _19523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18607_ _19486_/CLK _18607_/D vssd1 vssd1 vccd1 vccd1 _18607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15819_ _19886_/Q _15819_/B vssd1 vssd1 vccd1 vccd1 _15819_/Y sky130_fd_sc_hd__nor2_4
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19587_ _19963_/CLK _19587_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16799_ _16818_/A _16799_/B vssd1 vssd1 vccd1 vccd1 _16799_/Y sky130_fd_sc_hd__nor2_1
X_09340_ _15819_/B _16809_/B _12739_/A vssd1 vssd1 vccd1 vccd1 _12678_/A sky130_fd_sc_hd__a21oi_2
XFILLER_80_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18538_ _19577_/CLK _18538_/D vssd1 vssd1 vccd1 vccd1 _18538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09271_ _09191_/B _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09329_/A sky130_fd_sc_hd__nand3b_2
X_18469_ _19671_/CLK _18469_/D vssd1 vssd1 vccd1 vccd1 _18469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10278__S1 _09887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17504__A0 _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12592__A2 _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11227__S0 _11085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17807__B2 _11972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15833__A3 _15819_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15273__A _15273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10202__S1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09607_ _09608_/A _09282_/X _09287_/X _09295_/X _18928_/Q vssd1 vssd1 vccd1 vccd1
+ _09617_/A sky130_fd_sc_hd__o2111a_4
XFILLER_113_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09538_ _10416_/S vssd1 vssd1 vccd1 vccd1 _10195_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16816__B _17346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ _18968_/Q vssd1 vssd1 vccd1 vccd1 _09470_/A sky130_fd_sc_hd__inv_2
XFILLER_106_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11500_ _18601_/Q _18862_/Q _18761_/Q _19096_/Q _10119_/X _10054_/A vssd1 vssd1 vccd1
+ vccd1 _11500_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12480_ _12480_/A vssd1 vssd1 vccd1 vccd1 _18068_/B sky130_fd_sc_hd__buf_2
XFILLER_138_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11431_ _09814_/A _11428_/X _11430_/X vssd1 vssd1 vccd1 vccd1 _11431_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12137__A _12137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14150_ _14844_/C _16809_/C _14000_/B vssd1 vssd1 vccd1 vccd1 _16371_/C sky130_fd_sc_hd__o21ai_1
XFILLER_164_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11362_ _11362_/A _11362_/B vssd1 vssd1 vccd1 vccd1 _11362_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13101_ _19329_/Q _12707_/X _13099_/X _19519_/Q _13100_/X vssd1 vssd1 vccd1 vccd1
+ _13101_/X sky130_fd_sc_hd__a221o_1
X_10313_ _19504_/Q _18916_/Q _18953_/Q _18527_/Q _10302_/X _10312_/X vssd1 vssd1 vccd1
+ vccd1 _10313_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14081_ _18668_/Q _13618_/X _14087_/S vssd1 vssd1 vccd1 vccd1 _14082_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16043__S _16045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ _11170_/A _11292_/X _10988_/A vssd1 vssd1 vccd1 vccd1 _11293_/Y sky130_fd_sc_hd__o21ai_1
X_13032_ input12/X _12988_/X _13031_/X _13007_/X vssd1 vssd1 vccd1 vccd1 _15203_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_98_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input52_A io_ibus_inst[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ _18816_/Q _19151_/Q _10244_/S vssd1 vssd1 vccd1 vccd1 _10244_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13532__B2 _19544_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09446__A _17331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15882__S _15890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17840_ _17624_/X _17835_/X _17839_/X _18007_/A _12024_/Y vssd1 vssd1 vccd1 vccd1
+ _17840_/X sky130_fd_sc_hd__a32o_1
X_10175_ _18818_/Q _19153_/Q _10175_/S vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__mux2_1
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17771_ _17791_/A vssd1 vssd1 vccd1 vccd1 _17771_/X sky130_fd_sc_hd__clkbuf_2
X_14983_ _19031_/Q _14465_/X _14983_/S vssd1 vssd1 vccd1 vccd1 _14984_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output139_A _12643_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19510_ _19510_/CLK _19510_/D vssd1 vssd1 vccd1 vccd1 _19510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16722_ _19678_/Q _16718_/C _16721_/Y vssd1 vssd1 vccd1 vccd1 _19678_/D sky130_fd_sc_hd__o21a_1
X_13934_ _13934_/A vssd1 vssd1 vccd1 vccd1 _18604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12600__A _12600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16234__B1 _12444_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19441_ _19566_/CLK _19441_/D vssd1 vssd1 vccd1 vccd1 _19441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16653_ _19659_/Q _16653_/B _16653_/C vssd1 vssd1 vccd1 vccd1 _16655_/B sky130_fd_sc_hd__and3_1
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13865_ _13761_/X _18574_/Q _13867_/S vssd1 vssd1 vccd1 vccd1 _13866_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11216__A _11216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15604_ _15604_/A vssd1 vssd1 vccd1 vccd1 _19295_/D sky130_fd_sc_hd__clkbuf_1
X_19372_ _19561_/CLK _19372_/D vssd1 vssd1 vccd1 vccd1 _19372_/Q sky130_fd_sc_hd__dfxtp_1
X_12816_ _15700_/A _12815_/Y _12853_/A vssd1 vssd1 vccd1 vccd1 _12816_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16584_ _19635_/Q _16584_/B vssd1 vssd1 vccd1 vccd1 _16590_/C sky130_fd_sc_hd__and2_1
X_13796_ _14621_/A vssd1 vssd1 vccd1 vccd1 _13796_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_90_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18323_ _18323_/A vssd1 vssd1 vccd1 vccd1 _18323_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ _19265_/Q _15222_/X _15539_/S vssd1 vssd1 vccd1 vccd1 _15536_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12747_/A vssd1 vssd1 vccd1 vccd1 _17319_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17734__B1 _18019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _18254_/A vssd1 vssd1 vccd1 vccd1 _19981_/D sky130_fd_sc_hd__clkbuf_1
X_12678_ _12678_/A vssd1 vssd1 vccd1 vccd1 _17149_/A sky130_fd_sc_hd__clkbuf_2
X_15466_ _15466_/A vssd1 vssd1 vccd1 vccd1 _19234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10774__B _12647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17205_ _17205_/A _17210_/B vssd1 vssd1 vccd1 vccd1 _17205_/X sky130_fd_sc_hd__or2_1
X_14417_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14417_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11629_ _11629_/A vssd1 vssd1 vccd1 vccd1 _12595_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14961__S _14961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18185_ _18185_/A vssd1 vssd1 vccd1 vccd1 _19950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15397_ _15443_/S vssd1 vssd1 vccd1 vccd1 _15406_/S sky130_fd_sc_hd__buf_6
XFILLER_156_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17136_ input68/X _17138_/B vssd1 vssd1 vccd1 vccd1 _17136_/X sky130_fd_sc_hd__or2_1
XANTENNA__11231__C1 _09736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14348_ _18785_/Q _13706_/X _14352_/S vssd1 vssd1 vccd1 vccd1 _14349_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16461__B _16461_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15358__A _15358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14279_ _13828_/X _18755_/Q _14279_/S vssd1 vssd1 vccd1 vccd1 _14280_/A sky130_fd_sc_hd__mux2_1
X_17067_ _19783_/Q hold19/X _17066_/Y vssd1 vssd1 vccd1 vccd1 _19783_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16018_ _16018_/A vssd1 vssd1 vccd1 vccd1 _19431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17969_ _12260_/A _17844_/X _17968_/X _17858_/X vssd1 vssd1 vccd1 vccd1 _17969_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19708_ _19718_/CLK _19708_/D vssd1 vssd1 vccd1 vccd1 _19708_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11298__C1 _10994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19639_ _19769_/CLK _19639_/D vssd1 vssd1 vccd1 vccd1 _19639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16917__A _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10030__A _10030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09323_ _19885_/Q vssd1 vssd1 vccd1 vccd1 _15819_/B sky130_fd_sc_hd__buf_2
XFILLER_80_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16128__S _16128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10499__S1 _10397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14437__A _14453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ _09425_/B vssd1 vssd1 vccd1 vccd1 _11645_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09185_ _20035_/Q vssd1 vssd1 vccd1 vccd1 _09272_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_153_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13514__B2 _19846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10205__A _10205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_168_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15207__S _15213_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11828__A1 _19517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11980_ _11885_/B _11917_/Y _11953_/Y _11954_/Y _11956_/A vssd1 vssd1 vccd1 vccd1
+ _11980_/Y sky130_fd_sc_hd__a311oi_2
XFILLER_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16216__B1 _13597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10931_ _10051_/A _10930_/X _09999_/A vssd1 vssd1 vccd1 vccd1 _10931_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13950__S _13950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10862_ _11399_/A _10862_/B vssd1 vssd1 vccd1 vccd1 _10862_/Y sky130_fd_sc_hd__nor2_1
X_13650_ _15228_/A vssd1 vssd1 vccd1 vccd1 _14605_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14839__A2_N _16315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12601_ _12601_/A _12601_/B vssd1 vssd1 vccd1 vccd1 _12601_/Y sky130_fd_sc_hd__nor2_2
XFILLER_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _18438_/Q _13029_/X _13579_/Y _13580_/X vssd1 vssd1 vccd1 vccd1 _13581_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13450__A0 _19918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _19366_/Q _18980_/Q _19430_/Q _18549_/Q _10849_/S _11496_/A vssd1 vssd1 vccd1
+ vccd1 _10794_/B sky130_fd_sc_hd__mux4_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12532_ _12532_/A _12532_/B vssd1 vssd1 vccd1 vccd1 _12534_/C sky130_fd_sc_hd__nand2_1
X_15320_ _15320_/A vssd1 vssd1 vccd1 vccd1 _19169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15877__S _15879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11439__S0 _10690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15251_ _15251_/A vssd1 vssd1 vccd1 vccd1 _15251_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12463_ _12463_/A vssd1 vssd1 vccd1 vccd1 _12463_/Y sky130_fd_sc_hd__inv_4
XFILLER_12_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14202_ _14202_/A vssd1 vssd1 vccd1 vccd1 _18720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11414_ _11565_/A _11568_/A _11565_/C _10556_/A _11413_/X vssd1 vssd1 vccd1 vccd1
+ _11560_/C sky130_fd_sc_hd__a311o_1
X_15182_ _15182_/A vssd1 vssd1 vccd1 vccd1 _19122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12394_ _12394_/A _12438_/C vssd1 vssd1 vccd1 vccd1 _12394_/Y sky130_fd_sc_hd__nor2_1
X_14133_ _14133_/A vssd1 vssd1 vccd1 vccd1 _14142_/S sky130_fd_sc_hd__buf_4
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ _11338_/Y _11340_/Y _11342_/Y _11344_/Y _10994_/A vssd1 vssd1 vccd1 vccd1
+ _11345_/X sky130_fd_sc_hd__o221a_2
XFILLER_125_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19990_ _20027_/CLK _19990_/D vssd1 vssd1 vccd1 vccd1 _19990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14064_ _18662_/Q _13727_/X _14068_/S vssd1 vssd1 vccd1 vccd1 _14065_/A sky130_fd_sc_hd__mux2_1
X_18941_ _19204_/CLK _18941_/D vssd1 vssd1 vccd1 vccd1 _18941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11276_ _10875_/A _11269_/X _11271_/X _11275_/X _09599_/A vssd1 vssd1 vccd1 vccd1
+ _11276_/X sky130_fd_sc_hd__a311o_4
X_13015_ _19887_/Q _13748_/B vssd1 vssd1 vccd1 vccd1 _14000_/B sky130_fd_sc_hd__and2_1
X_10227_ _10220_/X _10222_/Y _10224_/Y _10226_/Y _09741_/X vssd1 vssd1 vccd1 vccd1
+ _10227_/X sky130_fd_sc_hd__o221a_2
XANTENNA__10414__S1 _09841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18872_ _19288_/CLK _18872_/D vssd1 vssd1 vccd1 vccd1 _18872_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14810__A _14810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17823_ _17765_/X _17812_/X _17822_/X _17619_/A vssd1 vssd1 vccd1 vccd1 _17823_/X
+ sky130_fd_sc_hd__a211o_1
X_10158_ _09479_/A _10150_/X _10153_/X _10157_/X _09605_/X vssd1 vssd1 vccd1 vccd1
+ _10158_/X sky130_fd_sc_hd__a311o_1
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_12_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17754_ _17754_/A vssd1 vssd1 vccd1 vccd1 _17755_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14966_ _19023_/Q _14440_/X _14972_/S vssd1 vssd1 vccd1 vccd1 _14967_/A sky130_fd_sc_hd__mux2_1
X_10089_ _10746_/A _10086_/X _10088_/X _10621_/A vssd1 vssd1 vccd1 vccd1 _10090_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16207__B1 _13592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16705_ _19803_/Q _19802_/Q _19804_/Q _17115_/A vssd1 vssd1 vccd1 vccd1 _16710_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_63_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13917_ _13917_/A vssd1 vssd1 vccd1 vccd1 _18597_/D sky130_fd_sc_hd__clkbuf_1
X_17685_ _17569_/X _17573_/X _17685_/S vssd1 vssd1 vccd1 vccd1 _17685_/X sky130_fd_sc_hd__mux2_1
X_14897_ _14897_/A vssd1 vssd1 vccd1 vccd1 _18992_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09893__C1 _09719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19424_ _19455_/CLK _19424_/D vssd1 vssd1 vccd1 vccd1 _19424_/Q sky130_fd_sc_hd__dfxtp_1
X_16636_ _19653_/Q _16636_/B _16636_/C vssd1 vssd1 vccd1 vccd1 _16638_/B sky130_fd_sc_hd__and3_1
X_13848_ _13847_/X _18569_/Q _13851_/S vssd1 vssd1 vccd1 vccd1 _13849_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19355_ _19762_/CLK _19355_/D vssd1 vssd1 vccd1 vccd1 _19355_/Q sky130_fd_sc_hd__dfxtp_1
X_16567_ _16593_/A _16572_/C vssd1 vssd1 vccd1 vccd1 _16567_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13779_ _13779_/A vssd1 vssd1 vccd1 vccd1 _18547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18306_ _18306_/A _18331_/B vssd1 vssd1 vccd1 vccd1 _18306_/Y sky130_fd_sc_hd__nand2_1
X_15518_ _15574_/A vssd1 vssd1 vccd1 vccd1 _15587_/S sky130_fd_sc_hd__buf_6
XFILLER_148_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19286_ _19286_/CLK _19286_/D vssd1 vssd1 vccd1 vccd1 _19286_/Q sky130_fd_sc_hd__dfxtp_1
X_16498_ _19653_/Q _19652_/Q _19654_/Q _16630_/A vssd1 vssd1 vccd1 vccd1 _16640_/A
+ sky130_fd_sc_hd__and4_1
X_18237_ _18237_/A vssd1 vssd1 vccd1 vccd1 _19973_/D sky130_fd_sc_hd__clkbuf_1
X_15449_ _15449_/A vssd1 vssd1 vccd1 vccd1 _19226_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14691__S _14691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18132__A0 _16206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18168_ _16301_/B _19975_/Q _18170_/S vssd1 vssd1 vccd1 vccd1 _18169_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17119_ _17120_/B _17120_/C _17118_/Y vssd1 vssd1 vccd1 vccd1 _19802_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18099_ _17945_/A _18097_/B _17814_/X _18098_/X vssd1 vssd1 vccd1 vccd1 _18099_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16694__B1 _16667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09941_ _19476_/Q _19314_/Q _18723_/Q _18493_/Q _10218_/S _10271_/A vssd1 vssd1 vccd1
+ vccd1 _09941_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17507__S _17507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16411__S _16415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09872_ _10270_/S vssd1 vssd1 vccd1 vccd1 _09872_/X sky130_fd_sc_hd__clkbuf_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09814__A _09814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10191__C1 _09719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15027__S _15033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16647__A _16672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09306_ _17391_/A _17393_/B _17393_/A _11622_/A vssd1 vssd1 vccd1 vccd1 _11699_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_167_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17174__A1 _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10797__A1 _09693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _11629_/A _11729_/A vssd1 vssd1 vccd1 vccd1 _11650_/A sky130_fd_sc_hd__nor2_1
XANTENNA__17478__A _17507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_94_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11210__A2 _11199_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11130_ _19456_/Q _19294_/Q _18703_/Q _18473_/Q _11129_/X _11061_/A vssd1 vssd1 vccd1
+ vccd1 _11130_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11061_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11061_/X sky130_fd_sc_hd__and2_1
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10012_ _11395_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10012_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11973__B _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10182__C1 _09741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14820_ _14820_/A vssd1 vssd1 vccd1 vccd1 _18962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A io_dbus_rdata[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14751_ _14751_/A vssd1 vssd1 vccd1 vccd1 _18927_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11277__A2 _11267_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11963_ _12069_/A _12639_/B _12039_/C _18340_/A vssd1 vssd1 vccd1 vccd1 _17792_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13702_ _14644_/A vssd1 vssd1 vccd1 vccd1 _13702_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17470_ _17456_/X _17469_/X _17802_/B vssd1 vssd1 vccd1 vccd1 _17470_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10914_ _11026_/S vssd1 vssd1 vccd1 vccd1 _10914_/X sky130_fd_sc_hd__buf_4
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14682_ _14750_/S vssd1 vssd1 vccd1 vccd1 _14691_/S sky130_fd_sc_hd__buf_2
X_11894_ _11894_/A vssd1 vssd1 vccd1 vccd1 _11961_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16421_ _16421_/A vssd1 vssd1 vccd1 vccd1 _19567_/D sky130_fd_sc_hd__clkbuf_1
X_10845_ _19107_/Q _18873_/Q _19555_/Q _19203_/Q _10702_/S _09662_/A vssd1 vssd1 vccd1
+ vccd1 _10846_/B sky130_fd_sc_hd__mux4_1
X_13633_ _15215_/A vssd1 vssd1 vccd1 vccd1 _14592_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14077__A _14133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19140_ _19268_/CLK _19140_/D vssd1 vssd1 vccd1 vccd1 _19140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16352_ _19953_/Q _16353_/B vssd1 vssd1 vccd1 vccd1 _16361_/C sky130_fd_sc_hd__or2_2
X_10776_ _19172_/Q vssd1 vssd1 vccd1 vccd1 _10776_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17165__A1 _15688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13564_ _12214_/A _13561_/Y _13563_/Y vssd1 vssd1 vccd1 vccd1 _13605_/S sky130_fd_sc_hd__a21o_1
XFILLER_158_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10788__A1 _09693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15303_ _15371_/S vssd1 vssd1 vccd1 vccd1 _15312_/S sky130_fd_sc_hd__buf_2
X_12515_ _19844_/Q vssd1 vssd1 vccd1 vccd1 _17234_/A sky130_fd_sc_hd__clkbuf_2
X_19071_ _19293_/CLK _19071_/D vssd1 vssd1 vccd1 vccd1 _19071_/Q sky130_fd_sc_hd__dfxtp_1
X_13495_ _19802_/Q vssd1 vssd1 vccd1 vccd1 _17120_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16283_ _16278_/A _16282_/C _13282_/A vssd1 vssd1 vccd1 vccd1 _16283_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_157_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15400__S _15406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18022_ _18020_/Y _18021_/X _18110_/S vssd1 vssd1 vccd1 vccd1 _18022_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ _15234_/A vssd1 vssd1 vccd1 vccd1 _19140_/D sky130_fd_sc_hd__clkbuf_1
X_12446_ _17223_/A _12470_/C _12445_/Y vssd1 vssd1 vccd1 vccd1 _12446_/X sky130_fd_sc_hd__o21a_1
XFILLER_173_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11737__A0 _19957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15165_ _19114_/Q vssd1 vssd1 vccd1 vccd1 _15166_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_153_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12377_ _12377_/A vssd1 vssd1 vccd1 vccd1 _12474_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14016__S _14024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16676__B1 _16667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output83_A _12336_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14116_ _18684_/Q _13685_/X _14120_/S vssd1 vssd1 vccd1 vccd1 _14117_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _11328_/A vssd1 vssd1 vccd1 vccd1 _11328_/Y sky130_fd_sc_hd__inv_2
X_15096_ _15118_/A vssd1 vssd1 vccd1 vccd1 _15105_/S sky130_fd_sc_hd__buf_2
X_19973_ _19978_/CLK _19973_/D vssd1 vssd1 vccd1 vccd1 _19973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18924_ _19480_/CLK _18924_/D vssd1 vssd1 vccd1 vccd1 _18924_/Q sky130_fd_sc_hd__dfxtp_1
X_14047_ _14047_/A vssd1 vssd1 vccd1 vccd1 _18654_/D sky130_fd_sc_hd__clkbuf_1
X_11259_ _18796_/Q _19131_/Q _11259_/S vssd1 vssd1 vccd1 vccd1 _11260_/B sky130_fd_sc_hd__mux2_1
XFILLER_68_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18855_ _19313_/CLK _18855_/D vssd1 vssd1 vccd1 vccd1 _18855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17806_ _18083_/A _17806_/B vssd1 vssd1 vccd1 vccd1 _17806_/X sky130_fd_sc_hd__or2_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18786_ _19411_/CLK _18786_/D vssd1 vssd1 vccd1 vccd1 _18786_/Q sky130_fd_sc_hd__dfxtp_1
X_15998_ _15998_/A vssd1 vssd1 vccd1 vccd1 _19422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17737_ _17571_/X _17584_/X _17760_/S vssd1 vssd1 vccd1 vccd1 _17737_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14949_ _14949_/A vssd1 vssd1 vccd1 vccd1 _19015_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_161_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19803_/CLK sky130_fd_sc_hd__clkbuf_16
X_17668_ _17668_/A _17721_/C vssd1 vssd1 vccd1 vccd1 _17754_/A sky130_fd_sc_hd__nor2_2
XFILLER_165_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19407_ _19407_/CLK _19407_/D vssd1 vssd1 vccd1 vccd1 _19407_/Q sky130_fd_sc_hd__dfxtp_1
X_16619_ _16629_/A _16619_/B _16619_/C vssd1 vssd1 vccd1 vccd1 _19647_/D sky130_fd_sc_hd__nor3_1
XANTENNA__13603__B _13603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17599_ _17690_/A vssd1 vssd1 vccd1 vccd1 _17923_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_176_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19873_/CLK sky130_fd_sc_hd__clkbuf_16
X_19338_ _19844_/CLK _19338_/D vssd1 vssd1 vccd1 vccd1 _19338_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_116_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19269_ _19272_/CLK _19269_/D vssd1 vssd1 vccd1 vccd1 _19269_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10874__S1 _10084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14715__A _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09809__A _09809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10626__S1 _10604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13765__S _13765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09924_ _18691_/Q _19186_/Q _09924_/S vssd1 vssd1 vccd1 vccd1 _09925_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_114_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19577_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_120_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16141__S _16145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20044_ _20044_/CLK _20044_/D vssd1 vssd1 vccd1 vccd1 _20044_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09544__A _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input7_A io_dbus_rdata[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _09855_/A vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__buf_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15980__S _15984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09786_ _09786_/A vssd1 vssd1 vccd1 vccd1 _09786_/Y sky130_fd_sc_hd__inv_2
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_129_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19042_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _10630_/A vssd1 vssd1 vccd1 vccd1 _10632_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17700__S _18109_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11967__A0 _19964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10561_ _10294_/A _10560_/X _10296_/A vssd1 vssd1 vccd1 vccd1 _10561_/X sky130_fd_sc_hd__a21o_1
XANTENNA__14625__A _14657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12300_ _17977_/B _12300_/B vssd1 vssd1 vccd1 vccd1 _12301_/B sky130_fd_sc_hd__and2_1
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17001__A _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13280_ input7/X _13172_/A _13175_/A vssd1 vssd1 vccd1 vccd1 _13292_/A sky130_fd_sc_hd__a21o_1
X_10492_ _10486_/A _10491_/X _09709_/A vssd1 vssd1 vccd1 vccd1 _10492_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11968__B _17412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ _12174_/A _12174_/B _12203_/A _12230_/Y vssd1 vssd1 vccd1 vccd1 _12232_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_135_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12162_ _12602_/A _12189_/A _12190_/A vssd1 vssd1 vccd1 vccd1 _12162_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_162_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11290__S1 _10978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__A1 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ _11113_/A vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_111_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16970_ _19749_/Q _16970_/B vssd1 vssd1 vccd1 vccd1 _16973_/B sky130_fd_sc_hd__nor2_1
X_12093_ _15760_/A _12091_/Y _12157_/C _12066_/B vssd1 vssd1 vccd1 vccd1 _12093_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15921_ _19388_/Q _15197_/X _15929_/S vssd1 vssd1 vccd1 vccd1 _15922_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11044_ _11216_/A _11043_/X _10056_/A vssd1 vssd1 vccd1 vccd1 _11044_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__15890__S _15890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18640_ _19491_/CLK _18640_/D vssd1 vssd1 vccd1 vccd1 _18640_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18280__C1 _17243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15852_ _15852_/A vssd1 vssd1 vccd1 vccd1 _19357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14803_ _14803_/A vssd1 vssd1 vccd1 vccd1 _18954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18571_ _19389_/CLK _18571_/D vssd1 vssd1 vccd1 vccd1 _18571_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output121_A _12657_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15783_ _15783_/A _18458_/Q vssd1 vssd1 vccd1 vccd1 _15783_/Y sky130_fd_sc_hd__nand2_1
X_12995_ _12995_/A vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17522_ _17538_/C _17721_/A _17668_/A vssd1 vssd1 vccd1 vccd1 _17919_/A sky130_fd_sc_hd__and3b_1
X_14734_ _14734_/A vssd1 vssd1 vccd1 vccd1 _18919_/D sky130_fd_sc_hd__clkbuf_1
X_11946_ _19520_/Q _12155_/B _15760_/A vssd1 vssd1 vccd1 vccd1 _11946_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19272_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17453_ _17899_/B _17973_/B _17465_/S vssd1 vssd1 vccd1 vccd1 _17453_/X sky130_fd_sc_hd__mux2_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _14665_/A vssd1 vssd1 vccd1 vccd1 _18891_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _11877_/A vssd1 vssd1 vccd1 vccd1 _13172_/A sky130_fd_sc_hd__buf_4
X_16404_ _13277_/X _19560_/Q _16404_/S vssd1 vssd1 vccd1 vccd1 _16405_/A sky130_fd_sc_hd__mux2_1
X_13616_ _13616_/A vssd1 vssd1 vccd1 vccd1 _18507_/D sky130_fd_sc_hd__clkbuf_1
X_10828_ _19107_/Q _18873_/Q _19555_/Q _19203_/Q _11372_/S _09515_/A vssd1 vssd1 vccd1
+ vccd1 _10828_/X sky130_fd_sc_hd__mux4_1
X_17384_ _17392_/C _17384_/B vssd1 vssd1 vccd1 vccd1 _17534_/B sky130_fd_sc_hd__nor2_2
XFILLER_60_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14596_ _14596_/A vssd1 vssd1 vccd1 vccd1 _14596_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19123_ _19313_/CLK _19123_/D vssd1 vssd1 vccd1 vccd1 _19123_/Q sky130_fd_sc_hd__dfxtp_1
X_16335_ _12127_/X _15799_/A _16300_/A vssd1 vssd1 vccd1 vccd1 _16335_/Y sky130_fd_sc_hd__o21ai_1
X_13547_ _19355_/Q _12864_/X _13099_/A _19545_/Q _13546_/X vssd1 vssd1 vccd1 vccd1
+ _13547_/X sky130_fd_sc_hd__a221o_1
XFILLER_146_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10759_ _18774_/Q _19045_/Q _19269_/Q _19013_/Q _11449_/S _10718_/A vssd1 vssd1 vccd1
+ vccd1 _10759_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19054_ _19504_/CLK _19054_/D vssd1 vssd1 vccd1 vccd1 _19054_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09629__A _11046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16266_ _16265_/A _16265_/C _16265_/B vssd1 vssd1 vccd1 vccd1 _16267_/B sky130_fd_sc_hd__o21ai_1
X_13478_ _19351_/Q _12759_/X _12758_/A _19541_/Q _13477_/X vssd1 vssd1 vccd1 vccd1
+ _13478_/X sky130_fd_sc_hd__a221o_1
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18005_ _12336_/A _17844_/X _18004_/X _17858_/X vssd1 vssd1 vccd1 vccd1 _18005_/X
+ sky130_fd_sc_hd__o211a_1
X_15217_ _19135_/Q _15215_/X _15229_/S vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__mux2_1
X_12429_ _12429_/A _12429_/B vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__nand2_2
X_16197_ _16197_/A vssd1 vssd1 vccd1 vccd1 _19511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_31_clock clkbuf_opt_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19305_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_126_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15148_ _15148_/A vssd1 vssd1 vccd1 vccd1 _19105_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14270__A _14281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19956_ _19956_/CLK _19956_/D vssd1 vssd1 vccd1 vccd1 _19956_/Q sky130_fd_sc_hd__dfxtp_2
X_15079_ _14599_/X _19073_/Q _15083_/S vssd1 vssd1 vccd1 vccd1 _15080_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18907_ _19495_/CLK _18907_/D vssd1 vssd1 vccd1 vccd1 _18907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_42_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_46_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19508_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19887_ _19888_/CLK _19887_/D vssd1 vssd1 vccd1 vccd1 _19887_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_132_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09640_ _18827_/Q vssd1 vssd1 vccd1 vccd1 _11280_/S sky130_fd_sc_hd__clkbuf_2
X_18838_ _19200_/CLK _18838_/D vssd1 vssd1 vccd1 vccd1 _18838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09571_ _18602_/Q _18863_/Q _18762_/Q _19097_/Q _09761_/S _09569_/A vssd1 vssd1 vccd1
+ vccd1 _09572_/B sky130_fd_sc_hd__mux4_1
XFILLER_83_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18827__D _18827_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18769_ _19490_/CLK _18769_/D vssd1 vssd1 vccd1 vccd1 _18769_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13614__A _13744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10973__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09539__A _10195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10385__C1 _09826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15276__A _15276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09907_ _18595_/Q _18856_/Q _18755_/Q _19090_/Q _10197_/S _09899_/X vssd1 vssd1 vccd1
+ vccd1 _09908_/B sky130_fd_sc_hd__mux4_1
XFILLER_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11024__S1 _10974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20027_ _20027_/CLK _20027_/D vssd1 vssd1 vccd1 vccd1 _20027_/Q sky130_fd_sc_hd__dfxtp_1
X_09838_ _09904_/S vssd1 vssd1 vccd1 vccd1 _10160_/S sky130_fd_sc_hd__buf_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09769_ _10166_/A _09769_/B vssd1 vssd1 vccd1 vccd1 _09769_/X sky130_fd_sc_hd__or2_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _17467_/A _11712_/C _11849_/C _11688_/A vssd1 vssd1 vccd1 vccd1 _11807_/A
+ sky130_fd_sc_hd__o31a_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12864_/A vssd1 vssd1 vccd1 vccd1 _12802_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ _12601_/A _09266_/B _11730_/X _17378_/A _09304_/A vssd1 vssd1 vccd1 vccd1
+ _12598_/B sky130_fd_sc_hd__o32a_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18419__A1_N _12475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _18819_/Q _14449_/X _14450_/S vssd1 vssd1 vccd1 vccd1 _14451_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10860__B1 _10056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11662_ _16208_/S vssd1 vssd1 vccd1 vccd1 _12444_/A sky130_fd_sc_hd__buf_2
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _19728_/Q vssd1 vssd1 vccd1 vccd1 _16923_/C sky130_fd_sc_hd__clkbuf_2
X_10613_ _10613_/A vssd1 vssd1 vccd1 vccd1 _11440_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11404__A2 _11393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ _11553_/X _11554_/Y _11555_/X _11556_/Y _11592_/X vssd1 vssd1 vccd1 vccd1
+ _11593_/X sky130_fd_sc_hd__a221o_1
X_14381_ _14381_/A vssd1 vssd1 vccd1 vccd1 _18797_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10883__A _11250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16120_ _13453_/X _19477_/Q _16128_/S vssd1 vssd1 vccd1 vccd1 _16121_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13332_ _18487_/Q _13331_/X _13358_/S vssd1 vssd1 vccd1 vccd1 _13333_/A sky130_fd_sc_hd__mux2_1
X_10544_ _10544_/A _10544_/B vssd1 vssd1 vccd1 vccd1 _10544_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14074__B _14074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16051_ _16051_/A vssd1 vssd1 vccd1 vccd1 _19446_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13157__A2 _13560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10475_ _19373_/Q _18987_/Q _19437_/Q _18556_/Q _10382_/X _10462_/X vssd1 vssd1 vccd1
+ vccd1 _10476_/B sky130_fd_sc_hd__mux4_1
X_13263_ _19720_/Q vssd1 vssd1 vccd1 vccd1 _16920_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_170_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15002_ _15059_/S vssd1 vssd1 vccd1 vccd1 _15011_/S sky130_fd_sc_hd__buf_2
X_12214_ _12214_/A vssd1 vssd1 vccd1 vccd1 _12314_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13194_ _13194_/A _13194_/B vssd1 vssd1 vccd1 vccd1 _15228_/A sky130_fd_sc_hd__and2_2
XFILLER_29_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12145_ _12145_/A vssd1 vssd1 vccd1 vccd1 _17884_/B sky130_fd_sc_hd__buf_2
X_19810_ _20018_/CLK _19810_/D vssd1 vssd1 vccd1 vccd1 _19810_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09781__B2 _19921_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16953_ _19745_/Q _16957_/B _19741_/Q _19740_/Q vssd1 vssd1 vccd1 vccd1 _16955_/B
+ sky130_fd_sc_hd__and4_1
X_19741_ _19745_/CLK _19741_/D vssd1 vssd1 vccd1 vccd1 _19741_/Q sky130_fd_sc_hd__dfxtp_1
X_12076_ _12076_/A vssd1 vssd1 vccd1 vccd1 _12076_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11015__S1 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15904_ _13453_/X _19381_/Q _15912_/S vssd1 vssd1 vccd1 vccd1 _15905_/A sky130_fd_sc_hd__mux2_1
X_11027_ _11027_/A vssd1 vssd1 vccd1 vccd1 _11027_/Y sky130_fd_sc_hd__inv_2
X_19672_ _19804_/CLK _19672_/D vssd1 vssd1 vccd1 vccd1 _19672_/Q sky130_fd_sc_hd__dfxtp_1
X_16884_ _16897_/A _16884_/B _16891_/D vssd1 vssd1 vccd1 vccd1 _19725_/D sky130_fd_sc_hd__nor3_1
XFILLER_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18623_ _19409_/CLK _18623_/D vssd1 vssd1 vccd1 vccd1 _18623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15835_ _15834_/X _19353_/Q _15835_/S vssd1 vssd1 vccd1 vccd1 _15836_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11653__S _11657_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15125__S _15127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18554_ _19305_/CLK _18554_/D vssd1 vssd1 vccd1 vccd1 _18554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _15765_/X _19342_/Q _15772_/S vssd1 vssd1 vccd1 vccd1 _15767_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13093__A1 _16219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ _18463_/Q _12973_/X _10139_/A _12976_/X vssd1 vssd1 vccd1 vccd1 _18463_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17503_/X _17802_/C _17508_/S vssd1 vssd1 vccd1 vccd1 _17505_/X sky130_fd_sc_hd__mux2_1
X_14717_ _14717_/A vssd1 vssd1 vccd1 vccd1 _18911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18485_ _19563_/CLK _18485_/D vssd1 vssd1 vccd1 vccd1 _18485_/Q sky130_fd_sc_hd__dfxtp_1
X_11929_ _11990_/A _11990_/C _12194_/A vssd1 vssd1 vccd1 vccd1 _11930_/B sky130_fd_sc_hd__o21ai_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15697_ _19899_/Q _15668_/X _16235_/A vssd1 vssd1 vccd1 vccd1 _15697_/X sky130_fd_sc_hd__a21o_1
XFILLER_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17436_ _17508_/S vssd1 vssd1 vccd1 vccd1 _17565_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14648_ _14647_/X _18886_/Q _14654_/S vssd1 vssd1 vccd1 vccd1 _14649_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17367_ _17373_/A _17367_/B vssd1 vssd1 vccd1 vccd1 _17368_/A sky130_fd_sc_hd__and2_1
XFILLER_159_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14579_ _14579_/A vssd1 vssd1 vccd1 vccd1 _18864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19106_ _19288_/CLK _19106_/D vssd1 vssd1 vccd1 vccd1 _19106_/Q sky130_fd_sc_hd__dfxtp_1
X_16318_ _15784_/X _16317_/X _16318_/S vssd1 vssd1 vccd1 vccd1 _16318_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17298_ _17217_/Y _19872_/Q _17302_/S vssd1 vssd1 vccd1 vccd1 _17299_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19037_ _19487_/CLK _19037_/D vssd1 vssd1 vccd1 vccd1 _19037_/Q sky130_fd_sc_hd__dfxtp_1
X_16249_ _16248_/A _16248_/C _13191_/A vssd1 vssd1 vccd1 vccd1 _16250_/B sky130_fd_sc_hd__o21ai_1
XFILLER_115_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11159__A1 _11082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput102 _12024_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[9] sky130_fd_sc_hd__buf_2
Xoutput113 _12649_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[13] sky130_fd_sc_hd__buf_2
Xoutput124 _12661_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[23] sky130_fd_sc_hd__buf_2
XFILLER_127_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput135 _12636_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[4] sky130_fd_sc_hd__buf_2
XFILLER_99_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput146 _12161_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[13] sky130_fd_sc_hd__buf_2
Xoutput157 _12424_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[23] sky130_fd_sc_hd__buf_2
XANTENNA__15096__A _15118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput168 _11893_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[4] sky130_fd_sc_hd__buf_2
XANTENNA__13609__A _14074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__B _12667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19939_ _19987_/CLK _19939_/D vssd1 vssd1 vccd1 vccd1 _19939_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11006__S1 _11236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11331__A1 _10024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18200__A _18268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__S0 _11451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09822__A _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _09623_/A vssd1 vssd1 vccd1 vccd1 _09623_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09554_ _11315_/A vssd1 vssd1 vccd1 vccd1 _11204_/A sky130_fd_sc_hd__buf_2
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14874__S _14878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09485_ _11473_/A vssd1 vssd1 vccd1 vccd1 _10840_/A sky130_fd_sc_hd__buf_2
XANTENNA__16655__A _16672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10907__S _11085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _10147_/A _10257_/X _10259_/X _09580_/A vssd1 vssd1 vccd1 vccd1 _10260_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11245__S1 _11115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _10184_/Y _10186_/Y _10188_/Y _10190_/Y _09719_/X vssd1 vssd1 vccd1 vccd1
+ _10191_/X sky130_fd_sc_hd__o221a_1
XANTENNA__14114__S _14120_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13953__S _13961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13950_ _18612_/Q _13651_/X _13950_/S vssd1 vssd1 vccd1 vccd1 _13951_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10756__S0 _09647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ _18460_/Q _12901_/B vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__or2_1
XFILLER_59_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13881_ _13783_/X _18581_/Q _13889_/S vssd1 vssd1 vccd1 vccd1 _13882_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15620_ _14618_/X _19303_/Q _15622_/S vssd1 vssd1 vccd1 vccd1 _15621_/A sky130_fd_sc_hd__mux2_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _13116_/A vssd1 vssd1 vccd1 vccd1 _12832_/X sky130_fd_sc_hd__buf_2
XFILLER_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15551_/A vssd1 vssd1 vccd1 vccd1 _19272_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14784__S _14786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12763_ _19755_/Q _12692_/X _12762_/X _12714_/X vssd1 vssd1 vccd1 vccd1 _12763_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14502_/A _15589_/B vssd1 vssd1 vccd1 vccd1 _14559_/A sky130_fd_sc_hd__or2_4
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _09328_/D _19989_/Q _18273_/S vssd1 vssd1 vccd1 vccd1 _18271_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11764_/A _11764_/B _11764_/C vssd1 vssd1 vccd1 vccd1 _11717_/A sky130_fd_sc_hd__o21ai_1
X_15482_ _15482_/A vssd1 vssd1 vccd1 vccd1 _19241_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _13205_/A vssd1 vssd1 vccd1 vccd1 _12695_/A sky130_fd_sc_hd__buf_2
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17221_ _19840_/Q _17226_/B vssd1 vssd1 vccd1 vccd1 _17221_/X sky130_fd_sc_hd__or2_1
XFILLER_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14637_/A vssd1 vssd1 vccd1 vccd1 _14433_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11645_ _11675_/A _11645_/B vssd1 vssd1 vccd1 vccd1 _17337_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17152_ _17152_/A vssd1 vssd1 vccd1 vccd1 _17152_/Y sky130_fd_sc_hd__inv_2
Xinput15 io_dbus_rdata[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_4
X_14364_ _14364_/A vssd1 vssd1 vccd1 vccd1 _18792_/D sky130_fd_sc_hd__clkbuf_1
Xinput26 io_dbus_rdata[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_4
X_11576_ _11570_/B _11573_/Y _11574_/Y _11575_/Y vssd1 vssd1 vccd1 vccd1 _11576_/Y
+ sky130_fd_sc_hd__a22oi_1
Xinput37 io_ibus_inst[12] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_2
XFILLER_168_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16103_ _16103_/A vssd1 vssd1 vccd1 vccd1 _19469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput48 io_ibus_inst[22] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_2
XFILLER_128_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput59 io_ibus_inst[3] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13315_ _13335_/C _13315_/B vssd1 vssd1 vccd1 vccd1 _13315_/Y sky130_fd_sc_hd__nor2_1
X_10527_ _10521_/A _10524_/X _10526_/X _10307_/A vssd1 vssd1 vccd1 vccd1 _10527_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17083_ _17108_/A _17087_/C vssd1 vssd1 vccd1 vccd1 _17083_/Y sky130_fd_sc_hd__nor2_1
X_14295_ _14295_/A vssd1 vssd1 vccd1 vccd1 _18762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16034_ _13357_/X _19439_/Q _16034_/S vssd1 vssd1 vccd1 vccd1 _16035_/A sky130_fd_sc_hd__mux2_1
X_10458_ _10459_/A _12655_/B vssd1 vssd1 vccd1 vccd1 _10460_/A sky130_fd_sc_hd__and2_1
XFILLER_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13246_ _19863_/Q _12699_/A _13205_/X _19830_/Q vssd1 vssd1 vccd1 vccd1 _13246_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10389_ _10448_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _10389_/Y sky130_fd_sc_hd__nor2_1
X_13177_ _13060_/X _13167_/X _13171_/X _13176_/X vssd1 vssd1 vccd1 vccd1 _15225_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14024__S _14024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15827__A1 _18465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12128_ _19829_/Q vssd1 vssd1 vccd1 vccd1 _17187_/A sky130_fd_sc_hd__buf_2
X_17985_ _17985_/A _17985_/B vssd1 vssd1 vccd1 vccd1 _17985_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14959__S _14961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13863__S _13867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13302__A2 _19909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19724_ _19726_/CLK _19724_/D vssd1 vssd1 vccd1 vccd1 _19724_/Q sky130_fd_sc_hd__dfxtp_1
X_16936_ _19741_/Q _16936_/B vssd1 vssd1 vccd1 vccd1 _16939_/B sky130_fd_sc_hd__or2_1
XFILLER_42_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12059_ _12086_/A _12086_/C vssd1 vssd1 vccd1 vccd1 _12059_/X sky130_fd_sc_hd__xor2_1
XFILLER_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11313__A1 _10949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__B1 _19605_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16867_ _16920_/B _16920_/C _16866_/X vssd1 vssd1 vccd1 vccd1 _19720_/D sky130_fd_sc_hd__o21ba_1
X_19655_ _19789_/CLK _19655_/D vssd1 vssd1 vccd1 vccd1 _19655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15818_ _15818_/A vssd1 vssd1 vccd1 vccd1 _15818_/X sky130_fd_sc_hd__clkbuf_4
X_18606_ _19487_/CLK _18606_/D vssd1 vssd1 vccd1 vccd1 _18606_/Q sky130_fd_sc_hd__dfxtp_1
X_19586_ _19594_/CLK _19586_/D vssd1 vssd1 vccd1 vccd1 _19586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16798_ _19704_/Q _16798_/B vssd1 vssd1 vccd1 vccd1 _16799_/B sky130_fd_sc_hd__and2_1
XFILLER_53_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18537_ _19204_/CLK _18537_/D vssd1 vssd1 vccd1 vccd1 _18537_/Q sky130_fd_sc_hd__dfxtp_1
X_15749_ _15811_/A _18452_/Q vssd1 vssd1 vccd1 vccd1 _15749_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14694__S _14702_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09270_ _09303_/A _11684_/A _09301_/A _09298_/A vssd1 vssd1 vccd1 vccd1 _09277_/C
+ sky130_fd_sc_hd__o211a_1
X_18468_ _19938_/CLK _18468_/D vssd1 vssd1 vccd1 vccd1 _18468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17419_ _17419_/A vssd1 vssd1 vccd1 vccd1 _17450_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18399_ _18308_/A _12880_/A _14481_/X _18398_/Y vssd1 vssd1 vccd1 vccd1 _18400_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11227__S1 _09659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17245__S _17245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16491__A1 _19606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09606_ _09591_/X _09593_/X _09595_/X _09597_/X _09605_/X vssd1 vssd1 vccd1 vccd1
+ _09606_/X sky130_fd_sc_hd__a221o_1
XFILLER_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09537_ _10417_/S vssd1 vssd1 vccd1 vccd1 _10416_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_58_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ _17323_/B vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_164_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ _18338_/A _12702_/A _12701_/A _09391_/B _12797_/B vssd1 vssd1 vccd1 vccd1
+ _09399_/X sky130_fd_sc_hd__a2111o_1
XFILLER_156_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11430_ _10734_/A _11429_/X _09989_/A vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__a21o_1
XFILLER_165_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13948__S _13950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11361_ _19369_/Q _18983_/Q _19433_/Q _18552_/Q _10614_/X _11371_/A vssd1 vssd1 vccd1
+ vccd1 _11362_/B sky130_fd_sc_hd__mux4_1
XFILLER_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10312_ _10312_/A vssd1 vssd1 vccd1 vccd1 _10312_/X sky130_fd_sc_hd__buf_2
XFILLER_137_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13100_ _19855_/Q _12992_/X _12695_/A _19822_/Q vssd1 vssd1 vccd1 vccd1 _13100_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11292_ _19485_/Q _18897_/Q _18934_/Q _18508_/Q _10977_/A _10006_/A vssd1 vssd1 vccd1
+ vccd1 _11292_/X sky130_fd_sc_hd__mux4_1
X_14080_ _14080_/A vssd1 vssd1 vccd1 vccd1 _18667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10243_ _10243_/A _10243_/B vssd1 vssd1 vccd1 vccd1 _10243_/X sky130_fd_sc_hd__or2_1
XFILLER_106_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13031_ _19926_/Q _13030_/X _13554_/S vssd1 vssd1 vccd1 vccd1 _13031_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input45_A io_ibus_inst[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ _10174_/A vssd1 vssd1 vccd1 vccd1 _10174_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17770_ _17768_/Y _17769_/X _18110_/S vssd1 vssd1 vccd1 vccd1 _17770_/X sky130_fd_sc_hd__mux2_1
X_14982_ _14982_/A vssd1 vssd1 vccd1 vccd1 _19030_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10729__S0 _10608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_89_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16721_ _16731_/A _16727_/C vssd1 vssd1 vccd1 vccd1 _16721_/Y sky130_fd_sc_hd__nor2_1
X_13933_ _18604_/Q _13618_/X _13939_/S vssd1 vssd1 vccd1 vccd1 _13934_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19440_ _19566_/CLK _19440_/D vssd1 vssd1 vccd1 vccd1 _19440_/Q sky130_fd_sc_hd__dfxtp_1
X_16652_ _16653_/B _16653_/C _16651_/Y vssd1 vssd1 vccd1 vccd1 _19658_/D sky130_fd_sc_hd__o21a_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13864_ _13864_/A vssd1 vssd1 vccd1 vccd1 _18573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15603_ _14592_/X _19295_/Q _15611_/S vssd1 vssd1 vccd1 vccd1 _15604_/A sky130_fd_sc_hd__mux2_1
X_19371_ _19500_/CLK _19371_/D vssd1 vssd1 vccd1 vccd1 _19371_/Q sky130_fd_sc_hd__dfxtp_1
X_12815_ _13578_/A _18440_/Q vssd1 vssd1 vccd1 vccd1 _12815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16583_ _16629_/A _16583_/B _16584_/B vssd1 vssd1 vccd1 vccd1 _19634_/D sky130_fd_sc_hd__nor3_1
XFILLER_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13795_ _13795_/A vssd1 vssd1 vccd1 vccd1 _18552_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11154__S0 _11224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18322_ _20008_/Q _18310_/X _18321_/X _18317_/X vssd1 vssd1 vccd1 vccd1 _20008_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _15534_/A vssd1 vssd1 vccd1 vccd1 _19264_/D sky130_fd_sc_hd__clkbuf_1
X_12746_ _12686_/Y _12741_/X _12745_/X vssd1 vssd1 vccd1 vccd1 _19809_/D sky130_fd_sc_hd__o21a_1
XFILLER_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17734__A1 _11864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12271__A2 _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _19981_/Q _19602_/Q _18253_/S vssd1 vssd1 vccd1 vccd1 _18254_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15465_ _19234_/Q _15225_/X _15467_/S vssd1 vssd1 vccd1 vccd1 _15466_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12328__A _12328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12677_ _12677_/A vssd1 vssd1 vccd1 vccd1 _17140_/C sky130_fd_sc_hd__buf_2
X_17204_ _12772_/B _17197_/X _17203_/X _17201_/X vssd1 vssd1 vccd1 vccd1 _19834_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11232__A _19896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14416_ _14416_/A vssd1 vssd1 vccd1 vccd1 _18808_/D sky130_fd_sc_hd__clkbuf_1
X_18184_ _19950_/Q _19982_/Q _18192_/S vssd1 vssd1 vccd1 vccd1 _18185_/A sky130_fd_sc_hd__mux2_1
X_11628_ _11623_/Y _17342_/B _11625_/X _12596_/B vssd1 vssd1 vccd1 vccd1 _11628_/X
+ sky130_fd_sc_hd__a31o_1
X_15396_ _15396_/A vssd1 vssd1 vccd1 vccd1 _19203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17498__A0 _12480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17135_ _19812_/Q _12880_/X _17134_/X _16480_/X vssd1 vssd1 vccd1 vccd1 _19812_/D
+ sky130_fd_sc_hd__o211a_1
X_14347_ _14347_/A vssd1 vssd1 vccd1 vccd1 _18784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11559_ _11563_/A _11560_/C _11560_/A vssd1 vssd1 vccd1 vccd1 _11559_/X sky130_fd_sc_hd__a21o_1
XFILLER_143_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17066_ _17066_/A _17070_/C vssd1 vssd1 vccd1 vccd1 _17066_/Y sky130_fd_sc_hd__nor2_1
X_14278_ _14278_/A vssd1 vssd1 vccd1 vccd1 _18754_/D sky130_fd_sc_hd__clkbuf_1
X_16017_ _13230_/X _19431_/Q _16023_/S vssd1 vssd1 vccd1 vccd1 _16018_/A sky130_fd_sc_hd__mux2_1
X_13229_ _11656_/X _13227_/X _13228_/X vssd1 vssd1 vccd1 vccd1 _15235_/A sky130_fd_sc_hd__o21a_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14689__S _14691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15374__A _15430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17968_ _17619_/X _17912_/Y _17967_/X vssd1 vssd1 vccd1 vccd1 _17968_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19707_ _19877_/CLK _19707_/D vssd1 vssd1 vccd1 vccd1 _19707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16919_ _16919_/A _16919_/B _16955_/A vssd1 vssd1 vccd1 vccd1 _19737_/D sky130_fd_sc_hd__nor3_1
XANTENNA__17422__A0 _17749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17899_ _18033_/A _17899_/B vssd1 vssd1 vccd1 vccd1 _17899_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19638_ _19769_/CLK _19638_/D vssd1 vssd1 vccd1 vccd1 _19638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16917__B _16930_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19569_ _19569_/CLK _19569_/D vssd1 vssd1 vccd1 vccd1 _19569_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16409__S _16415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11145__S0 _11030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ _11615_/A _11699_/A _09321_/X vssd1 vssd1 vccd1 vccd1 _09322_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09253_ _09303_/A _11724_/D _09214_/C _12594_/C vssd1 vssd1 vccd1 vccd1 _11624_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_09184_ _11680_/C _11646_/C vssd1 vssd1 vccd1 vccd1 _17331_/A sky130_fd_sc_hd__nand2_1
XFILLER_159_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14453__A _14453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11773__A1 _19813_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13069__A _15209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_90_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__A _15198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17413__A0 _17792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10930_ _18643_/Q _19234_/Q _19396_/Q _18611_/Q _11493_/S _09660_/A vssd1 vssd1 vccd1
+ vccd1 _10930_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10861_ _18644_/Q _19235_/Q _19397_/Q _18612_/Q _10777_/A _10010_/X vssd1 vssd1 vccd1
+ vccd1 _10862_/B sky130_fd_sc_hd__mux4_2
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14628__A _14628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11136__S0 _11035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12600_ _12600_/A vssd1 vssd1 vccd1 vccd1 _17323_/A sky130_fd_sc_hd__buf_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17004__A _17046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ _13580_/A vssd1 vssd1 vccd1 vccd1 _13580_/X sky130_fd_sc_hd__buf_2
X_10792_ _10792_/A _10792_/B vssd1 vssd1 vccd1 vccd1 _10792_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13450__A1 _13449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12531_/A _18090_/B vssd1 vssd1 vccd1 vccd1 _12532_/B sky130_fd_sc_hd__or2_1
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10367__S _10367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _15250_/A vssd1 vssd1 vccd1 vccd1 _19145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12462_ _12482_/B _12462_/B vssd1 vssd1 vccd1 vccd1 _12463_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11439__S1 _10691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14201_ _13819_/X _18720_/Q _14207_/S vssd1 vssd1 vccd1 vccd1 _14202_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13678__S _13694_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ _11562_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _11413_/X sky130_fd_sc_hd__and2_1
XANTENNA__11987__A _11987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15181_ _19122_/Q vssd1 vssd1 vccd1 vccd1 _15182_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__16054__S _16056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10891__A _18965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ _19600_/Q _12393_/B vssd1 vssd1 vccd1 vccd1 _12438_/C sky130_fd_sc_hd__and2_1
XFILLER_137_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14132_ _14132_/A vssd1 vssd1 vccd1 vccd1 _18691_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12961__B1 _10672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ _10986_/A _11343_/X _10920_/A vssd1 vssd1 vccd1 vccd1 _11344_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15893__S _15901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14063_ _14063_/A vssd1 vssd1 vccd1 vccd1 _18661_/D sky130_fd_sc_hd__clkbuf_1
X_18940_ _19042_/CLK _18940_/D vssd1 vssd1 vccd1 vccd1 _18940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11275_ _10941_/X _11272_/X _11274_/X _09574_/A vssd1 vssd1 vccd1 vccd1 _11275_/X
+ sky130_fd_sc_hd__o211a_1
X_13014_ _14844_/C vssd1 vssd1 vccd1 vccd1 _18295_/A sky130_fd_sc_hd__clkinv_4
X_10226_ _10233_/A _10225_/X _09891_/X vssd1 vssd1 vccd1 vccd1 _10226_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_output151_A _12297_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18871_ _19201_/CLK _18871_/D vssd1 vssd1 vccd1 vccd1 _18871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10157_ _10209_/A _10154_/X _10156_/X _09826_/X vssd1 vssd1 vccd1 vccd1 _10157_/X
+ sky130_fd_sc_hd__o211a_1
X_17822_ _17816_/X _17818_/Y _17821_/X vssd1 vssd1 vccd1 vccd1 _17822_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14302__S _14308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14965_ _14965_/A vssd1 vssd1 vccd1 vccd1 _19022_/D sky130_fd_sc_hd__clkbuf_1
X_10088_ _10817_/A _10088_/B vssd1 vssd1 vccd1 vccd1 _10088_/X sky130_fd_sc_hd__or2_1
XFILLER_47_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17753_ _17560_/X _17743_/X _17752_/X _17598_/X vssd1 vssd1 vccd1 vccd1 _17753_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16207__A1 _11890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13916_ _13835_/X _18597_/Q _13922_/S vssd1 vssd1 vccd1 vccd1 _13917_/A sky130_fd_sc_hd__mux2_1
X_16704_ _19799_/Q _19801_/Q _19800_/Q _17107_/A vssd1 vssd1 vccd1 vccd1 _17115_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17684_ _17682_/X _17683_/X _17759_/S vssd1 vssd1 vccd1 vccd1 _17684_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14896_ _14647_/X _18992_/Q _14900_/S vssd1 vssd1 vccd1 vccd1 _14897_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17955__A1 _12234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16635_ _16635_/A vssd1 vssd1 vccd1 vccd1 _16672_/A sky130_fd_sc_hd__buf_2
X_19423_ _19455_/CLK _19423_/D vssd1 vssd1 vccd1 vccd1 _19423_/Q sky130_fd_sc_hd__dfxtp_1
X_13847_ _14672_/A vssd1 vssd1 vccd1 vccd1 _13847_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19354_ _19762_/CLK _19354_/D vssd1 vssd1 vccd1 vccd1 _19354_/Q sky130_fd_sc_hd__dfxtp_1
X_16566_ _19629_/Q _16566_/B vssd1 vssd1 vccd1 vccd1 _16572_/C sky130_fd_sc_hd__and2_1
XFILLER_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13778_ _13777_/X _18547_/Q _13781_/S vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15517_ _15918_/B _15517_/B vssd1 vssd1 vccd1 vccd1 _15574_/A sky130_fd_sc_hd__nor2_4
X_18305_ _18323_/A vssd1 vssd1 vccd1 vccd1 _18331_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_19285_ _19285_/CLK _19285_/D vssd1 vssd1 vccd1 vccd1 _19285_/Q sky130_fd_sc_hd__dfxtp_1
X_12729_ _13117_/A vssd1 vssd1 vccd1 vccd1 _12729_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16497_ _19649_/Q _19651_/Q _19650_/Q _16620_/A vssd1 vssd1 vccd1 vccd1 _16630_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_148_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18236_ _19973_/Q _16474_/A _18242_/S vssd1 vssd1 vccd1 vccd1 _18237_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15448_ _19226_/Q _15197_/X _15456_/S vssd1 vssd1 vccd1 vccd1 _15449_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18167_ _18167_/A vssd1 vssd1 vccd1 vccd1 _19942_/D sky130_fd_sc_hd__clkbuf_1
X_15379_ _15379_/A vssd1 vssd1 vccd1 vccd1 _19195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18132__A1 _19959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11755__A1 _18316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17118_ _17120_/B _17120_/C _17101_/X vssd1 vssd1 vccd1 vccd1 _17118_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12952__B1 _11355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18098_ _18118_/A _18098_/B vssd1 vssd1 vccd1 vccd1 _18098_/X sky130_fd_sc_hd__or2_1
X_09940_ _10283_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _09940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17049_ _19777_/Q _17046_/B _17048_/Y vssd1 vssd1 vccd1 vccd1 _19777_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17891__B1 _12117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09871_ _10279_/A vssd1 vssd1 vccd1 vccd1 _10229_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_112_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09581__C1 _09580_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13617__A _15203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14212__S _14218_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16139__S _16145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10246__A1 _10368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15978__S _15984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ _11627_/C _12595_/C _11724_/D vssd1 vssd1 vccd1 vccd1 _17393_/B sky130_fd_sc_hd__or3_1
XANTENNA__09731__S0 _09726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16663__A _16672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_37_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09236_ _09275_/C _11730_/B _11730_/C vssd1 vssd1 vccd1 vccd1 _11729_/A sky130_fd_sc_hd__or3_2
XFILLER_142_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16214__A_N _16206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15279__A _15279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09277__A _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11210__A3 _11209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17494__A _17675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11060_ _18800_/Q _19135_/Q _11114_/S vssd1 vssd1 vccd1 vccd1 _11061_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10706__C1 _11383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10011_ _19124_/Q _18890_/Q _19572_/Q _19220_/Q _10777_/A _10010_/X vssd1 vssd1 vccd1
+ vccd1 _10012_/B sky130_fd_sc_hd__mux4_1
XFILLER_103_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13961__S _13961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ _18927_/Q _14471_/X _14750_/S vssd1 vssd1 vccd1 vccd1 _14751_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11962_ _11962_/A vssd1 vssd1 vccd1 vccd1 _12039_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11277__A3 _11276_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ _15267_/A vssd1 vssd1 vccd1 vccd1 _14644_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09740__A _09740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ _11035_/A vssd1 vssd1 vccd1 vccd1 _11026_/S sky130_fd_sc_hd__buf_4
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14681_ _14737_/A vssd1 vssd1 vccd1 vccd1 _14750_/S sky130_fd_sc_hd__buf_6
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11893_ _11893_/A vssd1 vssd1 vccd1 vccd1 _11893_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11109__S0 _11000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16420_ _13393_/X _19567_/Q _16426_/S vssd1 vssd1 vccd1 vccd1 _16421_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13632_ _13632_/A vssd1 vssd1 vccd1 vccd1 _18511_/D sky130_fd_sc_hd__clkbuf_1
X_10844_ _09613_/A _10834_/X _10843_/X _09996_/X _19902_/Q vssd1 vssd1 vccd1 vccd1
+ _10869_/A sky130_fd_sc_hd__a32o_4
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15888__S _15890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16351_ _19541_/Q _16300_/X _16349_/Y _16350_/X vssd1 vssd1 vccd1 vccd1 _19541_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13563_ _12420_/A _13562_/Y _12857_/A vssd1 vssd1 vccd1 vccd1 _13563_/Y sky130_fd_sc_hd__o21ai_1
X_10775_ _19903_/Q vssd1 vssd1 vccd1 vccd1 _10775_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_13_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15302_ _15358_/A vssd1 vssd1 vccd1 vccd1 _15371_/S sky130_fd_sc_hd__buf_6
X_19070_ _19292_/CLK _19070_/D vssd1 vssd1 vccd1 vccd1 _19070_/Q sky130_fd_sc_hd__dfxtp_1
X_12514_ _19541_/Q _12122_/X _12262_/X _12513_/X _12123_/X vssd1 vssd1 vccd1 vccd1
+ _12514_/X sky130_fd_sc_hd__o221a_1
X_16282_ _19939_/Q _19940_/Q _16282_/C vssd1 vssd1 vccd1 vccd1 _16290_/B sky130_fd_sc_hd__or3_1
X_13494_ _19670_/Q vssd1 vssd1 vccd1 vccd1 _16689_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18021_ _18023_/A _18023_/B _18088_/S vssd1 vssd1 vccd1 vccd1 _18021_/X sky130_fd_sc_hd__mux2_1
X_15233_ _19140_/Q _15231_/X _15245_/S vssd1 vssd1 vccd1 vccd1 _15234_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12445_ _17223_/A _12470_/C _12444_/X vssd1 vssd1 vccd1 vccd1 _12445_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_172_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12606__A _12606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11737__A1 _11324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15164_ _15164_/A vssd1 vssd1 vccd1 vccd1 _19113_/D sky130_fd_sc_hd__clkbuf_1
X_12376_ _12376_/A vssd1 vssd1 vccd1 vccd1 _12473_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__10945__C1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14115_ _14115_/A vssd1 vssd1 vccd1 vccd1 _18683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11327_ _18667_/Q _19162_/Q _11327_/S vssd1 vssd1 vccd1 vccd1 _11328_/A sky130_fd_sc_hd__mux2_1
X_15095_ _15095_/A vssd1 vssd1 vccd1 vccd1 _19080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19972_ _19978_/CLK _19972_/D vssd1 vssd1 vccd1 vccd1 _19972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output76_A _12175_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18923_ _19092_/CLK _18923_/D vssd1 vssd1 vccd1 vccd1 _18923_/Q sky130_fd_sc_hd__dfxtp_1
X_14046_ _18654_/Q _13693_/X _14046_/S vssd1 vssd1 vccd1 vccd1 _14047_/A sky130_fd_sc_hd__mux2_1
X_11258_ _18668_/Q _19163_/Q _11306_/S vssd1 vssd1 vccd1 vccd1 _11258_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12162__A1 _12602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10209_ _10209_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10209_/X sky130_fd_sc_hd__or2_1
XANTENNA__10560__S _10560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18854_ _19476_/CLK _18854_/D vssd1 vssd1 vccd1 vccd1 _18854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11189_ _18669_/Q _19164_/Q _11191_/S vssd1 vssd1 vccd1 vccd1 _11190_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17805_ _17801_/X _17804_/X _17805_/S vssd1 vssd1 vccd1 vccd1 _17806_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17851__B _17853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18785_ _19411_/CLK _18785_/D vssd1 vssd1 vccd1 vccd1 _18785_/Q sky130_fd_sc_hd__dfxtp_1
X_15997_ _13056_/X _19422_/Q _16001_/S vssd1 vssd1 vccd1 vccd1 _15998_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14948_ _19015_/Q _14414_/X _14950_/S vssd1 vssd1 vccd1 vccd1 _14949_/A sky130_fd_sc_hd__mux2_1
X_17736_ _17574_/X _17563_/X _17759_/S vssd1 vssd1 vccd1 vccd1 _17736_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09650__A _10496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14879_ _14879_/A vssd1 vssd1 vccd1 vccd1 _18984_/D sky130_fd_sc_hd__clkbuf_1
X_17667_ _17667_/A _17667_/B vssd1 vssd1 vccd1 vccd1 _17667_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13172__A _13172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19406_ _19406_/CLK _19406_/D vssd1 vssd1 vccd1 vccd1 _19406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16618_ _16617_/B _16617_/C _19647_/Q vssd1 vssd1 vccd1 vccd1 _16619_/C sky130_fd_sc_hd__a21oi_1
X_17598_ _17953_/A vssd1 vssd1 vccd1 vccd1 _17598_/X sky130_fd_sc_hd__clkbuf_2
X_16549_ _19623_/Q _19622_/Q _19621_/Q _16549_/D vssd1 vssd1 vccd1 vccd1 _16555_/C
+ sky130_fd_sc_hd__and4_1
X_19337_ _19783_/CLK _19337_/D vssd1 vssd1 vccd1 vccd1 _19337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16364__A0 _15839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19268_ _19268_/CLK _19268_/D vssd1 vssd1 vccd1 vccd1 _19268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ _18219_/A vssd1 vssd1 vccd1 vccd1 _19965_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10735__S _10735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19199_ _19201_/CLK _19199_/D vssd1 vssd1 vccd1 vccd1 _19199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13111__S _13196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10087__S0 _11483_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16422__S _16426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09923_ _10279_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09923_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13350__A0 _19912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20043_ _20052_/CLK _20043_/D vssd1 vssd1 vccd1 vccd1 _20043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09854_ _10396_/A vssd1 vssd1 vccd1 vccd1 _09855_/A sky130_fd_sc_hd__buf_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__A1 _12097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _18695_/Q _19190_/Q _09787_/S vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11339__S0 _11030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10467__A1 _10294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__S0 _10777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11967__A1 _10961_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__S0 _11384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ _18682_/Q _19177_/Q _10560_/S vssd1 vssd1 vccd1 vccd1 _10560_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09219_ _19888_/Q _09349_/B vssd1 vssd1 vccd1 vccd1 _09325_/A sky130_fd_sc_hd__or2_4
XFILLER_154_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10491_ _19469_/Q _19307_/Q _18716_/Q _18486_/Q _10390_/S _10333_/A vssd1 vssd1 vccd1
+ vccd1 _10491_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11330__A _11330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12230_ _12170_/A _12201_/A _12229_/Y vssd1 vssd1 vccd1 vccd1 _12230_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12161_ _12161_/A vssd1 vssd1 vccd1 vccd1 _12161_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__14641__A _14657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11112_ _18966_/Q vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__clkbuf_2
X_12092_ _19828_/Q _19827_/Q _12092_/C vssd1 vssd1 vccd1 vccd1 _12157_/C sky130_fd_sc_hd__and3_2
XFILLER_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15920_ _15988_/S vssd1 vssd1 vccd1 vccd1 _15929_/S sky130_fd_sc_hd__clkbuf_4
X_11043_ _19490_/Q _18902_/Q _18939_/Q _18513_/Q _10903_/A _10974_/X vssd1 vssd1 vccd1
+ vccd1 _11043_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12161__A _12161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15851_ _13033_/X _19357_/Q _15857_/S vssd1 vssd1 vccd1 vccd1 _15852_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14802_ _18954_/Q _14440_/X _14808_/S vssd1 vssd1 vccd1 vccd1 _14803_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18570_ _19576_/CLK _18570_/D vssd1 vssd1 vccd1 vccd1 _18570_/Q sky130_fd_sc_hd__dfxtp_1
X_15782_ _18458_/Q _15782_/B vssd1 vssd1 vccd1 vccd1 _15782_/X sky130_fd_sc_hd__or2_1
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12994_ _18502_/Q _13546_/B _12707_/X _19324_/Q _12993_/X vssd1 vssd1 vccd1 vccd1
+ _12994_/X sky130_fd_sc_hd__a221o_1
XFILLER_29_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14733_ _18919_/Q _14446_/X _14735_/S vssd1 vssd1 vccd1 vccd1 _14734_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17521_ _18054_/A vssd1 vssd1 vccd1 vccd1 _17521_/X sky130_fd_sc_hd__clkbuf_2
X_11945_ _12032_/A vssd1 vssd1 vccd1 vccd1 _15760_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output114_A _12650_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17452_/A vssd1 vssd1 vccd1 vccd1 _17973_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _14663_/X _18891_/Q _14670_/S vssd1 vssd1 vccd1 vccd1 _14665_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11876_ _19820_/Q _11842_/B _11843_/X vssd1 vssd1 vccd1 vccd1 _11917_/A sky130_fd_sc_hd__a21bo_1
XFILLER_60_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16403_ _16403_/A vssd1 vssd1 vccd1 vccd1 _19559_/D sky130_fd_sc_hd__clkbuf_1
X_13615_ _18507_/Q _13608_/X _13631_/S vssd1 vssd1 vccd1 vccd1 _13616_/A sky130_fd_sc_hd__mux2_1
X_10827_ _09985_/X _10826_/X _10606_/A vssd1 vssd1 vccd1 vccd1 _10827_/X sky130_fd_sc_hd__a21o_1
X_17383_ _09304_/A _09266_/X _12641_/A _17382_/X _17325_/X vssd1 vssd1 vccd1 vccd1
+ _17384_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14595_ _14595_/A vssd1 vssd1 vccd1 vccd1 _18869_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15411__S _15417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19122_ _19508_/CLK _19122_/D vssd1 vssd1 vccd1 vccd1 _19122_/Q sky130_fd_sc_hd__dfxtp_1
X_16334_ _16338_/B _16333_/Y _16303_/X vssd1 vssd1 vccd1 vccd1 _16334_/Y sky130_fd_sc_hd__a21oi_1
X_13546_ _18506_/Q _13546_/B vssd1 vssd1 vccd1 vccd1 _13546_/X sky130_fd_sc_hd__and2_1
X_10758_ _18582_/Q _18843_/Q _18742_/Q _19077_/Q _09647_/A _10030_/A vssd1 vssd1 vccd1
+ vccd1 _10758_/X sky130_fd_sc_hd__mux4_2
XFILLER_13_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19053_ _19053_/CLK _19053_/D vssd1 vssd1 vccd1 vccd1 _19053_/Q sky130_fd_sc_hd__dfxtp_1
X_16265_ _16265_/A _16265_/B _16265_/C vssd1 vssd1 vccd1 vccd1 _16273_/B sky130_fd_sc_hd__or3_1
XANTENNA__14027__S _14035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13477_ _19877_/Q _12699_/A _13343_/X _19844_/Q vssd1 vssd1 vccd1 vccd1 _13477_/X
+ sky130_fd_sc_hd__a22o_1
X_10689_ _11362_/A _10689_/B vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__or2_1
X_15216_ _15299_/S vssd1 vssd1 vccd1 vccd1 _15229_/S sky130_fd_sc_hd__buf_2
X_18004_ _17619_/X _17862_/Y _18003_/X vssd1 vssd1 vccd1 vccd1 _18004_/X sky130_fd_sc_hd__a21o_1
XFILLER_173_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12428_ _12428_/A _18033_/B vssd1 vssd1 vccd1 vccd1 _12429_/B sky130_fd_sc_hd__nand2_1
X_16196_ _19511_/Q _14663_/A _16200_/S vssd1 vssd1 vccd1 vccd1 _16197_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15147_ _19105_/Q vssd1 vssd1 vccd1 vccd1 _15148_/A sky130_fd_sc_hd__clkbuf_1
X_12359_ _12390_/A _12359_/B vssd1 vssd1 vccd1 vccd1 _12361_/A sky130_fd_sc_hd__nand2_2
XFILLER_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19955_ _19987_/CLK _19955_/D vssd1 vssd1 vccd1 vccd1 _19955_/Q sky130_fd_sc_hd__dfxtp_1
X_15078_ _15078_/A vssd1 vssd1 vccd1 vccd1 _19072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14029_ _18646_/Q _13660_/X _14035_/S vssd1 vssd1 vccd1 vccd1 _14030_/A sky130_fd_sc_hd__mux2_1
X_18906_ _19366_/CLK _18906_/D vssd1 vssd1 vccd1 vccd1 _18906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19886_ _20044_/CLK _19886_/D vssd1 vssd1 vccd1 vccd1 _19886_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18837_ _18973_/CLK _18837_/D vssd1 vssd1 vccd1 vccd1 _18837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09570_ _18794_/Q _19065_/Q _19289_/Q _19033_/Q _09568_/X _09762_/A vssd1 vssd1 vccd1
+ vccd1 _09570_/X sky130_fd_sc_hd__mux4_1
X_18768_ _19489_/CLK _18768_/D vssd1 vssd1 vccd1 vccd1 _18768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17719_ _17719_/A vssd1 vssd1 vccd1 vccd1 _17719_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18699_ _19734_/CLK _18699_/D vssd1 vssd1 vccd1 vccd1 _18699_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11415__A _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14726__A _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13630__A _14589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10465__S _10465_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clock_A clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09555__A _11204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10480__S0 _10559_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09906_ _10254_/A _09900_/X _09903_/X _09905_/X vssd1 vssd1 vccd1 vccd1 _09906_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17772__A _17772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09274__B _17331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20026_ _20027_/CLK _20026_/D vssd1 vssd1 vccd1 vccd1 _20026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09837_ _09901_/A vssd1 vssd1 vccd1 vccd1 _09904_/S sky130_fd_sc_hd__buf_4
XANTENNA__10232__S0 _09872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15292__A _15292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09768_ _18599_/Q _18860_/Q _18759_/Q _19094_/Q _09761_/S _09569_/A vssd1 vssd1 vccd1
+ vccd1 _09769_/B sky130_fd_sc_hd__mux4_1
XFILLER_100_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _09699_/A _09699_/B vssd1 vssd1 vccd1 vccd1 _09699_/Y sky130_fd_sc_hd__nor2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _11730_/A _11730_/B _11730_/C vssd1 vssd1 vccd1 vccd1 _11730_/X sky130_fd_sc_hd__or3_1
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10860__A1 _10052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11661_/A vssd1 vssd1 vccd1 vccd1 _11661_/X sky130_fd_sc_hd__clkbuf_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _19796_/Q vssd1 vssd1 vccd1 vccd1 _17104_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13540__A _15295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10612_ _10604_/X _10607_/X _10610_/X _11362_/A _09475_/A vssd1 vssd1 vccd1 vccd1
+ _10623_/B sky130_fd_sc_hd__o221a_1
X_14380_ _18797_/Q _14379_/X _14386_/S vssd1 vssd1 vccd1 vccd1 _14381_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11404__A3 _11402_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11592_ _11557_/X _11558_/Y _11559_/X _11560_/Y _11591_/X vssd1 vssd1 vccd1 vccd1
+ _11592_/X sky130_fd_sc_hd__a221o_1
XFILLER_128_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ _15257_/A vssd1 vssd1 vccd1 vccd1 _13331_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10543_ _19372_/Q _18986_/Q _19436_/Q _18555_/Q _10337_/A _09855_/A vssd1 vssd1 vccd1
+ vccd1 _10544_/B sky130_fd_sc_hd__mux4_1
XFILLER_109_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16050_ _13471_/X _19446_/Q _16056_/S vssd1 vssd1 vccd1 vccd1 _16051_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13262_ input6/X _13172_/A _13175_/A vssd1 vssd1 vccd1 vccd1 _13276_/A sky130_fd_sc_hd__a21o_1
X_10474_ _10314_/X _10464_/X _10468_/X _10473_/X _10519_/A vssd1 vssd1 vccd1 vccd1
+ _10474_/X sky130_fd_sc_hd__a311o_1
XFILLER_108_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_160_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19805_/CLK sky130_fd_sc_hd__clkbuf_16
X_15001_ _15001_/A vssd1 vssd1 vccd1 vccd1 _19038_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13686__S _13694_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09766__C1 _09479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12213_ _19529_/Q _12206_/X _12208_/X _12211_/X _12212_/X vssd1 vssd1 vccd1 vccd1
+ _12213_/X sky130_fd_sc_hd__o221a_1
XFILLER_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13193_ _13337_/A _13189_/X _13191_/Y _13192_/X _13351_/A vssd1 vssd1 vccd1 vccd1
+ _13194_/B sky130_fd_sc_hd__a221o_1
XFILLER_155_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10471__S0 _10470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12144_ _12144_/A _12172_/A vssd1 vssd1 vccd1 vccd1 _12147_/A sky130_fd_sc_hd__nor2_1
XFILLER_123_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_2_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13314__B1 _13299_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19740_ _19852_/CLK _19740_/D vssd1 vssd1 vccd1 vccd1 _19740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16952_ _16957_/B _16946_/B _19745_/Q vssd1 vssd1 vccd1 vccd1 _16956_/B sky130_fd_sc_hd__a21oi_1
X_12075_ _19968_/Q vssd1 vssd1 vccd1 vccd1 _12075_/Y sky130_fd_sc_hd__clkinv_2
Xclkbuf_leaf_175_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19865_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_6_clock_A _19998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_159_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10223__S0 _09872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15903_ _15903_/A vssd1 vssd1 vccd1 vccd1 _15912_/S sky130_fd_sc_hd__clkbuf_4
X_11026_ _18673_/Q _19168_/Q _11026_/S vssd1 vssd1 vccd1 vccd1 _11027_/A sky130_fd_sc_hd__mux2_1
X_19671_ _19671_/CLK _19671_/D vssd1 vssd1 vccd1 vccd1 _19671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16883_ _16922_/C _19724_/Q _19723_/Q _16883_/D vssd1 vssd1 vccd1 vccd1 _16891_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15406__S _15406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18622_ _19503_/CLK _18622_/D vssd1 vssd1 vccd1 vccd1 _18622_/Q sky130_fd_sc_hd__dfxtp_1
X_15834_ _19922_/Q _15833_/X _15840_/S vssd1 vssd1 vccd1 vccd1 _15834_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18553_ _19575_/CLK _18553_/D vssd1 vssd1 vccd1 vccd1 _18553_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09916__S0 _10244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ _18462_/Q _12973_/X _09947_/A _12976_/X vssd1 vssd1 vccd1 vccd1 _18462_/D
+ sky130_fd_sc_hd__a22o_1
X_15765_ _19911_/Q _15764_/Y _15800_/S vssd1 vssd1 vccd1 vccd1 _15765_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09297__A1 _11704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _12614_/B _12673_/B _17504_/S vssd1 vssd1 vccd1 vccd1 _17802_/C sky130_fd_sc_hd__mux2_2
X_14716_ _18911_/Q _14420_/X _14724_/S vssd1 vssd1 vccd1 vccd1 _14717_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11928_ _11928_/A vssd1 vssd1 vccd1 vccd1 _12194_/A sky130_fd_sc_hd__clkbuf_2
X_18484_ _19561_/CLK _18484_/D vssd1 vssd1 vccd1 vccd1 _18484_/Q sky130_fd_sc_hd__dfxtp_1
X_15696_ _15814_/A _17166_/A vssd1 vssd1 vccd1 vccd1 _16235_/A sky130_fd_sc_hd__nor2_1
XFILLER_75_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14647_ _14647_/A vssd1 vssd1 vccd1 vccd1 _14647_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10851__A1 _10665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17435_ _17610_/B _12574_/A _17465_/S vssd1 vssd1 vccd1 vccd1 _17435_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11859_ _11860_/A _17418_/A vssd1 vssd1 vccd1 vccd1 _11861_/A sky130_fd_sc_hd__and2_1
XFILLER_159_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_113_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19576_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16319__A0 _19535_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14578_ _14574_/X _18864_/Q _14590_/S vssd1 vssd1 vccd1 vccd1 _14579_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15790__A1 _18459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _09209_/Y _18301_/A _17358_/X _13173_/B vssd1 vssd1 vccd1 vccd1 _17367_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10064__C1 _10063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19105_ _19201_/CLK _19105_/D vssd1 vssd1 vccd1 vccd1 _19105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13529_ _19804_/Q _13117_/A _12805_/Y _19640_/Q _13528_/X vssd1 vssd1 vccd1 vccd1
+ _13529_/X sky130_fd_sc_hd__a221o_2
X_16317_ _16317_/A _16317_/B vssd1 vssd1 vccd1 vccd1 _16317_/X sky130_fd_sc_hd__xor2_1
XFILLER_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17297_ _17297_/A vssd1 vssd1 vccd1 vccd1 _19871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19036_ _19484_/CLK _19036_/D vssd1 vssd1 vccd1 vccd1 _19036_/Q sky130_fd_sc_hd__dfxtp_1
X_16248_ _16248_/A _19934_/Q _16248_/C vssd1 vssd1 vccd1 vccd1 _16255_/B sky130_fd_sc_hd__or3_1
XFILLER_174_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_128_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19490_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13553__A0 _19924_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11159__A2 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput103 _09202_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[0] sky130_fd_sc_hd__buf_2
XFILLER_115_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput114 _12650_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[14] sky130_fd_sc_hd__buf_2
XFILLER_161_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16179_ _16179_/A vssd1 vssd1 vccd1 vccd1 _19503_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09221__A1 _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14281__A _14281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput125 _12662_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[24] sky130_fd_sc_hd__buf_2
XFILLER_154_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput136 _12637_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[5] sky130_fd_sc_hd__buf_2
XFILLER_126_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput147 _16471_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[14] sky130_fd_sc_hd__buf_2
Xoutput158 _12448_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[24] sky130_fd_sc_hd__buf_2
XFILLER_115_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput169 _11924_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19938_ _19938_/CLK _19938_/D vssd1 vssd1 vccd1 vccd1 _19938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19869_ _19873_/CLK _19869_/D vssd1 vssd1 vccd1 vccd1 _19869_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10765__S1 _10037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ _09622_/A vssd1 vssd1 vccd1 vccd1 _09623_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13625__A _15209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14220__S _14222_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _11116_/A vssd1 vssd1 vccd1 vccd1 _11315_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09484_ _11489_/A vssd1 vssd1 vccd1 vccd1 _11473_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_102_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10842__A1 _10730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15051__S _15055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15986__S _15988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__S _10195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10453__S0 _10325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ _10184_/A _10189_/X _09712_/A vssd1 vssd1 vccd1 vccd1 _10190_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_92_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _18845_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16494__C1 _12749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_160_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11858__A0 _19961_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10756__S1 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12900_ _19665_/Q _12887_/X _12889_/X _19797_/Q _12899_/X vssd1 vssd1 vccd1 vccd1
+ _12901_/B sky130_fd_sc_hd__a221o_4
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09920__C1 _09605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20009_ _20020_/CLK _20009_/D vssd1 vssd1 vccd1 vccd1 _20009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13880_ _13926_/S vssd1 vssd1 vccd1 vccd1 _13889_/S sky130_fd_sc_hd__buf_4
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12831_ _18198_/A vssd1 vssd1 vccd1 vccd1 _16315_/A sky130_fd_sc_hd__buf_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _19272_/Q _15244_/X _15550_/S vssd1 vssd1 vccd1 vccd1 _15551_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11086__A1 _10914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_30_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19561_/CLK sky130_fd_sc_hd__clkbuf_16
X_12762_ _19808_/Q _12684_/C _12696_/X _19834_/Q _12761_/X vssd1 vssd1 vccd1 vccd1
+ _12762_/X sky130_fd_sc_hd__a221o_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _18293_/A _14501_/B vssd1 vssd1 vccd1 vccd1 _15589_/B sky130_fd_sc_hd__nand2_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10833__A1 _09989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _19958_/Q _11302_/A _11809_/A vssd1 vssd1 vccd1 vccd1 _11764_/C sky130_fd_sc_hd__mux2_4
X_15481_ _19241_/Q _15247_/X _15489_/S vssd1 vssd1 vccd1 vccd1 _15482_/A sky130_fd_sc_hd__mux2_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _13136_/D _12693_/C vssd1 vssd1 vccd1 vccd1 _13205_/A sky130_fd_sc_hd__and3_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _14432_/A vssd1 vssd1 vccd1 vccd1 _18813_/D sky130_fd_sc_hd__clkbuf_1
X_17220_ _17220_/A vssd1 vssd1 vccd1 vccd1 _17220_/Y sky130_fd_sc_hd__inv_2
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11704_/B vssd1 vssd1 vccd1 vccd1 _11901_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10046__C1 _09738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17151_ _13572_/X _17164_/B _17150_/X _18412_/A vssd1 vssd1 vccd1 vccd1 _19817_/D
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_45_clock clkbuf_opt_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19476_/CLK sky130_fd_sc_hd__clkbuf_16
X_14363_ _18792_/Q _13735_/X _14363_/S vssd1 vssd1 vccd1 vccd1 _14364_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput16 io_dbus_rdata[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_85_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11575_ _11575_/A _11578_/A _11575_/C vssd1 vssd1 vccd1 vccd1 _11575_/Y sky130_fd_sc_hd__nand3_1
XFILLER_11_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput27 io_dbus_rdata[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_2
X_16102_ _13321_/X _19469_/Q _16106_/S vssd1 vssd1 vccd1 vccd1 _16103_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput38 io_ibus_inst[13] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13314_ _16301_/A _13312_/B _13299_/C vssd1 vssd1 vccd1 vccd1 _13315_/B sky130_fd_sc_hd__o21ai_1
X_10526_ _10571_/A _10526_/B vssd1 vssd1 vccd1 vccd1 _10526_/X sky130_fd_sc_hd__or2_1
XFILLER_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput49 io_ibus_inst[23] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
X_17082_ _17082_/A vssd1 vssd1 vccd1 vccd1 _17087_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10692__S0 _10690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14294_ _13850_/X _18762_/Q _14294_/S vssd1 vssd1 vccd1 vccd1 _14295_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16033_ _16033_/A vssd1 vssd1 vccd1 vccd1 _19438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15197__A _15197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ _13245_/A vssd1 vssd1 vccd1 vccd1 _13245_/X sky130_fd_sc_hd__clkbuf_2
X_10457_ _09749_/A _10446_/X _10455_/X _09756_/A _10456_/Y vssd1 vssd1 vccd1 vccd1
+ _12655_/B sky130_fd_sc_hd__o32a_4
XFILLER_171_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13176_ input31/X _13172_/X _13175_/X vssd1 vssd1 vccd1 vccd1 _13176_/X sky130_fd_sc_hd__a21o_1
X_10388_ _19117_/Q _18883_/Q _19565_/Q _19213_/Q _09651_/A _10440_/A vssd1 vssd1 vccd1
+ vccd1 _10389_/B sky130_fd_sc_hd__mux4_1
XFILLER_123_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12127_ _12127_/A vssd1 vssd1 vccd1 vccd1 _12127_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__15827__A2 _13502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17984_ _17989_/B _17985_/B vssd1 vssd1 vccd1 vccd1 _17988_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10134__A _19920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18301__A _18301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19723_ _19737_/CLK _19723_/D vssd1 vssd1 vccd1 vccd1 _19723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16935_ _16936_/B _16935_/B vssd1 vssd1 vccd1 vccd1 _19740_/D sky130_fd_sc_hd__nor2_1
X_12058_ _19588_/Q vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11009_ _18577_/Q _18838_/Q _18737_/Q _19072_/Q _10937_/S _09954_/A vssd1 vssd1 vccd1
+ vccd1 _11010_/B sky130_fd_sc_hd__mux4_1
XANTENNA__14040__S _14046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19654_ _19789_/CLK _19654_/D vssd1 vssd1 vccd1 vccd1 _19654_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_6_0_clock_A clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16866_ _16920_/B _16865_/A _16870_/D _18365_/A vssd1 vssd1 vccd1 vccd1 _16866_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_93_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18605_ _19484_/CLK _18605_/D vssd1 vssd1 vccd1 vccd1 _18605_/Q sky130_fd_sc_hd__dfxtp_1
X_15817_ _15817_/A vssd1 vssd1 vccd1 vccd1 _19350_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13164__B _19901_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14975__S _14983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19585_ _19966_/CLK _19585_/D vssd1 vssd1 vccd1 vccd1 _19585_/Q sky130_fd_sc_hd__dfxtp_1
X_16797_ _19703_/Q _16793_/B _16796_/Y vssd1 vssd1 vccd1 vccd1 _19703_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18536_ _19063_/CLK _18536_/D vssd1 vssd1 vccd1 vccd1 _18536_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _15748_/A vssd1 vssd1 vccd1 vccd1 _19338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ _19938_/CLK _18467_/D vssd1 vssd1 vccd1 vccd1 _18467_/Q sky130_fd_sc_hd__dfxtp_1
X_15679_ _18441_/Q _15679_/B vssd1 vssd1 vccd1 vccd1 _15679_/X sky130_fd_sc_hd__or2_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17418_ _17418_/A vssd1 vssd1 vccd1 vccd1 _17729_/B sky130_fd_sc_hd__buf_2
XFILLER_21_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18398_ input39/X vssd1 vssd1 vccd1 vccd1 _18398_/Y sky130_fd_sc_hd__inv_12
XANTENNA__16960__B1 _16833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17349_ _17349_/A vssd1 vssd1 vccd1 vccd1 _19884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10683__S0 _10608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19019_ _19501_/CLK _19019_/D vssd1 vssd1 vccd1 vccd1 _19019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10435__S0 _10325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10760__B1 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18211__A _18268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10512__B1 _10296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ _09605_/A vssd1 vssd1 vccd1 vccd1 _09605_/X sky130_fd_sc_hd__buf_2
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14885__S _14889_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09536_ _10382_/A vssd1 vssd1 vccd1 vccd1 _10417_/S sky130_fd_sc_hd__buf_2
XFILLER_58_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09467_ _11680_/C _09467_/B vssd1 vssd1 vccd1 vccd1 _17323_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_107_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ _09398_/A _09398_/B _11833_/A vssd1 vssd1 vccd1 vccd1 _12701_/A sky130_fd_sc_hd__or3b_1
XFILLER_8_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10219__A _10219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16832__C _16832_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11360_ _11575_/A _11578_/A _11575_/C _11574_/A _11359_/X vssd1 vssd1 vccd1 vccd1
+ _11570_/C sky130_fd_sc_hd__a311o_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10311_ _10380_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10311_/X sky130_fd_sc_hd__or2_1
XFILLER_3_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14125__S _14131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11291_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13030_ _09345_/X _13029_/X _13553_/S vssd1 vssd1 vccd1 vccd1 _13030_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10242_ _19119_/Q _18885_/Q _19567_/Q _19215_/Q _09902_/S _09822_/A vssd1 vssd1 vccd1
+ vccd1 _10243_/B sky130_fd_sc_hd__mux4_1
XFILLER_105_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13964__S _13972_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10173_ _18690_/Q _19185_/Q _10173_/S vssd1 vssd1 vccd1 vccd1 _10174_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input38_A io_ibus_inst[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14981_ _19030_/Q _14462_/X _14983_/S vssd1 vssd1 vccd1 vccd1 _14982_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10729__S1 _10609_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_opt_5_0_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16720_ _16729_/D vssd1 vssd1 vccd1 vccd1 _16727_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13932_ _13932_/A vssd1 vssd1 vccd1 vccd1 _18603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13863_ _13758_/X _18573_/Q _13867_/S vssd1 vssd1 vccd1 vccd1 _13864_/A sky130_fd_sc_hd__mux2_1
X_16651_ _16653_/B _16653_/C _16624_/X vssd1 vssd1 vccd1 vccd1 _16651_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14795__S _14797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17982__A2 _17861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15480__A _15502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ _12853_/A _12814_/B vssd1 vssd1 vccd1 vccd1 _12814_/Y sky130_fd_sc_hd__nor2_4
X_15602_ _15659_/S vssd1 vssd1 vccd1 vccd1 _15611_/S sky130_fd_sc_hd__buf_2
XFILLER_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19370_ _19560_/CLK _19370_/D vssd1 vssd1 vccd1 vccd1 _19370_/Q sky130_fd_sc_hd__dfxtp_1
X_13794_ _13793_/X _18552_/Q _13797_/S vssd1 vssd1 vccd1 vccd1 _13795_/A sky130_fd_sc_hd__mux2_1
X_16582_ _19634_/Q _19633_/Q _16582_/C vssd1 vssd1 vccd1 vccd1 _16584_/B sky130_fd_sc_hd__and3_1
XFILLER_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18321_ _18321_/A _18333_/B vssd1 vssd1 vccd1 vccd1 _18321_/X sky130_fd_sc_hd__or2_1
XANTENNA__11154__S1 _11330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12745_ _19809_/Q _18281_/B _17245_/S vssd1 vssd1 vccd1 vccd1 _12745_/X sky130_fd_sc_hd__or3_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15533_ _19264_/Q _15219_/X _15539_/S vssd1 vssd1 vccd1 vccd1 _15534_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12609__A _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ _15464_/A vssd1 vssd1 vccd1 vccd1 _19233_/D sky130_fd_sc_hd__clkbuf_1
X_18252_ _18252_/A vssd1 vssd1 vccd1 vccd1 _19980_/D sky130_fd_sc_hd__clkbuf_1
X_12676_ _12914_/B vssd1 vssd1 vccd1 vccd1 _12893_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _18808_/Q _14414_/X _14418_/S vssd1 vssd1 vccd1 vccd1 _14416_/A sky130_fd_sc_hd__mux2_1
X_17203_ _19834_/Q _17210_/B vssd1 vssd1 vccd1 vccd1 _17203_/X sky130_fd_sc_hd__or2_1
XANTENNA__17396__A_N _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11627_ _11645_/B _11627_/B _11627_/C _11682_/A vssd1 vssd1 vccd1 vccd1 _12596_/B
+ sky130_fd_sc_hd__and4_2
X_15395_ _14605_/X _19203_/Q _15395_/S vssd1 vssd1 vccd1 vccd1 _15396_/A sky130_fd_sc_hd__mux2_1
X_18183_ _18183_/A vssd1 vssd1 vccd1 vccd1 _18192_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_156_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17498__A1 _17749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14346_ _18784_/Q _13702_/X _14352_/S vssd1 vssd1 vccd1 vccd1 _14347_/A sky130_fd_sc_hd__mux2_1
X_17134_ input67/X _17138_/B vssd1 vssd1 vccd1 vccd1 _17134_/X sky130_fd_sc_hd__or2_1
XANTENNA__11231__A1 _10920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11558_ _11558_/A _11558_/B vssd1 vssd1 vccd1 vccd1 _11558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10509_ _18811_/Q _19146_/Q _10509_/S vssd1 vssd1 vccd1 vccd1 _10510_/B sky130_fd_sc_hd__mux2_1
X_17065_ _17065_/A vssd1 vssd1 vccd1 vccd1 _17070_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14277_ _13825_/X _18754_/Q _14279_/S vssd1 vssd1 vccd1 vccd1 _14278_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14035__S _14035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16170__A1 _14624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11489_ _11489_/A _11489_/B vssd1 vssd1 vccd1 vccd1 _11489_/X sky130_fd_sc_hd__or2_1
XFILLER_143_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16016_ _16016_/A vssd1 vssd1 vccd1 vccd1 _19430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13228_ input3/X _13172_/X _13175_/X vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13874__S _13878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _19618_/Q vssd1 vssd1 vccd1 vccd1 _16538_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11090__S0 _11147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09653__A _09653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16473__A2 _16449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17670__B2 _11767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17967_ _17560_/A _17957_/Y _17965_/X _17966_/Y vssd1 vssd1 vccd1 vccd1 _17967_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_111_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19706_ _19877_/CLK _19706_/D vssd1 vssd1 vccd1 vccd1 _19706_/Q sky130_fd_sc_hd__dfxtp_1
X_16918_ _19737_/Q _19736_/Q _16925_/B _16918_/D vssd1 vssd1 vccd1 vccd1 _16955_/A
+ sky130_fd_sc_hd__and4_4
X_17898_ _17914_/A vssd1 vssd1 vccd1 vccd1 _18033_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17422__A1 _12480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19637_ _19637_/CLK _19637_/D vssd1 vssd1 vccd1 vccd1 _19637_/Q sky130_fd_sc_hd__dfxtp_1
X_16849_ _16946_/A _16857_/D vssd1 vssd1 vccd1 vccd1 _16849_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19568_ _19569_/CLK _19568_/D vssd1 vssd1 vccd1 vccd1 _19568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11145__S1 _09658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09321_ _12611_/A _09751_/B _09751_/C vssd1 vssd1 vccd1 vccd1 _09321_/X sky130_fd_sc_hd__or3_1
X_18519_ _19498_/CLK _18519_/D vssd1 vssd1 vccd1 vccd1 _18519_/Q sky130_fd_sc_hd__dfxtp_1
X_19499_ _19500_/CLK _19499_/D vssd1 vssd1 vccd1 vccd1 _19499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09252_ _11648_/A _11648_/C vssd1 vssd1 vccd1 vccd1 _12594_/C sky130_fd_sc_hd__nor2_2
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09183_ _11785_/A _11787_/A _11786_/A vssd1 vssd1 vccd1 vccd1 _11646_/C sky130_fd_sc_hd__nor3b_1
XANTENNA__10039__A _10039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09828__A _10205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12970__A1 _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10981__B1 _10980_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10408__S0 _10268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11525__A2 _11534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17110__B1 _17101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_33_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15672__B1 _13592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17413__A1 _12432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__B1 _13353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10860_ _10052_/X _10859_/X _10056_/X vssd1 vssd1 vccd1 vccd1 _10860_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11136__S1 _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ _09841_/A vssd1 vssd1 vccd1 vccd1 _09520_/A sky130_fd_sc_hd__buf_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12789__B2 _18455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ _19462_/Q _19300_/Q _18709_/Q _18479_/Q _10048_/A _10037_/A vssd1 vssd1 vccd1
+ vccd1 _10792_/B sky130_fd_sc_hd__mux4_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12429__A _12429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12531_/A _18090_/B vssd1 vssd1 vccd1 vccd1 _12532_/A sky130_fd_sc_hd__nand2_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13959__S _13961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12461_ _12482_/A _12436_/B _12460_/Y vssd1 vssd1 vccd1 vccd1 _12462_/B sky130_fd_sc_hd__o21a_1
X_14200_ _14200_/A vssd1 vssd1 vccd1 vccd1 _18719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11412_ _10674_/Y _11569_/B _11567_/A _10673_/A vssd1 vssd1 vccd1 vccd1 _11565_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15180_ _15180_/A vssd1 vssd1 vccd1 vccd1 _19121_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09738__A _09738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ _19600_/Q _12393_/B vssd1 vssd1 vccd1 vccd1 _12394_/A sky130_fd_sc_hd__nor2_1
XFILLER_137_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14131_ _18691_/Q _13714_/X _14131_/S vssd1 vssd1 vccd1 vccd1 _14132_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12961__A1 _18451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ _18635_/Q _19226_/Q _19388_/Q _18603_/Q _11030_/A _09658_/A vssd1 vssd1 vccd1
+ vccd1 _11343_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09457__B _17346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16152__A1 _14599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14062_ _18661_/Q _13723_/X _14068_/S vssd1 vssd1 vccd1 vccd1 _14063_/A sky130_fd_sc_hd__mux2_1
X_11274_ _11274_/A _11274_/B vssd1 vssd1 vccd1 vccd1 _11274_/X sky130_fd_sc_hd__or2_1
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13694__S _13694_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13013_ _19998_/Q vssd1 vssd1 vccd1 vccd1 _14844_/C sky130_fd_sc_hd__clkbuf_4
X_10225_ _18785_/Q _19056_/Q _19280_/Q _19024_/Q _09653_/A _09927_/A vssd1 vssd1 vccd1
+ vccd1 _10225_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11072__S0 _11000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18870_ _19200_/CLK _18870_/D vssd1 vssd1 vccd1 vccd1 _18870_/Q sky130_fd_sc_hd__dfxtp_1
X_17821_ _18000_/A _17817_/X _17820_/X _17533_/A vssd1 vssd1 vccd1 vccd1 _17821_/X
+ sky130_fd_sc_hd__o211a_1
X_10156_ _10156_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _10156_/X sky130_fd_sc_hd__or2_1
XFILLER_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12477__B1 _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17752_ _17524_/X _17745_/Y _17751_/X _17667_/A vssd1 vssd1 vccd1 vccd1 _17752_/X
+ sky130_fd_sc_hd__a211o_1
X_10087_ _18598_/Q _18859_/Q _18758_/Q _19093_/Q _11483_/S _10618_/A vssd1 vssd1 vccd1
+ vccd1 _10088_/B sky130_fd_sc_hd__mux4_1
X_14964_ _19022_/Q _14436_/X _14972_/S vssd1 vssd1 vccd1 vccd1 _14965_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16703_ _19797_/Q _19796_/Q _19798_/Q _17098_/A vssd1 vssd1 vccd1 vccd1 _17107_/A
+ sky130_fd_sc_hd__and4_1
X_13915_ _13915_/A vssd1 vssd1 vccd1 vccd1 _18596_/D sky130_fd_sc_hd__clkbuf_1
X_17683_ _17562_/X _17564_/X _17802_/D vssd1 vssd1 vccd1 vccd1 _17683_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14895_ _14895_/A vssd1 vssd1 vccd1 vccd1 _18991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19422_ _19666_/CLK _19422_/D vssd1 vssd1 vccd1 vccd1 _19422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16634_ _16636_/B _16636_/C _16633_/Y vssd1 vssd1 vccd1 vccd1 _19652_/D sky130_fd_sc_hd__o21a_1
XFILLER_63_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13846_ _13846_/A vssd1 vssd1 vccd1 vccd1 _18568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19353_ _19879_/CLK _19353_/D vssd1 vssd1 vccd1 vccd1 _19353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16565_ _16573_/A _16565_/B _16566_/B vssd1 vssd1 vccd1 vccd1 _19628_/D sky130_fd_sc_hd__nor3_1
X_13777_ _14602_/A vssd1 vssd1 vccd1 vccd1 _13777_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10989_ _11216_/A _10987_/X _10988_/X vssd1 vssd1 vccd1 vccd1 _10989_/Y sky130_fd_sc_hd__o21ai_1
X_18304_ _20001_/Q _18285_/X _18302_/Y _18303_/X vssd1 vssd1 vccd1 vccd1 _20001_/D
+ sky130_fd_sc_hd__o211a_1
X_15516_ _15516_/A vssd1 vssd1 vccd1 vccd1 _19257_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19284_ _19510_/CLK _19284_/D vssd1 vssd1 vccd1 vccd1 _19284_/Q sky130_fd_sc_hd__dfxtp_1
X_12728_ _12888_/A vssd1 vssd1 vccd1 vccd1 _13117_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10886__S0 _09983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16496_ _19647_/Q _19646_/Q _19648_/Q _16612_/A vssd1 vssd1 vccd1 vccd1 _16620_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_31_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18235_ _18235_/A vssd1 vssd1 vccd1 vccd1 _19972_/D sky130_fd_sc_hd__clkbuf_1
X_12659_ _12663_/A _12659_/B vssd1 vssd1 vccd1 vccd1 _12659_/Y sky130_fd_sc_hd__nor2_2
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15447_ _15515_/S vssd1 vssd1 vccd1 vccd1 _15456_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_129_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18166_ _16301_/A _19974_/Q _18170_/S vssd1 vssd1 vccd1 vccd1 _18167_/A sky130_fd_sc_hd__mux2_1
X_15378_ _14580_/X _19195_/Q _15384_/S vssd1 vssd1 vccd1 vccd1 _15379_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11755__A2 _12937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17117_ _19801_/Q _17114_/B _17116_/Y vssd1 vssd1 vccd1 vccd1 _19801_/D sky130_fd_sc_hd__o21a_1
XFILLER_172_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10293__S _10417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14329_ _14329_/A vssd1 vssd1 vccd1 vccd1 _18776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18097_ _18098_/B _18097_/B vssd1 vssd1 vccd1 vccd1 _18101_/B sky130_fd_sc_hd__nand2_1
XFILLER_143_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17048_ _17066_/A _17053_/C vssd1 vssd1 vccd1 vccd1 _17048_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09870_ _10403_/A vssd1 vssd1 vccd1 vccd1 _10279_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ _19481_/CLK _18999_/D vssd1 vssd1 vccd1 vccd1 _18999_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11676__D1 _12602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17946__A2 _17949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13633__A _15215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09304_ _09304_/A _11684_/A vssd1 vssd1 vccd1 vccd1 _17391_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10877__S0 _09983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09731__S1 _09730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12640__B1 _12670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09235_ _09238_/A vssd1 vssd1 vccd1 vccd1 _11730_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12943__A1 _12942_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15295__A _15295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__S0 _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12712__A _12837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10010_ _10054_/A vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13527__B _13527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09999_ _09999_/A vssd1 vssd1 vccd1 vccd1 _10655_/A sky130_fd_sc_hd__buf_2
XFILLER_135_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13120__B2 _19520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15742__B _18451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11961_ _11961_/A vssd1 vssd1 vccd1 vccd1 _12069_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13700_ _13700_/A vssd1 vssd1 vccd1 vccd1 _18527_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17015__A _17073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10912_ _18579_/Q _18840_/Q _18739_/Q _19074_/Q _11493_/S _09660_/A vssd1 vssd1 vccd1
+ vccd1 _10912_/X sky130_fd_sc_hd__mux4_1
X_14680_ _15445_/B _16134_/B vssd1 vssd1 vccd1 vccd1 _14737_/A sky130_fd_sc_hd__nor2_8
X_11892_ _11892_/A _11892_/B vssd1 vssd1 vccd1 vccd1 _11893_/A sky130_fd_sc_hd__and2_2
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11109__S1 _11065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13631_ _18511_/Q _13630_/X _13631_/S vssd1 vssd1 vccd1 vccd1 _13632_/A sky130_fd_sc_hd__mux2_1
X_10843_ _10836_/X _10838_/X _10840_/X _10842_/X _09602_/A vssd1 vssd1 vccd1 vccd1
+ _10843_/X sky130_fd_sc_hd__a221o_1
XFILLER_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13562_ _13562_/A _13562_/B vssd1 vssd1 vccd1 vccd1 _13562_/Y sky130_fd_sc_hd__nand2_1
X_16350_ _12215_/X _15822_/X _16223_/S vssd1 vssd1 vccd1 vccd1 _16350_/X sky130_fd_sc_hd__a21bo_1
XFILLER_158_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10774_ _12076_/A _12647_/A vssd1 vssd1 vccd1 vccd1 _11570_/B sky130_fd_sc_hd__or2_1
XFILLER_157_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15301_ _15301_/A _15373_/C _15445_/B vssd1 vssd1 vccd1 vccd1 _15358_/A sky130_fd_sc_hd__nor3_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12513_ _12509_/Y _12512_/Y _12562_/S vssd1 vssd1 vccd1 vccd1 _12513_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10642__C1 _10757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16281_ _16281_/A vssd1 vssd1 vccd1 vccd1 _19528_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16065__S _16073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13493_ _13512_/B _13492_/Y _11607_/X vssd1 vssd1 vccd1 vccd1 _13493_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18020_ _18023_/A _18023_/B vssd1 vssd1 vccd1 vccd1 _18020_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15232_ _15299_/S vssd1 vssd1 vccd1 vccd1 _15245_/S sky130_fd_sc_hd__buf_2
X_12444_ _12444_/A vssd1 vssd1 vccd1 vccd1 _12444_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15163_ _19113_/Q vssd1 vssd1 vccd1 vccd1 _15164_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_60_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12375_ _19599_/Q _12363_/X _12371_/Y _12374_/Y vssd1 vssd1 vccd1 vccd1 _12375_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_154_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14114_ _18683_/Q _13681_/X _14120_/S vssd1 vssd1 vccd1 vccd1 _14115_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11326_ _11342_/A _11326_/B vssd1 vssd1 vccd1 vccd1 _11326_/Y sky130_fd_sc_hd__nor2_1
X_15094_ _14621_/X _19080_/Q _15094_/S vssd1 vssd1 vccd1 vccd1 _15095_/A sky130_fd_sc_hd__mux2_1
X_19971_ _19971_/CLK _19971_/D vssd1 vssd1 vccd1 vccd1 _19971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15409__S _15417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ _14045_/A vssd1 vssd1 vccd1 vccd1 _18653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18922_ _19478_/CLK _18922_/D vssd1 vssd1 vccd1 vccd1 _18922_/Q sky130_fd_sc_hd__dfxtp_1
X_11257_ _11317_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11257_/X sky130_fd_sc_hd__or2_1
XANTENNA__11045__S0 _10914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14313__S _14319_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ _19506_/Q _18918_/Q _18955_/Q _18529_/Q _10160_/S _09809_/A vssd1 vssd1 vccd1
+ vccd1 _10209_/B sky130_fd_sc_hd__mux4_1
XFILLER_122_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18853_ _19311_/CLK _18853_/D vssd1 vssd1 vccd1 vccd1 _18853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11188_ _09745_/A _11176_/X _11186_/X _09752_/A _11187_/Y vssd1 vssd1 vccd1 vccd1
+ _12633_/B sky130_fd_sc_hd__o32a_4
X_17804_ _17802_/X _17694_/X _17803_/X _17845_/A vssd1 vssd1 vccd1 vccd1 _17804_/X
+ sky130_fd_sc_hd__o22a_1
X_10139_ _10139_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _10139_/X sky130_fd_sc_hd__or2_1
XFILLER_95_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18784_ _19409_/CLK _18784_/D vssd1 vssd1 vccd1 vccd1 _18784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15996_ _15996_/A vssd1 vssd1 vccd1 vccd1 _19421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17735_ _19897_/Q _09419_/X _17733_/X _17734_/Y vssd1 vssd1 vccd1 vccd1 _19897_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14947_ _14947_/A vssd1 vssd1 vccd1 vccd1 _19014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13453__A _15279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17666_ _17656_/X _17664_/Y _17666_/S vssd1 vssd1 vccd1 vccd1 _17667_/B sky130_fd_sc_hd__mux2_1
X_14878_ _14621_/X _18984_/Q _14878_/S vssd1 vssd1 vccd1 vccd1 _14879_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19405_ _19405_/CLK _19405_/D vssd1 vssd1 vccd1 vccd1 _19405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16617_ _19647_/Q _16617_/B _16617_/C vssd1 vssd1 vccd1 vccd1 _16619_/B sky130_fd_sc_hd__and3_1
X_13829_ _13828_/X _18563_/Q _13829_/S vssd1 vssd1 vccd1 vccd1 _13830_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14983__S _14983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17597_ _18072_/A vssd1 vssd1 vccd1 vccd1 _17953_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19336_ _19881_/CLK _19336_/D vssd1 vssd1 vccd1 vccd1 _19336_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10859__S0 _10753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16548_ _16573_/A _16548_/B _16548_/C vssd1 vssd1 vccd1 vccd1 _19622_/D sky130_fd_sc_hd__nor3_1
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19267_ _19493_/CLK _19267_/D vssd1 vssd1 vccd1 vccd1 _19267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16479_ _12339_/C _16477_/X _12313_/X _12317_/Y _16468_/X vssd1 vssd1 vccd1 vccd1
+ _19597_/D sky130_fd_sc_hd__o221a_1
X_18218_ _19965_/Q _12027_/A _18220_/S vssd1 vssd1 vccd1 vccd1 _18219_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19198_ _19455_/CLK _19198_/D vssd1 vssd1 vccd1 vccd1 _19198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18149_ _18149_/A vssd1 vssd1 vccd1 vccd1 _19934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16930__C _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17864__A1 _17866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09922_ _19122_/Q _18888_/Q _19570_/Q _19218_/Q _10173_/S _10271_/A vssd1 vssd1 vccd1
+ vccd1 _09923_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10751__S _10751_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13350__A1 _15768_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09853_ _09926_/S vssd1 vssd1 vccd1 vccd1 _10175_/S sky130_fd_sc_hd__buf_4
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20042_ _20044_/CLK _20042_/D vssd1 vssd1 vccd1 vccd1 _20042_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16939__A _16939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _09800_/A _09784_/B vssd1 vssd1 vccd1 vccd1 _09784_/Y sky130_fd_sc_hd__nor2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11339__S1 _09658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09841__A _09841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18041__A1 _12414_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__S1 _10010_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16674__A _16674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12707__A _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09218_ _19890_/Q _19889_/Q vssd1 vssd1 vccd1 vccd1 _09349_/B sky130_fd_sc_hd__or2_1
XANTENNA__09288__A _12935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10490_ _10490_/A _10490_/B vssd1 vssd1 vccd1 vccd1 _10490_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12160_ _12160_/A _12160_/B vssd1 vssd1 vccd1 vccd1 _12161_/A sky130_fd_sc_hd__and2_2
XFILLER_107_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11111_ _18671_/Q _19166_/Q _11305_/S vssd1 vssd1 vccd1 vccd1 _11111_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_2_2_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12091_ _17180_/A _12092_/C _19828_/Q vssd1 vssd1 vccd1 vccd1 _12091_/Y sky130_fd_sc_hd__a21oi_1
X_11042_ _11046_/A _11042_/B vssd1 vssd1 vccd1 vccd1 _11042_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13972__S _13972_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16849__A _16946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15850_ _15850_/A vssd1 vssd1 vccd1 vccd1 _19356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input20_A io_dbus_rdata[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ _14801_/A vssd1 vssd1 vccd1 vccd1 _18953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _15781_/A vssd1 vssd1 vccd1 vccd1 _19344_/D sky130_fd_sc_hd__clkbuf_1
X_12993_ _19850_/Q _12992_/X _12695_/A _19817_/Q vssd1 vssd1 vccd1 vccd1 _12993_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17520_ _17798_/A vssd1 vssd1 vccd1 vccd1 _18054_/A sky130_fd_sc_hd__clkbuf_2
X_14732_ _14732_/A vssd1 vssd1 vccd1 vccd1 _18918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11944_ _19323_/D _11665_/B _11943_/Y _12155_/B vssd1 vssd1 vccd1 vccd1 _11944_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15899__S _15901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _17451_/A vssd1 vssd1 vccd1 vccd1 _17899_/B sky130_fd_sc_hd__buf_2
X_14663_ _14663_/A vssd1 vssd1 vccd1 vccd1 _14663_/X sky130_fd_sc_hd__clkbuf_2
X_11875_ _19821_/Q vssd1 vssd1 vccd1 vccd1 _17162_/A sky130_fd_sc_hd__inv_2
XFILLER_55_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output107_A _09188_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _13259_/X _19559_/Q _16404_/S vssd1 vssd1 vccd1 vccd1 _16403_/A sky130_fd_sc_hd__mux2_1
X_10826_ _18804_/Q _19139_/Q _10826_/S vssd1 vssd1 vccd1 vccd1 _10826_/X sky130_fd_sc_hd__mux2_1
X_13614_ _13744_/S vssd1 vssd1 vccd1 vccd1 _13631_/S sky130_fd_sc_hd__buf_2
X_17382_ _17382_/A _17382_/B _17382_/C vssd1 vssd1 vccd1 vccd1 _17382_/X sky130_fd_sc_hd__and3_1
X_14594_ _14592_/X _18869_/Q _14606_/S vssd1 vssd1 vccd1 vccd1 _14595_/A sky130_fd_sc_hd__mux2_1
X_19121_ _19313_/CLK _19121_/D vssd1 vssd1 vccd1 vccd1 _19121_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_2_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16333_ _16332_/A _16332_/C _13428_/A vssd1 vssd1 vccd1 vccd1 _16333_/Y sky130_fd_sc_hd__o21ai_1
X_10757_ _10757_/A _10757_/B vssd1 vssd1 vccd1 vccd1 _10757_/Y sky130_fd_sc_hd__nor2_1
X_13545_ _19805_/Q vssd1 vssd1 vccd1 vccd1 _16708_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14308__S _14308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11521__A _11538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19052_ _19406_/CLK _19052_/D vssd1 vssd1 vccd1 vccd1 _19052_/Q sky130_fd_sc_hd__dfxtp_1
X_16264_ _16264_/A vssd1 vssd1 vccd1 vccd1 _19525_/D sky130_fd_sc_hd__clkbuf_1
X_13476_ _16347_/B _13491_/C vssd1 vssd1 vccd1 vccd1 _13476_/Y sky130_fd_sc_hd__xnor2_1
X_10688_ _19368_/Q _18982_/Q _19432_/Q _18551_/Q _10614_/X _10682_/X vssd1 vssd1 vccd1
+ vccd1 _10689_/B sky130_fd_sc_hd__mux4_1
X_18003_ _17560_/A _17995_/Y _18002_/X _17966_/Y vssd1 vssd1 vccd1 vccd1 _18003_/X
+ sky130_fd_sc_hd__a31o_1
X_12427_ _12427_/A vssd1 vssd1 vccd1 vccd1 _18046_/A sky130_fd_sc_hd__buf_2
X_15215_ _15215_/A vssd1 vssd1 vccd1 vccd1 _15215_/X sky130_fd_sc_hd__clkbuf_2
X_16195_ _16195_/A vssd1 vssd1 vccd1 vccd1 _19510_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10137__A _10137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11040__C1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12358_ _12358_/A _18012_/B vssd1 vssd1 vccd1 vccd1 _12359_/B sky130_fd_sc_hd__nand2_1
X_15146_ _15146_/A vssd1 vssd1 vccd1 vccd1 _19104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11309_ _18571_/Q _18832_/Q _18731_/Q _19066_/Q _11129_/X _11115_/A vssd1 vssd1 vccd1
+ vccd1 _11309_/X sky130_fd_sc_hd__mux4_2
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15077_ _14596_/X _19072_/Q _15083_/S vssd1 vssd1 vccd1 vccd1 _15078_/A sky130_fd_sc_hd__mux2_1
X_19954_ _19954_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 _19954_/Q sky130_fd_sc_hd__dfxtp_1
X_12289_ _12263_/A _12288_/C _12339_/B vssd1 vssd1 vccd1 vccd1 _12290_/C sky130_fd_sc_hd__a21o_1
XFILLER_99_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12135__A2 _12649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ _14028_/A vssd1 vssd1 vccd1 vccd1 _18645_/D sky130_fd_sc_hd__clkbuf_1
X_18905_ _19204_/CLK _18905_/D vssd1 vssd1 vccd1 vccd1 _18905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19885_ _20044_/CLK _19885_/D vssd1 vssd1 vccd1 vccd1 _19885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18836_ _18836_/CLK _18836_/D vssd1 vssd1 vccd1 vccd1 _18836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18767_ _19486_/CLK _18767_/D vssd1 vssd1 vccd1 vccd1 _18767_/Q sky130_fd_sc_hd__dfxtp_1
X_15979_ _15979_/A vssd1 vssd1 vccd1 vccd1 _19414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17718_ _17679_/Y _17604_/B _17741_/S vssd1 vssd1 vccd1 vccd1 _17871_/A sky130_fd_sc_hd__mux2_1
X_18698_ _19952_/CLK _18698_/D vssd1 vssd1 vccd1 vccd1 _18698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11415__B _12656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17649_ _17649_/A vssd1 vssd1 vccd1 vccd1 _17800_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19319_ _19481_/CLK _19319_/D vssd1 vssd1 vccd1 vccd1 _19319_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12071__A1 _18349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14218__S _14218_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16433__S _16437_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09775__B1 _09479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09836__A _10367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15049__S _15055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11009__S0 _10937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12262__A _14477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09905_ _09822_/X _09904_/X _10256_/A vssd1 vssd1 vccd1 vccd1 _09905_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17772__B _17772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18262__A1 _19606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20025_ _20049_/CLK _20025_/D vssd1 vssd1 vccd1 vccd1 _20025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09836_ _10367_/S vssd1 vssd1 vccd1 vccd1 _09901_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10232__S1 _09874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09767_ _18791_/Q _19062_/Q _19286_/Q _19030_/Q _09763_/S _09526_/A vssd1 vssd1 vccd1
+ vccd1 _09767_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _18666_/Q _19257_/Q _19419_/Q _18634_/Q _09655_/X _09727_/A vssd1 vssd1 vccd1
+ vccd1 _09699_/B sky130_fd_sc_hd__mux4_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14917__A _18299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11660_ _17391_/B _17346_/A vssd1 vssd1 vccd1 vccd1 _11661_/A sky130_fd_sc_hd__and2_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09689__S0 _09726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10611_ _10805_/A vssd1 vssd1 vccd1 vccd1 _11362_/A sky130_fd_sc_hd__clkbuf_2
X_11591_ _11561_/X _11563_/Y _11564_/X _11565_/Y _11590_/X vssd1 vssd1 vccd1 vccd1
+ _11591_/X sky130_fd_sc_hd__a221o_1
X_13330_ _13324_/X _13328_/X _13329_/X vssd1 vssd1 vccd1 vccd1 _15257_/A sky130_fd_sc_hd__o21a_4
X_10542_ _10323_/A _10535_/X _10537_/Y _10541_/Y _09740_/A vssd1 vssd1 vccd1 vccd1
+ _10542_/X sky130_fd_sc_hd__o311a_2
XANTENNA__17947__B _17949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13261_ _13261_/A vssd1 vssd1 vccd1 vccd1 _18482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10473_ _10478_/A _10469_/X _10472_/X _10307_/X vssd1 vssd1 vccd1 vccd1 _10473_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15000_ _19038_/Q _14385_/X _15000_/S vssd1 vssd1 vccd1 vccd1 _15001_/A sky130_fd_sc_hd__mux2_1
X_12212_ _13591_/A vssd1 vssd1 vccd1 vccd1 _12212_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11022__C1 _09601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13192_ _13191_/A _13214_/C _13038_/A vssd1 vssd1 vccd1 vccd1 _13192_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input68_A io_irq_spi_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12143_ _12143_/A _17451_/A vssd1 vssd1 vccd1 vccd1 _12172_/A sky130_fd_sc_hd__nor2_1
XANTENNA__17963__A _17976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10471__S1 _10462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16951_ _17052_/A vssd1 vssd1 vccd1 vccd1 _16993_/A sky130_fd_sc_hd__clkbuf_2
X_12074_ _12074_/A _17866_/A vssd1 vssd1 vccd1 vccd1 _12080_/A sky130_fd_sc_hd__xor2_1
XFILLER_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15902_ _15902_/A vssd1 vssd1 vccd1 vccd1 _19380_/D sky130_fd_sc_hd__clkbuf_1
X_11025_ _11025_/A _11025_/B vssd1 vssd1 vccd1 vccd1 _11025_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18253__A1 _19602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19670_ _19671_/CLK _19670_/D vssd1 vssd1 vccd1 vccd1 _19670_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11876__A1 _19820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10223__S1 _09858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16882_ _16922_/C _16888_/D vssd1 vssd1 vccd1 vccd1 _16884_/B sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_3_6_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18621_ _19406_/CLK _18621_/D vssd1 vssd1 vccd1 vccd1 _18621_/Q sky130_fd_sc_hd__dfxtp_1
X_15833_ _15818_/X _18466_/Q _15819_/Y _13568_/X _15832_/X vssd1 vssd1 vccd1 vccd1
+ _15833_/X sky130_fd_sc_hd__a32o_2
XANTENNA__13078__B1 _12756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11516__A _11520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18552_ _18845_/CLK _18552_/D vssd1 vssd1 vccd1 vccd1 _18552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09916__S1 _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15764_ _15764_/A vssd1 vssd1 vccd1 vccd1 _15764_/Y sky130_fd_sc_hd__inv_2
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12976_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09297__A2 _11809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17503_ _12574_/A _11764_/C _17507_/S vssd1 vssd1 vccd1 vccd1 _17503_/X sky130_fd_sc_hd__mux2_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _14737_/A vssd1 vssd1 vccd1 vccd1 _14724_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_18_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _19063_/CLK _18483_/D vssd1 vssd1 vccd1 vccd1 _18483_/Q sky130_fd_sc_hd__dfxtp_1
X_11927_ _17594_/A _17749_/A vssd1 vssd1 vccd1 vccd1 _11990_/C sky130_fd_sc_hd__or2_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15695_ _13580_/X _15693_/X _15694_/Y _13577_/A _18443_/Q vssd1 vssd1 vccd1 vccd1
+ _17166_/A sky130_fd_sc_hd__a32oi_4
XFILLER_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15422__S _15428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17434_ _12673_/B _12614_/B _17549_/A vssd1 vssd1 vccd1 vccd1 _17434_/X sky130_fd_sc_hd__mux2_1
X_14646_ _14646_/A vssd1 vssd1 vccd1 vccd1 _18885_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _19961_/Q _11135_/X _11966_/A vssd1 vssd1 vccd1 vccd1 _17418_/A sky130_fd_sc_hd__mux2_2
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10809_ _19108_/Q _18874_/Q _19556_/Q _19204_/Q _10073_/X _09957_/A vssd1 vssd1 vccd1
+ vccd1 _10810_/B sky130_fd_sc_hd__mux4_2
X_17365_ _17365_/A vssd1 vssd1 vccd1 vccd1 _19888_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11487__S0 _09532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14038__S _14046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _11789_/A _11789_/B _11789_/C _11789_/D vssd1 vssd1 vccd1 vccd1 _11790_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14577_ _14676_/S vssd1 vssd1 vccd1 vccd1 _14590_/S sky130_fd_sc_hd__buf_2
XFILLER_41_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19104_ _19394_/CLK _19104_/D vssd1 vssd1 vccd1 vccd1 _19104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16316_ _19534_/Q _16300_/X _16314_/X _16315_/X vssd1 vssd1 vccd1 vccd1 _19534_/D
+ sky130_fd_sc_hd__o22a_1
X_13528_ _19736_/Q _13341_/A _12810_/Y _19704_/Q _13527_/X vssd1 vssd1 vccd1 vccd1
+ _13528_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11261__C1 _10941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17296_ _15784_/X _19871_/Q _17302_/S vssd1 vssd1 vccd1 vccd1 _17297_/A sky130_fd_sc_hd__mux2_1
X_19035_ _19485_/CLK _19035_/D vssd1 vssd1 vccd1 vccd1 _19035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16247_ _16247_/A vssd1 vssd1 vccd1 vccd1 _19522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13459_ _19951_/Q vssd1 vssd1 vccd1 vccd1 _16347_/A sky130_fd_sc_hd__buf_2
XFILLER_133_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13553__A1 _13600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput104 _09209_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[1] sky130_fd_sc_hd__buf_2
X_16178_ _19503_/Q _14637_/A _16178_/S vssd1 vssd1 vccd1 vccd1 _16179_/A sky130_fd_sc_hd__mux2_1
Xoutput115 _12651_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[15] sky130_fd_sc_hd__buf_2
XFILLER_142_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput126 _12663_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[25] sky130_fd_sc_hd__buf_2
Xoutput137 _12638_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[6] sky130_fd_sc_hd__buf_2
XANTENNA__13178__A _15225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput148 _12220_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[15] sky130_fd_sc_hd__buf_2
X_15129_ _14672_/X _19096_/Q _15131_/S vssd1 vssd1 vccd1 vccd1 _15130_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput159 _12472_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[25] sky130_fd_sc_hd__buf_2
XFILLER_114_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19937_ _19954_/CLK hold13/X vssd1 vssd1 vccd1 vccd1 _19937_/Q sky130_fd_sc_hd__dfxtp_1
X_19868_ _19873_/CLK _19868_/D vssd1 vssd1 vccd1 vccd1 _19868_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12810__A _17247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ _09621_/A vssd1 vssd1 vccd1 vccd1 _09622_/A sky130_fd_sc_hd__buf_4
XFILLER_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18819_ _19058_/CLK _18819_/D vssd1 vssd1 vccd1 vccd1 _18819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19799_ _19803_/CLK _19799_/D vssd1 vssd1 vccd1 vccd1 _19799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09552_ _18967_/Q vssd1 vssd1 vccd1 vccd1 _11116_/A sky130_fd_sc_hd__inv_2
XANTENNA__12816__B1 _12853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ _11014_/A vssd1 vssd1 vccd1 vccd1 _11489_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14737__A _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17507__A0 _12553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16163__S _16167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09843__S0 _09904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09285__B _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_103_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13816__A _13832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15507__S _15511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11858__A1 _11135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16246__A0 _19522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20008_ _20020_/CLK _20008_/D vssd1 vssd1 vccd1 vccd1 _20008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09819_ _19123_/Q _18889_/Q _19571_/Q _19219_/Q _09812_/X _10148_/A vssd1 vssd1 vccd1
+ vccd1 _09819_/X sky130_fd_sc_hd__mux4_2
XFILLER_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12830_ _13591_/A _12829_/X _12855_/B _18413_/A vssd1 vssd1 vccd1 vccd1 _17129_/S
+ sky130_fd_sc_hd__a31oi_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12807__B1 _13560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12761_ _19867_/Q _13560_/A _13562_/A _19531_/Q _12760_/X vssd1 vssd1 vccd1 vccd1
+ _12761_/X sky130_fd_sc_hd__a221o_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14500_ _14828_/A _18412_/B vssd1 vssd1 vccd1 vccd1 _18831_/D sky130_fd_sc_hd__nor2_4
XFILLER_43_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _17581_/S _11928_/A _11712_/C vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__and3_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _15502_/A vssd1 vssd1 vccd1 vccd1 _15489_/S sky130_fd_sc_hd__buf_2
X_12692_ _12692_/A vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14431_ _18813_/Q _14430_/X _14434_/S vssd1 vssd1 vccd1 vccd1 _14432_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12035__A1 _12855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11643_/A vssd1 vssd1 vccd1 vccd1 _11651_/C sky130_fd_sc_hd__inv_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11896__A2_N _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17150_ _19817_/Q _17229_/A vssd1 vssd1 vccd1 vccd1 _17150_/X sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_28_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14362_ _14362_/A vssd1 vssd1 vccd1 vccd1 _18791_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_opt_1_0_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_11574_ _11574_/A vssd1 vssd1 vccd1 vccd1 _11574_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_13_0_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 io_dbus_rdata[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_2
X_16101_ _16101_/A vssd1 vssd1 vccd1 vccd1 _19468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 io_dbus_rdata[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_4
Xinput39 io_ibus_inst[14] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_2
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10525_ _18651_/Q _19242_/Q _19404_/Q _18619_/Q _10509_/S _10461_/A vssd1 vssd1 vccd1
+ vccd1 _10526_/B sky130_fd_sc_hd__mux4_1
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13313_ _19942_/Q vssd1 vssd1 vccd1 vccd1 _16301_/A sky130_fd_sc_hd__clkbuf_2
X_17081_ _17089_/A _17081_/B _17081_/C vssd1 vssd1 vccd1 vccd1 _19788_/D sky130_fd_sc_hd__nor3_1
X_14293_ _14293_/A vssd1 vssd1 vccd1 vccd1 _18761_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10692__S1 _10691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16073__S _16073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16032_ _13331_/X _19438_/Q _16034_/S vssd1 vssd1 vccd1 vccd1 _16033_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09476__A _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13244_ _19719_/Q vssd1 vssd1 vccd1 vccd1 _16865_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10456_ _19911_/Q vssd1 vssd1 vccd1 vccd1 _10456_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11546__B1 _12662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12614__B _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13175_ _13175_/A vssd1 vssd1 vccd1 vccd1 _13175_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10387_ _09616_/A _10376_/X _10386_/X _09623_/A _19912_/Q vssd1 vssd1 vccd1 vccd1
+ _11415_/A sky130_fd_sc_hd__a32o_2
X_12126_ _16226_/A vssd1 vssd1 vccd1 vccd1 _12127_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17983_ _17995_/A _17983_/B vssd1 vssd1 vccd1 vccd1 _17983_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15417__S _15417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19722_ _19737_/CLK _19722_/D vssd1 vssd1 vccd1 vccd1 _19722_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13726__A _15286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16934_ _19740_/Q _16965_/C _16833_/X vssd1 vssd1 vccd1 vccd1 _16935_/B sky130_fd_sc_hd__o21ai_1
X_12057_ _11870_/C _12088_/B _12056_/A vssd1 vssd1 vccd1 vccd1 _12057_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11008_ _18769_/Q _19040_/Q _19264_/Q _19008_/Q _10893_/X _09512_/A vssd1 vssd1 vccd1
+ vccd1 _11008_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19653_ _19789_/CLK _19653_/D vssd1 vssd1 vccd1 vccd1 _19653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16865_ _16865_/A _19718_/Q _16868_/C _16865_/D vssd1 vssd1 vccd1 vccd1 _16920_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_19_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18604_ _19485_/CLK _18604_/D vssd1 vssd1 vccd1 vccd1 _18604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15816_ _15815_/X _19350_/Q _15835_/S vssd1 vssd1 vccd1 vccd1 _15817_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19584_ _19966_/CLK _19584_/D vssd1 vssd1 vccd1 vccd1 _19584_/Q sky130_fd_sc_hd__dfxtp_1
X_16796_ _16818_/A _16798_/B vssd1 vssd1 vccd1 vccd1 _16796_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18535_ _19512_/CLK _18535_/D vssd1 vssd1 vccd1 vccd1 _18535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _15746_/X _19338_/Q _15747_/S vssd1 vssd1 vccd1 vccd1 _15748_/A sky130_fd_sc_hd__mux2_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _17861_/A vssd1 vssd1 vccd1 vccd1 _12959_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18466_ _19952_/CLK _18466_/D vssd1 vssd1 vccd1 vccd1 _18466_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15678_ _16268_/A vssd1 vssd1 vccd1 vccd1 _15814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17417_ _17411_/X _17413_/X _17500_/S vssd1 vssd1 vccd1 vccd1 _17417_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14629_ _14628_/X _18880_/Q _14638_/S vssd1 vssd1 vccd1 vccd1 _14630_/A sky130_fd_sc_hd__mux2_1
X_18397_ _18401_/A vssd1 vssd1 vccd1 vccd1 _18426_/A sky130_fd_sc_hd__clkbuf_2
X_17348_ _17355_/A _17348_/B vssd1 vssd1 vccd1 vccd1 _17349_/A sky130_fd_sc_hd__and2_1
XFILLER_174_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17279_ _17279_/A vssd1 vssd1 vccd1 vccd1 _19863_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12805__A _12837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19018_ _19500_/CLK _19018_/D vssd1 vssd1 vccd1 vccd1 _19018_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13526__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10325__A _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14231__S _14235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__A _19606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10512__A1 _10294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09604_ _09604_/A vssd1 vssd1 vccd1 vccd1 _09605_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10060__A _11399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09535_ _10509_/S vssd1 vssd1 vccd1 vccd1 _10382_/A sky130_fd_sc_hd__buf_2
XANTENNA__12265__A1 _19531_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13462__B1 _13205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09466_ _13316_/A _09419_/X _09465_/X vssd1 vssd1 vccd1 vccd1 _18931_/D sky130_fd_sc_hd__o21ai_1
XFILLER_24_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15997__S _16001_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09397_ _12711_/A _12689_/B _09397_/C vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_174_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19831_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17900__B1 _17607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13310__S _13358_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _19376_/Q _18990_/Q _19440_/Q _18559_/Q _10302_/X _09817_/A vssd1 vssd1 vccd1
+ vccd1 _10311_/B sky130_fd_sc_hd__mux4_1
XFILLER_138_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11290_ _19357_/Q _18971_/Q _19421_/Q _18540_/Q _11329_/S _10978_/A vssd1 vssd1 vccd1
+ vccd1 _11291_/B sky130_fd_sc_hd__mux4_1
XFILLER_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_189_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _20018_/CLK sky130_fd_sc_hd__clkbuf_16
X_10241_ _10241_/A _10241_/B vssd1 vssd1 vccd1 vccd1 _11552_/A sky130_fd_sc_hd__nor2_1
XFILLER_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14930__A _14987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16467__B1 _16455_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10172_ _10184_/A _10172_/B vssd1 vssd1 vccd1 vccd1 _10172_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15745__B _17191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17018__A _17066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19555_/CLK sky130_fd_sc_hd__clkbuf_16
X_14980_ _14980_/A vssd1 vssd1 vccd1 vccd1 _19029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13931_ _18603_/Q _13608_/X _13939_/S vssd1 vssd1 vccd1 vccd1 _13932_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17960__B _17960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16650_ _19657_/Q _16647_/B _16649_/Y vssd1 vssd1 vccd1 vccd1 _19657_/D sky130_fd_sc_hd__o21a_1
X_13862_ _13862_/A vssd1 vssd1 vccd1 vccd1 _18572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15601_ _15601_/A vssd1 vssd1 vccd1 vccd1 _19294_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_127_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19395_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12813_ _12813_/A _12813_/B vssd1 vssd1 vccd1 vccd1 _12814_/B sky130_fd_sc_hd__nor2_4
XFILLER_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16581_ _19633_/Q _16582_/C _19634_/Q vssd1 vssd1 vccd1 vccd1 _16583_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13793_ _14618_/A vssd1 vssd1 vccd1 vccd1 _13793_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18320_ _20007_/Q _18310_/X _18319_/X _18317_/X vssd1 vssd1 vccd1 vccd1 _20007_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ _15532_/A vssd1 vssd1 vccd1 vccd1 _19263_/D sky130_fd_sc_hd__clkbuf_1
X_12744_ _16820_/A vssd1 vssd1 vccd1 vccd1 _18281_/B sky130_fd_sc_hd__buf_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12008__A1 _19522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18251_ _19980_/Q _12416_/A _18253_/S vssd1 vssd1 vccd1 vccd1 _18252_/A sky130_fd_sc_hd__mux2_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _19233_/Q _15222_/X _15467_/S vssd1 vssd1 vccd1 vccd1 _15464_/A sky130_fd_sc_hd__mux2_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12675_/A vssd1 vssd1 vccd1 vccd1 _12675_/X sky130_fd_sc_hd__buf_8
X_17202_ _12741_/X _17197_/X _17199_/X _17201_/X vssd1 vssd1 vccd1 vccd1 _19833_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14414_ _14618_/A vssd1 vssd1 vccd1 vccd1 _14414_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11626_ _11785_/A _11786_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _11682_/A sky130_fd_sc_hd__nor3b_1
X_18182_ _18182_/A vssd1 vssd1 vccd1 vccd1 _19949_/D sky130_fd_sc_hd__clkbuf_1
X_15394_ _15394_/A vssd1 vssd1 vccd1 vccd1 _19202_/D sky130_fd_sc_hd__clkbuf_1
X_17133_ _18413_/A vssd1 vssd1 vccd1 vccd1 _17138_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14345_ _14345_/A vssd1 vssd1 vccd1 vccd1 _18783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11557_ _11560_/A _11563_/A _11560_/C _10460_/A vssd1 vssd1 vccd1 vccd1 _11557_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ _11562_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _11563_/A sky130_fd_sc_hd__or2_1
X_17064_ _17089_/A hold19/A _17064_/C vssd1 vssd1 vccd1 vccd1 _19782_/D sky130_fd_sc_hd__nor3_1
X_14276_ _14276_/A vssd1 vssd1 vccd1 vccd1 _18753_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output99_A _11940_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11488_ _18601_/Q _18862_/Q _18761_/Q _19096_/Q _09967_/A _09513_/A vssd1 vssd1 vccd1
+ vccd1 _11489_/B sky130_fd_sc_hd__mux4_1
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16015_ _13219_/X _19430_/Q _16023_/S vssd1 vssd1 vccd1 vccd1 _16016_/A sky130_fd_sc_hd__mux2_1
X_10439_ _18813_/Q _19148_/Q _10439_/S vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__mux2_1
X_13227_ _13224_/Y _13254_/C _13226_/X _13418_/A vssd1 vssd1 vccd1 vccd1 _13227_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_170_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13158_ _19746_/Q _12692_/X _12696_/X _17176_/A _12714_/X vssd1 vssd1 vccd1 vccd1
+ _13158_/X sky130_fd_sc_hd__a221o_1
XFILLER_3_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11090__S1 _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _12050_/A _12079_/A _12081_/B vssd1 vssd1 vccd1 vccd1 _12109_/Y sky130_fd_sc_hd__a21oi_1
X_13089_ _15212_/A vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__clkbuf_1
X_17966_ _17966_/A _17966_/B vssd1 vssd1 vccd1 vccd1 _17966_/Y sky130_fd_sc_hd__nand2_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19705_ _19721_/CLK _19705_/D vssd1 vssd1 vccd1 vccd1 _19705_/Q sky130_fd_sc_hd__dfxtp_1
X_16917_ _19737_/Q _16930_/D vssd1 vssd1 vccd1 vccd1 _16919_/B sky130_fd_sc_hd__nor2_1
XFILLER_66_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12495__B2 _11771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17897_ _17985_/A vssd1 vssd1 vccd1 vccd1 _17945_/A sky130_fd_sc_hd__buf_2
XFILLER_77_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19636_ _19718_/CLK _19636_/D vssd1 vssd1 vccd1 vccd1 _19636_/Q sky130_fd_sc_hd__dfxtp_1
X_16848_ _19715_/Q _19714_/Q _16848_/C _16848_/D vssd1 vssd1 vccd1 vccd1 _16857_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_19_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19567_ _19570_/CLK _19567_/D vssd1 vssd1 vccd1 vccd1 _19567_/Q sky130_fd_sc_hd__dfxtp_1
X_16779_ _16898_/A vssd1 vssd1 vccd1 vccd1 _16874_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13444__B1 _13205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ _09320_/A _09320_/B _09320_/C _09319_/X vssd1 vssd1 vccd1 vccd1 _09751_/C
+ sky130_fd_sc_hd__or4b_2
X_18518_ _18777_/CLK _18518_/D vssd1 vssd1 vccd1 vccd1 _18518_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11704__A _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19498_ _19498_/CLK _19498_/D vssd1 vssd1 vccd1 vccd1 _19498_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17186__A1 _12854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18383__B1 _18374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19497_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09251_ _17382_/A _17393_/A vssd1 vssd1 vccd1 vccd1 _17336_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18449_ _19938_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09182_ _09271_/B vssd1 vssd1 vccd1 vccd1 _11786_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10408__S1 _10440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16441__S _16441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18222__A _18268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15057__S _15059_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15672__A1 _11187_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14896__S _14900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19314_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09518_ _10510_/A vssd1 vssd1 vccd1 vccd1 _09841_/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_59_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19416_/CLK sky130_fd_sc_hd__clkbuf_16
X_10790_ _10790_/A _10790_/B vssd1 vssd1 vccd1 vccd1 _10790_/Y sky130_fd_sc_hd__nor2_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _11723_/B _09449_/B _09453_/B vssd1 vssd1 vccd1 vccd1 _11790_/A sky130_fd_sc_hd__or3_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ _12460_/A _18046_/B vssd1 vssd1 vccd1 vccd1 _12460_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _11411_/A _12651_/A vssd1 vssd1 vccd1 vccd1 _11567_/A sky130_fd_sc_hd__and2_1
XFILLER_165_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12391_ _12391_/A _12391_/B vssd1 vssd1 vccd1 vccd1 _12391_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__14136__S _14142_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14130_ _14130_/A vssd1 vssd1 vccd1 vccd1 _18690_/D sky130_fd_sc_hd__clkbuf_1
X_11342_ _11342_/A _11342_/B vssd1 vssd1 vccd1 vccd1 _11342_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14061_ _14061_/A vssd1 vssd1 vccd1 vccd1 _18660_/D sky130_fd_sc_hd__clkbuf_1
X_11273_ _19453_/Q _19291_/Q _18700_/Q _18470_/Q _11002_/A _10880_/A vssd1 vssd1 vccd1
+ vccd1 _11274_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10224_ _10229_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10224_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13012_ _15061_/A _14917_/B vssd1 vssd1 vccd1 vccd1 _14151_/B sky130_fd_sc_hd__nand2_2
XANTENNA__09754__A _10065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input50_A io_ibus_inst[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11072__S1 _10083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17820_ _17820_/A _17820_/B vssd1 vssd1 vccd1 vccd1 _17820_/X sky130_fd_sc_hd__or2_1
X_10155_ _19475_/Q _19313_/Q _18722_/Q _18492_/Q _10244_/S _10148_/A vssd1 vssd1 vccd1
+ vccd1 _10156_/B sky130_fd_sc_hd__mux4_1
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17751_ _17697_/X _17748_/X _17750_/Y _17705_/X vssd1 vssd1 vccd1 vccd1 _17751_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14963_ _14974_/A vssd1 vssd1 vccd1 vccd1 _14972_/S sky130_fd_sc_hd__buf_2
X_10086_ _18790_/Q _19061_/Q _19285_/Q _19029_/Q _10081_/X _10691_/A vssd1 vssd1 vccd1
+ vccd1 _10086_/X sky130_fd_sc_hd__mux4_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output137_A _12638_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15491__A _15502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16702_ _19793_/Q _19795_/Q _19794_/Q _17090_/A vssd1 vssd1 vccd1 vccd1 _17098_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13914_ _13831_/X _18596_/Q _13922_/S vssd1 vssd1 vccd1 vccd1 _13915_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17404__A2 _12620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17682_ _17572_/X _17561_/X _17685_/S vssd1 vssd1 vccd1 vccd1 _17682_/X sky130_fd_sc_hd__mux2_1
X_14894_ _14644_/X _18991_/Q _14900_/S vssd1 vssd1 vccd1 vccd1 _14895_/A sky130_fd_sc_hd__mux2_1
X_19421_ _19727_/CLK _19421_/D vssd1 vssd1 vccd1 vccd1 _19421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16633_ _16636_/B _16636_/C _16624_/X vssd1 vssd1 vccd1 vccd1 _16633_/Y sky130_fd_sc_hd__a21oi_1
X_13845_ _13844_/X _18568_/Q _13845_/S vssd1 vssd1 vccd1 vccd1 _13846_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19352_ _19879_/CLK _19352_/D vssd1 vssd1 vccd1 vccd1 _19352_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11524__A _18302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16564_ _19628_/Q _19627_/Q _16564_/C vssd1 vssd1 vccd1 vccd1 _16566_/B sky130_fd_sc_hd__and3_1
X_13776_ _13776_/A vssd1 vssd1 vccd1 vccd1 _18546_/D sky130_fd_sc_hd__clkbuf_1
X_10988_ _10988_/A vssd1 vssd1 vccd1 vccd1 _10988_/X sky130_fd_sc_hd__clkbuf_2
X_18303_ _18341_/A vssd1 vssd1 vccd1 vccd1 _18303_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15515_ _19257_/Q _15298_/X _15515_/S vssd1 vssd1 vccd1 vccd1 _15516_/A sky130_fd_sc_hd__mux2_1
X_19283_ _19443_/CLK _19283_/D vssd1 vssd1 vccd1 vccd1 _19283_/Q sky130_fd_sc_hd__dfxtp_1
X_12727_ _13116_/A vssd1 vssd1 vccd1 vccd1 _12727_/X sky130_fd_sc_hd__clkbuf_2
X_16495_ _19642_/Q _19643_/Q _19645_/Q _19644_/Q vssd1 vssd1 vccd1 vccd1 _16612_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18234_ _19972_/Q _12338_/A _18242_/S vssd1 vssd1 vccd1 vccd1 _18235_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09929__A _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15446_ _15502_/A vssd1 vssd1 vccd1 vccd1 _15515_/S sky130_fd_sc_hd__buf_6
XFILLER_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12658_ _12664_/A vssd1 vssd1 vccd1 vccd1 _12663_/A sky130_fd_sc_hd__buf_8
XFILLER_129_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11609_ _11690_/B vssd1 vssd1 vccd1 vccd1 _17394_/B sky130_fd_sc_hd__clkbuf_2
X_18165_ _18165_/A vssd1 vssd1 vccd1 vccd1 _19941_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14046__S _14046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15377_ _15377_/A vssd1 vssd1 vccd1 vccd1 _19194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12589_ _12421_/X _12587_/X _12588_/Y _12131_/X vssd1 vssd1 vccd1 vccd1 _12589_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17116_ _17123_/A _17120_/C vssd1 vssd1 vccd1 vccd1 _17116_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14328_ _18776_/Q _13668_/X _14330_/S vssd1 vssd1 vccd1 vccd1 _14329_/A sky130_fd_sc_hd__mux2_1
X_18096_ _19921_/Q _18019_/X _18095_/X vssd1 vssd1 vccd1 vccd1 _19921_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17340__B2 _18302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13885__S _13889_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17047_ _17047_/A vssd1 vssd1 vccd1 vccd1 _17053_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14259_ _14281_/A vssd1 vssd1 vccd1 vccd1 _14268_/S sky130_fd_sc_hd__buf_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18998_ _19574_/CLK _18998_/D vssd1 vssd1 vccd1 vccd1 _18998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11418__B _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12468__A1 _19539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _17949_/A _17945_/B vssd1 vssd1 vccd1 vccd1 _17949_/X sky130_fd_sc_hd__or2b_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16603__B1 _16577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19619_ _19620_/CLK _19619_/D vssd1 vssd1 vccd1 vccd1 _19619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17159__A1 _19820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11979__B1 _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09303_ _09303_/A vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10877__S1 _10084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09234_ _09262_/A _09303_/A _11629_/A vssd1 vssd1 vccd1 vccd1 _17379_/B sky130_fd_sc_hd__a21oi_1
XFILLER_167_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14480__A _14831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11054__S1 _10083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12712__B _12837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09998_ _09998_/A vssd1 vssd1 vccd1 vccd1 _09998_/X sky130_fd_sc_hd__buf_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15515__S _15515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11960_ _11974_/A _12150_/B _11947_/Y _11959_/X vssd1 vssd1 vccd1 vccd1 _16458_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13408__A0 _19915_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ _10041_/A _10908_/Y _10910_/Y _10929_/A vssd1 vssd1 vccd1 vccd1 _10911_/X
+ sky130_fd_sc_hd__o211a_1
X_11891_ _11872_/Y _11874_/Y _11887_/X _11890_/X _16487_/A vssd1 vssd1 vccd1 vccd1
+ _11892_/B sky130_fd_sc_hd__o221ai_1
X_13630_ _14589_/A vssd1 vssd1 vccd1 vccd1 _13630_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10842_ _10730_/A _10841_/X _09976_/X vssd1 vssd1 vccd1 vccd1 _10842_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13561_ _13546_/B _13562_/A _13562_/B vssd1 vssd1 vccd1 vccd1 _13561_/Y sky130_fd_sc_hd__o21ai_1
X_10773_ _09748_/A _10762_/X _10771_/X _09755_/A _10772_/Y vssd1 vssd1 vccd1 vccd1
+ _12647_/A sky130_fd_sc_hd__o32a_4
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18127__A _18127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15300_ _15300_/A vssd1 vssd1 vccd1 vccd1 _19161_/D sky130_fd_sc_hd__clkbuf_1
X_12512_ _12512_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12512_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09749__A _09749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16280_ _19528_/Q _16279_/X _16280_/S vssd1 vssd1 vccd1 vccd1 _16281_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13492_ _16347_/B _13491_/C _19953_/Q vssd1 vssd1 vccd1 vccd1 _13492_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15231_ _15231_/A vssd1 vssd1 vccd1 vccd1 _15231_/X sky130_fd_sc_hd__clkbuf_2
X_12443_ _19841_/Q vssd1 vssd1 vccd1 vccd1 _17223_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11198__A1 _11204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12395__A0 _12391_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15162_ _15162_/A vssd1 vssd1 vccd1 vccd1 _19112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12374_ _12314_/X _12372_/Y _12419_/C _12218_/X vssd1 vssd1 vccd1 vccd1 _12374_/Y
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__10945__B2 _11250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14113_ _14113_/A vssd1 vssd1 vccd1 vccd1 _18682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11325_ _19098_/Q _18864_/Q _19546_/Q _19194_/Q _11030_/A _09658_/A vssd1 vssd1 vccd1
+ vccd1 _11326_/B sky130_fd_sc_hd__mux4_1
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15093_ _15093_/A vssd1 vssd1 vccd1 vccd1 _19079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19970_ _19971_/CLK _19970_/D vssd1 vssd1 vccd1 vccd1 _19970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18921_ _19449_/CLK _18921_/D vssd1 vssd1 vccd1 vccd1 _18921_/Q sky130_fd_sc_hd__dfxtp_1
X_14044_ _18653_/Q _13689_/X _14046_/S vssd1 vssd1 vccd1 vccd1 _14045_/A sky130_fd_sc_hd__mux2_1
X_11256_ _19099_/Q _18865_/Q _19547_/Q _19195_/Q _11003_/A _11059_/A vssd1 vssd1 vccd1
+ vccd1 _11257_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10158__C1 _09605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11045__S1 _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10207_ _10207_/A _10207_/B vssd1 vssd1 vccd1 vccd1 _10207_/X sky130_fd_sc_hd__or2_1
X_18852_ _19565_/CLK _18852_/D vssd1 vssd1 vccd1 vccd1 _18852_/Q sky130_fd_sc_hd__dfxtp_1
X_11187_ _19895_/Q vssd1 vssd1 vccd1 vccd1 _11187_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_151_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _11544_/A _11544_/B vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__nand2_1
X_17803_ _17674_/X _17677_/X _17803_/S vssd1 vssd1 vccd1 vccd1 _17803_/X sky130_fd_sc_hd__mux2_1
X_18783_ _19409_/CLK _18783_/D vssd1 vssd1 vccd1 vccd1 _18783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15995_ _13033_/X _19421_/Q _16001_/S vssd1 vssd1 vccd1 vccd1 _15996_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13734__A _15292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18035__C1 _17543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17734_ _11864_/A _17554_/B _18019_/A vssd1 vssd1 vccd1 vccd1 _17734_/Y sky130_fd_sc_hd__o21ai_1
X_14946_ _19014_/Q _14411_/X _14950_/S vssd1 vssd1 vccd1 vccd1 _14947_/A sky130_fd_sc_hd__mux2_1
X_10069_ _18694_/Q _19189_/Q _10812_/S vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17665_ _17888_/A vssd1 vssd1 vccd1 vccd1 _17666_/S sky130_fd_sc_hd__clkbuf_2
X_14877_ _14877_/A vssd1 vssd1 vccd1 vccd1 _18983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19404_ _19405_/CLK _19404_/D vssd1 vssd1 vccd1 vccd1 _19404_/Q sky130_fd_sc_hd__dfxtp_1
X_16616_ _16617_/B _16617_/C _16615_/Y vssd1 vssd1 vccd1 vccd1 _19646_/D sky130_fd_sc_hd__o21a_1
X_13828_ _14653_/A vssd1 vssd1 vccd1 vccd1 _13828_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17596_ _17966_/A _17596_/B vssd1 vssd1 vccd1 vccd1 _18072_/A sky130_fd_sc_hd__and2_1
XFILLER_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19335_ _19879_/CLK _19335_/D vssd1 vssd1 vccd1 vccd1 _19335_/Q sky130_fd_sc_hd__dfxtp_1
X_16547_ _19622_/Q _16547_/B _16547_/C vssd1 vssd1 vccd1 vccd1 _16548_/C sky130_fd_sc_hd__and3_1
X_13759_ _13758_/X _18541_/Q _13765_/S vssd1 vssd1 vccd1 vccd1 _13760_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10859__S1 _10014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17010__B1 _16860_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__A _09659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19266_ _19490_/CLK _19266_/D vssd1 vssd1 vccd1 vccd1 _19266_/Q sky130_fd_sc_hd__dfxtp_1
X_16478_ _12339_/B _16477_/X _12292_/X _12296_/X _16468_/X vssd1 vssd1 vccd1 vccd1
+ _19596_/D sky130_fd_sc_hd__o221a_1
X_18217_ _18217_/A vssd1 vssd1 vccd1 vccd1 _19964_/D sky130_fd_sc_hd__clkbuf_1
X_15429_ _15429_/A vssd1 vssd1 vccd1 vccd1 _19218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19197_ _19455_/CLK _19197_/D vssd1 vssd1 vccd1 vccd1 _19197_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_76_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12925__A2 _15799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18148_ _13191_/A _19966_/Q _18148_/S vssd1 vssd1 vccd1 vccd1 _18149_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18079_ _18079_/A _18079_/B vssd1 vssd1 vccd1 vccd1 _18079_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16930__D _16930_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09921_ _09616_/A _09911_/X _09920_/X _09623_/A _19917_/Q vssd1 vssd1 vccd1 vccd1
+ _10144_/A sky130_fd_sc_hd__a32o_2
XFILLER_160_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20041_ _20052_/CLK _20041_/D vssd1 vssd1 vccd1 vccd1 _20041_/Q sky130_fd_sc_hd__dfxtp_2
X_09852_ _09924_/S vssd1 vssd1 vccd1 vccd1 _09926_/S sky130_fd_sc_hd__clkbuf_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10333__A _10333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10795__S0 _10700_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _19126_/Q _18892_/Q _19574_/Q _19222_/Q _09724_/S _09688_/A vssd1 vssd1 vccd1
+ vccd1 _09784_/B sky130_fd_sc_hd__mux4_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17116__A _17123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10547__S0 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16955__A _16955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14475__A _18404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15070__S _15072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__A _09569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16355__A2 _15828_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09217_ _13163_/A vssd1 vssd1 vccd1 vccd1 _13316_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__17786__A _17792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10508__A _11562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ _11125_/A _11110_/B vssd1 vssd1 vccd1 vccd1 _11110_/X sky130_fd_sc_hd__or2_1
XFILLER_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12090_ _19525_/Q _12120_/A _12855_/A vssd1 vssd1 vccd1 vccd1 _12090_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11041_ _19362_/Q _18976_/Q _19426_/Q _18545_/Q _10914_/X _10969_/A vssd1 vssd1 vccd1
+ vccd1 _11042_/B sky130_fd_sc_hd__mux4_1
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18410__A _18412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10786__S0 _10048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14800_ _18953_/Q _14436_/X _14808_/S vssd1 vssd1 vccd1 vccd1 _14801_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17026__A _17046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _15778_/X _19344_/Q _15801_/S vssd1 vssd1 vccd1 vccd1 _15781_/A sky130_fd_sc_hd__mux2_1
X_12992_ _12992_/A vssd1 vssd1 vccd1 vccd1 _12992_/X sky130_fd_sc_hd__buf_2
XFILLER_76_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14731_ _18918_/Q _14443_/X _14735_/S vssd1 vssd1 vccd1 vccd1 _14732_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input13_A io_dbus_rdata[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11943_ _11974_/A _12240_/B vssd1 vssd1 vccd1 vccd1 _11943_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _17884_/B _17985_/B _17450_/S vssd1 vssd1 vccd1 vccd1 _17450_/X sky130_fd_sc_hd__mux2_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14662_/A vssd1 vssd1 vccd1 vccd1 _18890_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _19518_/Q _11782_/X _15719_/S vssd1 vssd1 vccd1 vccd1 _11874_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _16401_/A vssd1 vssd1 vccd1 vccd1 _19558_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _13719_/A vssd1 vssd1 vccd1 vccd1 _13744_/S sky130_fd_sc_hd__buf_6
XFILLER_38_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _10825_/A _10825_/B vssd1 vssd1 vccd1 vccd1 _10825_/X sky130_fd_sc_hd__and2_1
X_17381_ _17381_/A _17394_/B _17381_/C vssd1 vssd1 vccd1 vccd1 _17382_/C sky130_fd_sc_hd__and3_1
XFILLER_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14593_ _14676_/S vssd1 vssd1 vccd1 vccd1 _14606_/S sky130_fd_sc_hd__buf_2
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14385__A _14589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19120_ _19569_/CLK _19120_/D vssd1 vssd1 vccd1 vccd1 _19120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16332_ _16332_/A _19949_/Q _16332_/C vssd1 vssd1 vccd1 vccd1 _16338_/B sky130_fd_sc_hd__or3_1
X_13544_ _19673_/Q vssd1 vssd1 vccd1 vccd1 _16507_/B sky130_fd_sc_hd__clkbuf_2
X_10756_ _19109_/Q _18875_/Q _19557_/Q _19205_/Q _09647_/A _11387_/A vssd1 vssd1 vccd1
+ vccd1 _10757_/B sky130_fd_sc_hd__mux4_2
XFILLER_125_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10710__S0 _10753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19051_ _19051_/CLK _19051_/D vssd1 vssd1 vccd1 vccd1 _19051_/Q sky130_fd_sc_hd__dfxtp_1
X_16263_ _19525_/Q _16262_/X _16280_/S vssd1 vssd1 vccd1 vccd1 _16264_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13475_ _19952_/Q vssd1 vssd1 vccd1 vccd1 _16347_/B sky130_fd_sc_hd__buf_2
X_10687_ _09979_/X _10677_/X _10681_/X _10686_/X _10623_/A vssd1 vssd1 vccd1 vccd1
+ _10687_/X sky130_fd_sc_hd__a311o_2
X_18002_ _18002_/A _18002_/B _18002_/C _18002_/D vssd1 vssd1 vccd1 vccd1 _18002_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_127_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15214_ _15214_/A vssd1 vssd1 vccd1 vccd1 _19134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12426_ _12473_/A _12662_/B _12474_/A _12425_/X vssd1 vssd1 vccd1 vccd1 _12427_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12907__A2 _17122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16194_ _19510_/Q _14660_/A _16200_/S vssd1 vssd1 vccd1 vccd1 _16195_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10137__B _12666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15145_ _19104_/Q vssd1 vssd1 vccd1 vccd1 _15146_/A sky130_fd_sc_hd__clkbuf_1
X_12357_ _12358_/A _18012_/B vssd1 vssd1 vccd1 vccd1 _12390_/A sky130_fd_sc_hd__or2_2
XANTENNA__12633__A _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output81_A _12309_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11308_ _11482_/A _11305_/X _11307_/X vssd1 vssd1 vccd1 vccd1 _11308_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19953_ _19985_/CLK _19953_/D vssd1 vssd1 vccd1 vccd1 _19953_/Q sky130_fd_sc_hd__dfxtp_2
X_15076_ _15076_/A vssd1 vssd1 vccd1 vccd1 _19071_/D sky130_fd_sc_hd__clkbuf_1
X_12288_ _19595_/Q _19596_/Q _12288_/C vssd1 vssd1 vccd1 vccd1 _12365_/D sky130_fd_sc_hd__and3_1
XFILLER_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14027_ _18645_/Q _13655_/X _14035_/S vssd1 vssd1 vccd1 vccd1 _14028_/A sky130_fd_sc_hd__mux2_1
X_18904_ _19204_/CLK _18904_/D vssd1 vssd1 vccd1 vccd1 _18904_/Q sky130_fd_sc_hd__dfxtp_1
X_11239_ _11304_/A _11234_/X _11236_/X _11238_/X vssd1 vssd1 vccd1 vccd1 _11239_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_68_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19884_ _19892_/CLK _19884_/D vssd1 vssd1 vccd1 vccd1 _19884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18835_ _18836_/CLK _18835_/D vssd1 vssd1 vccd1 vccd1 _18835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10551__C1 _09718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15978_ _19414_/Q _15283_/X _15984_/S vssd1 vssd1 vccd1 vccd1 _15979_/A sky130_fd_sc_hd__mux2_1
X_18766_ _19488_/CLK _18766_/D vssd1 vssd1 vccd1 vccd1 _18766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14929_ _14929_/A vssd1 vssd1 vccd1 vccd1 _19006_/D sky130_fd_sc_hd__clkbuf_1
X_17717_ _17714_/X _17716_/X _17888_/A vssd1 vssd1 vccd1 vccd1 _17717_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14994__S _15000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18697_ _19556_/CLK _18697_/D vssd1 vssd1 vccd1 vccd1 _18697_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10854__B1 _10655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17648_ _17425_/X _17433_/X _17660_/S vssd1 vssd1 vccd1 vccd1 _17648_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17579_ _17476_/X _17495_/X _17590_/S vssd1 vssd1 vccd1 vccd1 _17579_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11712__A _17581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19318_ _19512_/CLK _19318_/D vssd1 vssd1 vccd1 vccd1 _19318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19249_ _19411_/CLK _19249_/D vssd1 vssd1 vccd1 vccd1 _19249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13639__A _14596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11009__S1 _09954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09904_ _18819_/Q _19154_/Q _09904_/S vssd1 vssd1 vccd1 vccd1 _09904_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10063__A _10063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20024_ _20027_/CLK _20024_/D vssd1 vssd1 vccd1 vccd1 _20024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09835_ _10559_/S vssd1 vssd1 vccd1 vccd1 _10367_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA_input5_A io_dbus_rdata[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10542__C1 _09740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _09762_/X _09764_/X _09765_/X _10166_/A _09479_/X vssd1 vssd1 vccd1 vccd1
+ _09771_/B sky130_fd_sc_hd__o221a_1
XFILLER_101_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09697_ _09699_/A _09689_/X _09696_/X vssd1 vssd1 vccd1 vccd1 _09697_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11193__S0 _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10937__S _10937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12718__A _12989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _19112_/Q _18878_/Q _19560_/Q _19208_/Q _10608_/X _10609_/X vssd1 vssd1 vccd1
+ vccd1 _10610_/X sky130_fd_sc_hd__mux4_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11590_ _11566_/X _11568_/Y _11569_/Y _11571_/Y _11589_/X vssd1 vssd1 vccd1 vccd1
+ _11590_/X sky130_fd_sc_hd__a2111o_1
XFILLER_10_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16328__A2 _16327_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _10544_/A _10538_/X _10540_/X vssd1 vssd1 vccd1 vccd1 _10541_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13260_ _18482_/Q _13259_/X _13278_/S vssd1 vssd1 vccd1 vccd1 _13261_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10472_ _10521_/A _10472_/B vssd1 vssd1 vccd1 vccd1 _10472_/X sky130_fd_sc_hd__or2_1
XFILLER_136_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12211_ _12204_/Y _12209_/X _12583_/S vssd1 vssd1 vccd1 vccd1 _12211_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09766__B2 _10166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14144__S _14146_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13191_ _13191_/A _13214_/C vssd1 vssd1 vccd1 vccd1 _13191_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15839__A1 _15818_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ _12143_/A _17451_/A vssd1 vssd1 vccd1 vccd1 _12144_/A sky130_fd_sc_hd__and2_1
XFILLER_124_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15764__A _15764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16950_ _16957_/B _16946_/B _16949_/Y vssd1 vssd1 vccd1 vccd1 _19744_/D sky130_fd_sc_hd__o21a_1
X_12073_ _12376_/A _12647_/A _12039_/C _12072_/X vssd1 vssd1 vccd1 vccd1 _17866_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_96_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10759__S0 _11449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15901_ _13433_/X _19380_/Q _15901_/S vssd1 vssd1 vccd1 vccd1 _15902_/A sky130_fd_sc_hd__mux2_1
X_11024_ _19104_/Q _18870_/Q _19552_/Q _19200_/Q _10903_/A _10974_/X vssd1 vssd1 vccd1
+ vccd1 _11025_/B sky130_fd_sc_hd__mux4_1
X_16881_ _16897_/A _16881_/B _16888_/D vssd1 vssd1 vccd1 vccd1 _19724_/D sky130_fd_sc_hd__nor3_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_24_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18620_ _19501_/CLK _18620_/D vssd1 vssd1 vccd1 vccd1 _18620_/Q sky130_fd_sc_hd__dfxtp_1
X_15832_ _13519_/X _09339_/A _18466_/Q vssd1 vssd1 vccd1 vccd1 _15832_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13078__B2 _19518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18551_ _19302_/CLK _18551_/D vssd1 vssd1 vccd1 vccd1 _18551_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11516__B _12669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15763_ _15763_/A vssd1 vssd1 vccd1 vccd1 _19341_/D sky130_fd_sc_hd__clkbuf_1
X_12975_ _18461_/Q _12973_/X _10144_/A _12969_/X vssd1 vssd1 vccd1 vccd1 _18461_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11628__A2 _17342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11184__S0 _11161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _14714_/A vssd1 vssd1 vccd1 vccd1 _18910_/D sky130_fd_sc_hd__clkbuf_1
X_17502_ _17497_/X _17500_/X _17686_/S vssd1 vssd1 vccd1 vccd1 _17502_/X sky130_fd_sc_hd__mux2_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _18845_/CLK _18482_/D vssd1 vssd1 vccd1 vccd1 _18482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11926_ _11926_/A vssd1 vssd1 vccd1 vccd1 _17772_/A sky130_fd_sc_hd__buf_2
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ _15818_/A _18443_/Q vssd1 vssd1 vccd1 vccd1 _15694_/Y sky130_fd_sc_hd__nand2_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17430_/X _17432_/X _17582_/S vssd1 vssd1 vccd1 vccd1 _17433_/X sky130_fd_sc_hd__mux2_1
X_14645_ _14644_/X _18885_/Q _14654_/S vssd1 vssd1 vccd1 vccd1 _14646_/A sky130_fd_sc_hd__mux2_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _11857_/A _17594_/A vssd1 vssd1 vccd1 vccd1 _11860_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__14319__S _14319_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12350__A1_N _12376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10808_ _10801_/X _10803_/X _10805_/X _10807_/X _09602_/A vssd1 vssd1 vccd1 vccd1
+ _10808_/X sky130_fd_sc_hd__a221o_2
X_17364_ _17373_/A _17364_/B vssd1 vssd1 vccd1 vccd1 _17365_/A sky130_fd_sc_hd__and2_1
X_14576_ _14657_/A vssd1 vssd1 vccd1 vccd1 _14676_/S sky130_fd_sc_hd__buf_4
X_11788_ _20028_/Q _18286_/A _18283_/A _12606_/D vssd1 vssd1 vccd1 vccd1 _11789_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_119_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16315_ _16315_/A _16315_/B _16315_/C vssd1 vssd1 vccd1 vccd1 _16315_/X sky130_fd_sc_hd__or3_4
X_19103_ _19293_/CLK _19103_/D vssd1 vssd1 vccd1 vccd1 _19103_/Q sky130_fd_sc_hd__dfxtp_1
X_13527_ _19672_/Q _13527_/B vssd1 vssd1 vccd1 vccd1 _13527_/X sky130_fd_sc_hd__and2_1
X_10739_ _09577_/A _10730_/X _10732_/X _10623_/A _10738_/X vssd1 vssd1 vccd1 vccd1
+ _10739_/X sky130_fd_sc_hd__a311o_1
X_17295_ _17295_/A vssd1 vssd1 vccd1 vccd1 _19870_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10148__A _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19034_ _19484_/CLK _19034_/D vssd1 vssd1 vccd1 vccd1 _19034_/Q sky130_fd_sc_hd__dfxtp_1
X_16246_ _19522_/Q _16245_/X _16252_/S vssd1 vssd1 vccd1 vccd1 _16247_/A sky130_fd_sc_hd__mux2_1
X_13458_ _19951_/Q _13460_/B vssd1 vssd1 vccd1 vccd1 _13491_/C sky130_fd_sc_hd__and2_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12409_ _12521_/A vssd1 vssd1 vccd1 vccd1 _12411_/A sky130_fd_sc_hd__inv_2
X_16177_ _16177_/A vssd1 vssd1 vccd1 vccd1 _19502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput105 _11673_/A vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[2] sky130_fd_sc_hd__buf_2
X_13389_ _19914_/Q _15782_/B _13483_/A vssd1 vssd1 vccd1 vccd1 _13389_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput116 _12653_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[16] sky130_fd_sc_hd__buf_2
Xoutput127 _12665_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[26] sky130_fd_sc_hd__buf_2
X_15128_ _15128_/A vssd1 vssd1 vccd1 vccd1 _19095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput138 _12639_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[7] sky130_fd_sc_hd__buf_2
Xoutput149 _12249_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[16] sky130_fd_sc_hd__buf_2
XFILLER_141_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15059_ _19065_/Q _14471_/X _15059_/S vssd1 vssd1 vccd1 vccd1 _15060_/A sky130_fd_sc_hd__mux2_1
X_19936_ _19954_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 _19936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12513__A0 _12509_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19867_ _19873_/CLK _19867_/D vssd1 vssd1 vccd1 vccd1 _19867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09620_ _09996_/A vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__buf_4
X_18818_ _19286_/CLK _18818_/D vssd1 vssd1 vccd1 vccd1 _18818_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10611__A _10805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19798_ _19803_/CLK _19798_/D vssd1 vssd1 vccd1 vccd1 _19798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09551_ _18698_/Q _19193_/Q _09763_/S vssd1 vssd1 vccd1 vccd1 _09551_/X sky130_fd_sc_hd__mux2_1
X_18749_ _19308_/CLK _18749_/D vssd1 vssd1 vccd1 vccd1 _18749_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12816__A1 _15700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10827__B1 _10606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09482_ _11202_/A vssd1 vssd1 vccd1 vccd1 _11014_/A sky130_fd_sc_hd__buf_2
XFILLER_51_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14229__S _14235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17507__A1 _17642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11252__B1 _10949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09843__S1 _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11307__A1 _10943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20007_ _20048_/CLK _20007_/D vssd1 vssd1 vccd1 vccd1 _20007_/Q sky130_fd_sc_hd__dfxtp_1
X_09818_ _09899_/A vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09749_ _09749_/A vssd1 vssd1 vccd1 vccd1 _09750_/A sky130_fd_sc_hd__buf_2
XFILLER_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10240__B _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13832__A _13832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17304__A _17304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12760_ _19813_/Q _17140_/C _12759_/X _19341_/Q vssd1 vssd1 vccd1 vccd1 _12760_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15757__A0 _19909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11928_/A _12673_/A _17581_/S vssd1 vssd1 vccd1 vccd1 _11764_/A sky130_fd_sc_hd__a21oi_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12691_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12692_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11352__A _11352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14430_ _14634_/A vssd1 vssd1 vccd1 vccd1 _14430_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11790_/A _11639_/X _11641_/X vssd1 vssd1 vccd1 vccd1 _11643_/A sky130_fd_sc_hd__o21a_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10046__A1 _10000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _18791_/Q _13731_/X _14363_/S vssd1 vssd1 vccd1 vccd1 _14362_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11573_ _12076_/A _12647_/A vssd1 vssd1 vccd1 vccd1 _11573_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput18 io_dbus_rdata[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_4
X_16100_ _13309_/X _19468_/Q _16106_/S vssd1 vssd1 vccd1 vccd1 _16101_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11794__A1 _19323_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ _19942_/Q _13312_/B vssd1 vssd1 vccd1 vccd1 _13335_/C sky130_fd_sc_hd__and2_1
Xinput29 io_dbus_rdata[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
X_10524_ _19468_/Q _19306_/Q _18715_/Q _18485_/Q _10559_/S _10510_/A vssd1 vssd1 vccd1
+ vccd1 _10524_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17080_ _17079_/A _17079_/C _19788_/Q vssd1 vssd1 vccd1 vccd1 _17081_/C sky130_fd_sc_hd__a21oi_1
X_14292_ _13847_/X _18761_/Q _14294_/S vssd1 vssd1 vccd1 vccd1 _14293_/A sky130_fd_sc_hd__mux2_1
X_16031_ _16031_/A vssd1 vssd1 vccd1 vccd1 _19437_/D sky130_fd_sc_hd__clkbuf_1
X_13243_ _19787_/Q vssd1 vssd1 vccd1 vccd1 _17079_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10455_ _10448_/Y _10450_/Y _10452_/Y _10454_/Y _09718_/A vssd1 vssd1 vccd1 vccd1
+ _10455_/X sky130_fd_sc_hd__o221a_1
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13174_ _13174_/A _13174_/B vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__or2_1
XFILLER_163_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10386_ _09820_/A _10378_/X _10380_/X _10385_/X _09605_/A vssd1 vssd1 vccd1 vccd1
+ _10386_/X sky130_fd_sc_hd__a311o_1
XANTENNA_output167_A _16453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ _12117_/Y _12121_/X _12124_/Y vssd1 vssd1 vccd1 vccd1 _12125_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17982_ _10456_/Y _17861_/X _17981_/X vssd1 vssd1 vccd1 vccd1 _19911_/D sky130_fd_sc_hd__a21oi_1
X_19721_ _19721_/CLK _19721_/D vssd1 vssd1 vccd1 vccd1 _19721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12056_ _12056_/A vssd1 vssd1 vccd1 vccd1 _12056_/Y sky130_fd_sc_hd__inv_2
X_16933_ _19740_/Q _16957_/C _16959_/B vssd1 vssd1 vccd1 vccd1 _16936_/B sky130_fd_sc_hd__and3_1
XFILLER_81_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11527__A _12606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _11001_/X _11005_/X _11006_/X _11014_/A _09472_/A vssd1 vssd1 vccd1 vccd1
+ _11012_/B sky130_fd_sc_hd__o221a_1
XFILLER_120_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19652_ _19789_/CLK _19652_/D vssd1 vssd1 vccd1 vccd1 _19652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16864_ _16864_/A _19715_/Q _16864_/C _16864_/D vssd1 vssd1 vccd1 vccd1 _16865_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18603_ _19485_/CLK _18603_/D vssd1 vssd1 vccd1 vccd1 _18603_/Q sky130_fd_sc_hd__dfxtp_1
X_15815_ _19919_/Q _12127_/A _15814_/Y vssd1 vssd1 vccd1 vccd1 _15815_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16795_ _19703_/Q _19702_/Q _16795_/C vssd1 vssd1 vccd1 vccd1 _16798_/B sky130_fd_sc_hd__and3_1
X_19583_ _19963_/CLK _19583_/D vssd1 vssd1 vccd1 vccd1 _19583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15433__S _15439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18534_ _19511_/CLK _18534_/D vssd1 vssd1 vccd1 vccd1 _18534_/Q sky130_fd_sc_hd__dfxtp_1
X_15746_ _19907_/Q _15708_/X _15745_/Y vssd1 vssd1 vccd1 vccd1 _15746_/X sky130_fd_sc_hd__a21o_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12958_ _18028_/A vssd1 vssd1 vccd1 vccd1 _17861_/A sky130_fd_sc_hd__buf_2
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10904__S0 _11493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11909_ _19583_/Q _11912_/B vssd1 vssd1 vccd1 vccd1 _12240_/B sky130_fd_sc_hd__and2_1
X_18465_ _19985_/CLK _18465_/D vssd1 vssd1 vccd1 vccd1 _18465_/Q sky130_fd_sc_hd__dfxtp_2
X_15677_ _15677_/A vssd1 vssd1 vccd1 vccd1 _19327_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _12889_/A vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__buf_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11262__A _18965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14628_ _14628_/A vssd1 vssd1 vccd1 vccd1 _14628_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17416_ _17486_/S vssd1 vssd1 vccd1 vccd1 _17500_/S sky130_fd_sc_hd__clkbuf_2
X_18396_ _18396_/A _18396_/B vssd1 vssd1 vccd1 vccd1 _20034_/D sky130_fd_sc_hd__nor2_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17347_ _17327_/A _12601_/Y _12824_/A _17358_/A _15818_/X vssd1 vssd1 vccd1 vccd1
+ _17348_/B sky130_fd_sc_hd__a32o_1
XFILLER_158_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14559_ _14559_/A vssd1 vssd1 vccd1 vccd1 _14568_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_147_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09667__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12982__B1 _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17278_ _15738_/X _19863_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17279_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19017_ _19500_/CLK _19017_/D vssd1 vssd1 vccd1 vccd1 _19017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16229_ _16369_/S vssd1 vssd1 vccd1 vccd1 _16252_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_173_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10606__A _10606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19919_ _19919_/CLK _19919_/D vssd1 vssd1 vccd1 vccd1 _19919_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10199__S1 _09822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__S0 _10702_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09603_ _09603_/A vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__buf_4
XFILLER_95_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16439__S _16441_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15343__S _15345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ _10678_/S vssd1 vssd1 vccd1 vccd1 _10509_/S sky130_fd_sc_hd__buf_6
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13462__B2 _19843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15739__A0 hold15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09465_ _11625_/B _12942_/S _17342_/B _09464_/X vssd1 vssd1 vccd1 vccd1 _09465_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09396_ _12689_/B _09397_/C vssd1 vssd1 vccd1 vccd1 _12810_/B sky130_fd_sc_hd__or2_4
XFILLER_149_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16174__S _16178_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18153__A1 _19968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__S0 _11003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09577__A _09577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11111__S _11305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10240_ _10240_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _10241_/B sky130_fd_sc_hd__nor2_1
XFILLER_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10171_ _19121_/Q _18887_/Q _19569_/Q _19217_/Q _09881_/X _10219_/A vssd1 vssd1 vccd1
+ vccd1 _10172_/B sky130_fd_sc_hd__mux4_2
XFILLER_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14422__S _14434_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13546__B _13546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13930_ _13998_/S vssd1 vssd1 vccd1 vccd1 _13939_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_120_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13861_ _13755_/X _18572_/Q _13867_/S vssd1 vssd1 vccd1 vccd1 _13862_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15600_ _14589_/X _19294_/Q _15600_/S vssd1 vssd1 vccd1 vccd1 _15601_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17034__A _17046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ _19645_/Q _13116_/A _12810_/Y _19677_/Q _12811_/X vssd1 vssd1 vccd1 vccd1
+ _12813_/B sky130_fd_sc_hd__a221o_1
XFILLER_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16580_ _16635_/A vssd1 vssd1 vccd1 vccd1 _16629_/A sky130_fd_sc_hd__buf_2
X_13792_ _13792_/A vssd1 vssd1 vccd1 vccd1 _18551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15531_ _19263_/Q _15215_/X _15539_/S vssd1 vssd1 vccd1 vccd1 _15532_/A sky130_fd_sc_hd__mux2_1
X_12743_ _12884_/A vssd1 vssd1 vccd1 vccd1 _16820_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18392__A1 _18302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18392__B2 _18391_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _18250_/A vssd1 vssd1 vccd1 vccd1 _19979_/D sky130_fd_sc_hd__clkbuf_1
X_15462_ _15462_/A vssd1 vssd1 vccd1 vccd1 _19232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12674_/A _12674_/B vssd1 vssd1 vccd1 vccd1 _12675_/A sky130_fd_sc_hd__and2_1
XFILLER_169_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _18289_/A vssd1 vssd1 vccd1 vccd1 _17201_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14413_/A vssd1 vssd1 vccd1 vccd1 _18807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11625_ _11625_/A _11625_/B _12942_/S vssd1 vssd1 vccd1 vccd1 _11625_/X sky130_fd_sc_hd__and3_1
X_18181_ _13428_/A _19981_/Q _18181_/S vssd1 vssd1 vccd1 vccd1 _18182_/A sky130_fd_sc_hd__mux2_1
X_15393_ _14602_/X _19202_/Q _15395_/S vssd1 vssd1 vccd1 vccd1 _15394_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18144__A1 _19964_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17132_ _17132_/A vssd1 vssd1 vccd1 vccd1 _19811_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12964__B1 _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09487__A _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14344_ _18783_/Q _13697_/X _14352_/S vssd1 vssd1 vccd1 vccd1 _14345_/A sky130_fd_sc_hd__mux2_1
X_11556_ _11556_/A _11558_/A _11556_/C vssd1 vssd1 vccd1 vccd1 _11556_/Y sky130_fd_sc_hd__nand3_1
XFILLER_129_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10507_ _09749_/A _10493_/X _10505_/X _09756_/A _10506_/Y vssd1 vssd1 vccd1 vccd1
+ _12654_/B sky130_fd_sc_hd__o32a_4
X_17063_ _17062_/A _17062_/C _19782_/Q vssd1 vssd1 vccd1 vccd1 _17064_/C sky130_fd_sc_hd__a21oi_1
X_14275_ _13822_/X _18753_/Q _14279_/S vssd1 vssd1 vccd1 vccd1 _14276_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11487_ _18793_/Q _19064_/Q _19288_/Q _19032_/Q _09532_/A _09514_/A vssd1 vssd1 vccd1
+ vccd1 _11487_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16014_ _16060_/S vssd1 vssd1 vccd1 vccd1 _16023_/S sky130_fd_sc_hd__buf_6
X_13226_ _19904_/Q _12851_/B _13520_/S vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ _10438_/A vssd1 vssd1 vccd1 vccd1 _10438_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15428__S _15428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _19858_/Q _13560_/A _13562_/A _19522_/Q vssd1 vssd1 vccd1 vccd1 _13157_/X
+ sky130_fd_sc_hd__a22o_1
X_10369_ _18814_/Q _19149_/Q _10465_/S vssd1 vssd1 vccd1 vccd1 _10369_/X sky130_fd_sc_hd__mux2_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12108_ _12108_/A _12145_/A vssd1 vssd1 vccd1 vccd1 _12111_/A sky130_fd_sc_hd__xor2_2
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ input27/X _12988_/X _13087_/X _13007_/X vssd1 vssd1 vccd1 vccd1 _15212_/A
+ sky130_fd_sc_hd__a22o_2
X_17965_ _18002_/A _17965_/B _17965_/C _17965_/D vssd1 vssd1 vccd1 vccd1 _17965_/X
+ sky130_fd_sc_hd__or4_1
X_19704_ _19721_/CLK _19704_/D vssd1 vssd1 vccd1 vccd1 _19704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16916_ _16919_/A _16916_/B _16930_/D vssd1 vssd1 vccd1 vccd1 _19736_/D sky130_fd_sc_hd__nor3_1
X_12039_ _18347_/A _12069_/A _12039_/C vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__and3_1
XANTENNA__10161__A _10161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17896_ _17914_/A vssd1 vssd1 vccd1 vccd1 _17985_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19635_ _19718_/CLK _19635_/D vssd1 vssd1 vccd1 vccd1 _19635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09991__S0 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16847_ _17073_/A vssd1 vssd1 vccd1 vccd1 _16946_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19566_ _19566_/CLK _19566_/D vssd1 vssd1 vccd1 vccd1 _19566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16778_ _19697_/Q _16781_/C _16777_/Y vssd1 vssd1 vccd1 vccd1 _19697_/D sky130_fd_sc_hd__o21a_1
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13444__B2 _19842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18517_ _19268_/CLK _18517_/D vssd1 vssd1 vccd1 vccd1 _18517_/Q sky130_fd_sc_hd__dfxtp_1
X_15729_ _15729_/A vssd1 vssd1 vccd1 vccd1 _19334_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11704__B _11704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19497_ _19497_/CLK _19497_/D vssd1 vssd1 vccd1 vccd1 _19497_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18383__B2 _18382_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09250_ _11675_/A _12595_/C _09263_/A _17378_/B _11724_/D vssd1 vssd1 vccd1 vccd1
+ _17393_/A sky130_fd_sc_hd__o32a_1
X_18448_ _19938_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _20026_/Q vssd1 vssd1 vccd1 vccd1 _09271_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14507__S _14513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_146_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18379_ _20029_/Q _18373_/X _18374_/X _18378_/Y vssd1 vssd1 vccd1 vccd1 _18380_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12955__B1 _10821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13647__A _14602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14242__S _14246_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15672__A2 _16303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14478__A _19323_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09517_ _10461_/A vssd1 vssd1 vccd1 vccd1 _10510_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11446__B1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ _17338_/B _18328_/A _09448_/C vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__or3_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09379_ _16809_/A _12797_/B vssd1 vssd1 vccd1 vccd1 _13136_/D sky130_fd_sc_hd__nor2_1
XANTENNA__12726__A _13527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18126__A1 _19924_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11410_ _11570_/A _11570_/B _11570_/C _11408_/Y _11409_/Y vssd1 vssd1 vccd1 vccd1
+ _11569_/B sky130_fd_sc_hd__a41o_4
XFILLER_137_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ _12390_/A _12390_/B vssd1 vssd1 vccd1 vccd1 _12391_/B sky130_fd_sc_hd__nand2_2
XFILLER_166_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11341_ _19452_/Q _19290_/Q _18699_/Q _18469_/Q _11161_/X _10974_/A vssd1 vssd1 vccd1
+ vccd1 _11342_/B sky130_fd_sc_hd__mux4_1
XFILLER_137_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14941__A _14987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18413__A _18413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14060_ _18660_/Q _13718_/X _14068_/S vssd1 vssd1 vccd1 vccd1 _14061_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11272_ _18636_/Q _19227_/Q _19389_/Q _18604_/Q _11262_/X _11113_/A vssd1 vssd1 vccd1
+ vccd1 _11272_/X sky130_fd_sc_hd__mux4_2
XFILLER_152_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13011_ _14074_/B vssd1 vssd1 vccd1 vccd1 _14917_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10223_ _18593_/Q _18854_/Q _18753_/Q _19088_/Q _09872_/X _09858_/X vssd1 vssd1 vccd1
+ vccd1 _10224_/B sky130_fd_sc_hd__mux4_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11921__A1 _12492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input43_A io_ibus_inst[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10280__S0 _10216_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _18658_/Q _19249_/Q _19411_/Q _18626_/Q _09508_/A _10148_/X vssd1 vssd1 vccd1
+ vccd1 _10154_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17971__B _17971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14962_ _14962_/A vssd1 vssd1 vccd1 vccd1 _19021_/D sky130_fd_sc_hd__clkbuf_1
X_17750_ _17616_/A _17746_/Y _17749_/Y vssd1 vssd1 vccd1 vccd1 _17750_/Y sky130_fd_sc_hd__a21oi_1
X_10085_ _10618_/A vssd1 vssd1 vccd1 vccd1 _10691_/A sky130_fd_sc_hd__clkbuf_4
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_102_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16701_ _19791_/Q _19790_/Q _19792_/Q _17082_/A vssd1 vssd1 vccd1 vccd1 _17090_/A
+ sky130_fd_sc_hd__and4_1
X_13913_ _13913_/A vssd1 vssd1 vccd1 vccd1 _13922_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__09973__S0 _10675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14893_ _14893_/A vssd1 vssd1 vccd1 vccd1 _18990_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17404__A3 _12620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17681_ _17681_/A vssd1 vssd1 vccd1 vccd1 _17681_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__14388__A _14592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19420_ _19727_/CLK _19420_/D vssd1 vssd1 vccd1 vccd1 _19420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13844_ _14669_/A vssd1 vssd1 vccd1 vccd1 _13844_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16632_ _19651_/Q _16629_/B _16631_/Y vssd1 vssd1 vccd1 vccd1 _19651_/D sky130_fd_sc_hd__o21a_1
XANTENNA__13426__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19351_ _19844_/CLK _19351_/D vssd1 vssd1 vccd1 vccd1 _19351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17699__A _18009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16563_ _19627_/Q _16564_/C _19628_/Q vssd1 vssd1 vccd1 vccd1 _16565_/B sky130_fd_sc_hd__a21oi_1
X_13775_ _13774_/X _18546_/Q _13781_/S vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__mux2_1
X_10987_ _19491_/Q _18903_/Q _18940_/Q _18514_/Q _11085_/A _09659_/A vssd1 vssd1 vccd1
+ vccd1 _10987_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18302_ _18302_/A _18302_/B vssd1 vssd1 vccd1 vccd1 _18302_/Y sky130_fd_sc_hd__nand2_1
X_15514_ _15514_/A vssd1 vssd1 vccd1 vccd1 _19256_/D sky130_fd_sc_hd__clkbuf_1
X_12726_ _13527_/B vssd1 vssd1 vccd1 vccd1 _13116_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11988__B2 _20049_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19282_ _19412_/CLK _19282_/D vssd1 vssd1 vccd1 vccd1 _19282_/Q sky130_fd_sc_hd__dfxtp_1
X_16494_ _19609_/Q _12628_/A _12625_/Y _12628_/Y _12749_/X vssd1 vssd1 vccd1 vccd1
+ _19609_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ _15918_/A _15445_/B vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__nor2_4
X_18233_ _18255_/A vssd1 vssd1 vccd1 vccd1 _18242_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_129_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12657_ _12657_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _12657_/Y sky130_fd_sc_hd__nor2_2
XFILLER_157_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12636__A _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18117__A1 _19923_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13231__S _13278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16108__A _16119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10099__S0 _11483_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11608_ _11608_/A vssd1 vssd1 vccd1 vccd1 _11619_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ _14574_/X _19194_/Q _15384_/S vssd1 vssd1 vccd1 vccd1 _15377_/A sky130_fd_sc_hd__mux2_1
X_18164_ _19941_/Q _19973_/Q _18170_/S vssd1 vssd1 vccd1 vccd1 _18165_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12588_ _17240_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _12588_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14327_ _14327_/A vssd1 vssd1 vccd1 vccd1 _18775_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17876__B1 _17875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17115_ _17115_/A vssd1 vssd1 vccd1 vccd1 _17120_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11539_ _11539_/A vssd1 vssd1 vccd1 vccd1 _11550_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18095_ _12538_/B _17755_/A _18094_/X _18028_/X vssd1 vssd1 vccd1 vccd1 _18095_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_144_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17046_ _17046_/A _17046_/B _17046_/C vssd1 vssd1 vccd1 vccd1 _19776_/D sky130_fd_sc_hd__nor3_1
XFILLER_172_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14258_ _14258_/A vssd1 vssd1 vccd1 vccd1 _18745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ _19620_/Q _13204_/X _13208_/X vssd1 vssd1 vccd1 vccd1 _13209_/X sky130_fd_sc_hd__o21a_1
XFILLER_143_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14062__S _14068_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14189_ _14189_/A vssd1 vssd1 vccd1 vccd1 _18714_/D sky130_fd_sc_hd__clkbuf_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18997_ _19317_/CLK _18997_/D vssd1 vssd1 vccd1 vccd1 _18997_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _17748_/S _17947_/X _17723_/X vssd1 vssd1 vccd1 vccd1 _17948_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_173_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19836_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_72_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14298__A _14354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17879_ _17884_/A _17884_/B vssd1 vssd1 vccd1 vccd1 _17883_/B sky130_fd_sc_hd__and2_1
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19618_ _19620_/CLK _19618_/D vssd1 vssd1 vccd1 vccd1 _19618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11715__A _11764_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_188_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19817_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19549_ _19551_/CLK _19549_/D vssd1 vssd1 vccd1 vccd1 _19549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11979__A1 _19521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09302_ _17394_/A _17381_/A _12664_/A vssd1 vssd1 vccd1 vccd1 _11615_/A sky130_fd_sc_hd__and3_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13930__A _13998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12640__A2 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09233_ _20052_/Q _11523_/A _09269_/B _11648_/C vssd1 vssd1 vccd1 vccd1 _11629_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA__12928__A0 _18311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19299_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10066__A _19919_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18233__A _18255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_126_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19394_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12156__A1 _17187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15068__S _15072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13377__A _13454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09997_ _09613_/A _09978_/X _09995_/X _09996_/X _19919_/Q vssd1 vssd1 vccd1 vccd1
+ _10139_/A sky130_fd_sc_hd__a32o_4
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14700__S _14702_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10910_ _10910_/A _10910_/B vssd1 vssd1 vccd1 vccd1 _10910_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11890_ _12214_/A vssd1 vssd1 vccd1 vccd1 _11890_/X sky130_fd_sc_hd__buf_2
XFILLER_72_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13408__A1 _13407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ _18644_/Q _19235_/Q _19397_/Q _18612_/Q _11429_/S _09985_/X vssd1 vssd1 vccd1
+ vccd1 _10841_/X sky130_fd_sc_hd__mux4_2
XFILLER_60_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15531__S _15539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13560_ _13560_/A _13560_/B _17247_/D vssd1 vssd1 vccd1 vccd1 _13562_/B sky130_fd_sc_hd__nor3_1
XFILLER_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10772_ _19904_/Q vssd1 vssd1 vccd1 vccd1 _10772_/Y sky130_fd_sc_hd__inv_2
X_12511_ _19604_/Q _19605_/Q _12511_/C vssd1 vssd1 vccd1 vccd1 _12540_/B sky130_fd_sc_hd__and3_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ _19952_/Q _19953_/Q _13491_/C vssd1 vssd1 vccd1 vccd1 _13512_/B sky130_fd_sc_hd__and3_1
XFILLER_157_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15230_ _15230_/A vssd1 vssd1 vccd1 vccd1 _19139_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12442_ _19538_/Q _11782_/X _13591_/A vssd1 vssd1 vccd1 vccd1 _12442_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12073__A1_N _12376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13986__S _13994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15161_ _19112_/Q vssd1 vssd1 vccd1 vccd1 _15162_/A sky130_fd_sc_hd__clkbuf_1
X_12373_ _19838_/Q _17210_/A _12373_/C vssd1 vssd1 vccd1 vccd1 _12419_/C sky130_fd_sc_hd__and3_1
XFILLER_138_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14112_ _18682_/Q _13676_/X _14120_/S vssd1 vssd1 vccd1 vccd1 _14113_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11324_ _11313_/X _11323_/X _09341_/X _09618_/A vssd1 vssd1 vccd1 vccd1 _11324_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15092_ _14618_/X _19079_/Q _15094_/S vssd1 vssd1 vccd1 vccd1 _15093_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18920_ _19377_/CLK _18920_/D vssd1 vssd1 vccd1 vccd1 _18920_/Q sky130_fd_sc_hd__dfxtp_1
X_14043_ _14043_/A vssd1 vssd1 vccd1 vccd1 _18652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11255_ _12633_/B _11348_/A _12634_/B _11254_/Y vssd1 vssd1 vccd1 vccd1 _11581_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_153_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10704__A _11046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ _19378_/Q _18992_/Q _19442_/Q _18561_/Q _10160_/S _10196_/A vssd1 vssd1 vccd1
+ vccd1 _10207_/B sky130_fd_sc_hd__mux4_1
X_18851_ _19565_/CLK _18851_/D vssd1 vssd1 vccd1 vccd1 _18851_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10253__S0 _09902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_90_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19369_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11186_ _11178_/Y _11181_/Y _11183_/Y _11185_/Y _10994_/A vssd1 vssd1 vccd1 vccd1
+ _11186_/X sky130_fd_sc_hd__o221a_2
XANTENNA__16598__A _16631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17802_ _17565_/S _17802_/B _17802_/C _17802_/D vssd1 vssd1 vccd1 vccd1 _17802_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10137_ _10137_/A _12666_/B vssd1 vssd1 vccd1 vccd1 _11544_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18782_ _19407_/CLK _18782_/D vssd1 vssd1 vccd1 vccd1 _18782_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14610__S _14622_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15994_ _15994_/A vssd1 vssd1 vccd1 vccd1 _19420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17733_ _17560_/X _17717_/X _17732_/X _17598_/X vssd1 vssd1 vccd1 vccd1 _17733_/X
+ sky130_fd_sc_hd__o211a_1
X_14945_ _14945_/A vssd1 vssd1 vccd1 vccd1 _19013_/D sky130_fd_sc_hd__clkbuf_1
X_10068_ _10139_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _11543_/A sky130_fd_sc_hd__and2_1
XFILLER_85_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09720__C1 _09719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17664_ _17664_/A vssd1 vssd1 vccd1 vccd1 _17664_/Y sky130_fd_sc_hd__inv_2
X_14876_ _14618_/X _18983_/Q _14878_/S vssd1 vssd1 vccd1 vccd1 _14877_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19403_ _19405_/CLK _19403_/D vssd1 vssd1 vccd1 vccd1 _19403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16615_ _16617_/B _16617_/C _16577_/X vssd1 vssd1 vccd1 vccd1 _16615_/Y sky130_fd_sc_hd__a21oi_1
X_13827_ _13827_/A vssd1 vssd1 vccd1 vccd1 _18562_/D sky130_fd_sc_hd__clkbuf_1
X_17595_ _17578_/X _17593_/X _17805_/S vssd1 vssd1 vccd1 vccd1 _17595_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14846__A _14902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13750__A _18299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15441__S _15443_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19334_ _19783_/CLK _19334_/D vssd1 vssd1 vccd1 vccd1 _19334_/Q sky130_fd_sc_hd__dfxtp_1
X_16546_ _16547_/B _16547_/C _19622_/Q vssd1 vssd1 vccd1 vccd1 _16548_/B sky130_fd_sc_hd__a21oi_1
X_13758_ _14583_/A vssd1 vssd1 vccd1 vccd1 _13758_/X sky130_fd_sc_hd__buf_2
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ _19866_/Q _12755_/A _12704_/X _19530_/Q _12708_/X vssd1 vssd1 vccd1 vccd1
+ _12709_/X sky130_fd_sc_hd__a221o_1
XFILLER_148_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19265_ _19491_/CLK _19265_/D vssd1 vssd1 vccd1 vccd1 _19265_/Q sky130_fd_sc_hd__dfxtp_1
X_13689_ _14634_/A vssd1 vssd1 vccd1 vccd1 _13689_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16477_ _16487_/A vssd1 vssd1 vccd1 vccd1 _16477_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18216_ _19964_/Q _19585_/Q _18220_/S vssd1 vssd1 vccd1 vccd1 _18217_/A sky130_fd_sc_hd__mux2_1
X_15428_ _14653_/X _19218_/Q _15428_/S vssd1 vssd1 vccd1 vccd1 _15429_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_19_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19196_ _19196_/CLK _19196_/D vssd1 vssd1 vccd1 vccd1 _19196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_43_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19570_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13896__S _13900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15359_ _19187_/Q _15279_/X _15367_/S vssd1 vssd1 vccd1 vccd1 _15360_/A sky130_fd_sc_hd__mux2_1
X_18147_ _18147_/A vssd1 vssd1 vccd1 vccd1 _19933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18078_ _18076_/Y _18077_/X _18078_/S vssd1 vssd1 vccd1 vccd1 _18078_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09920_ _09479_/A _09913_/X _09915_/X _09919_/X _09605_/A vssd1 vssd1 vccd1 vccd1
+ _09920_/X sky130_fd_sc_hd__a311o_1
XFILLER_116_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17029_ _19765_/Q _17026_/C _17028_/Y vssd1 vssd1 vccd1 vccd1 _19765_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10614__A _10824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_58_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19129_/CLK sky130_fd_sc_hd__clkbuf_16
X_20040_ _20052_/CLK _20040_/D vssd1 vssd1 vccd1 vccd1 _20040_/Q sky130_fd_sc_hd__dfxtp_1
X_09851_ _10392_/S vssd1 vssd1 vccd1 vccd1 _09924_/S sky130_fd_sc_hd__buf_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15616__S _15622_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10795__S1 _11496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _10184_/A vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14520__S _14524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09937__S0 _10173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _18931_/Q vssd1 vssd1 vccd1 vccd1 _13163_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17786__B _17792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10508__B _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14491__A _17123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09585__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11040_ _09999_/A _11025_/Y _11033_/X _11039_/Y _09737_/A vssd1 vssd1 vccd1 vccd1
+ _11040_/X sky130_fd_sc_hd__o311a_1
XFILLER_118_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10786__S1 _10037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18416__A1_N _18336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12991_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11355__A _11355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14730_ _14730_/A vssd1 vssd1 vccd1 vccd1 _18917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11942_ _11870_/C _11819_/X _11940_/A vssd1 vssd1 vccd1 vccd1 _11942_/X sky130_fd_sc_hd__a21o_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14660_/X _18890_/Q _14670_/S vssd1 vssd1 vccd1 vccd1 _14662_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _12444_/A vssd1 vssd1 vccd1 vccd1 _15719_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15261__S _15261_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18138__A _18138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16400_ _13239_/X _19558_/Q _16404_/S vssd1 vssd1 vccd1 vccd1 _16401_/A sky130_fd_sc_hd__mux2_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _15061_/A _18297_/A _15373_/A _14917_/D vssd1 vssd1 vccd1 vccd1 _13719_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _18676_/Q _19171_/Q _10824_/S vssd1 vssd1 vccd1 vccd1 _10825_/B sky130_fd_sc_hd__mux2_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _12610_/A _09269_/D _11648_/C _11619_/A _17331_/X vssd1 vssd1 vccd1 vccd1
+ _17382_/B sky130_fd_sc_hd__o311a_1
X_14592_ _14592_/A vssd1 vssd1 vccd1 vccd1 _14592_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16331_ _16331_/A vssd1 vssd1 vccd1 vccd1 _19537_/D sky130_fd_sc_hd__clkbuf_1
X_13543_ _19956_/Q _13543_/B vssd1 vssd1 vccd1 vccd1 _13543_/Y sky130_fd_sc_hd__xnor2_1
X_10755_ _10703_/A _10752_/Y _10754_/Y _10846_/A vssd1 vssd1 vccd1 vccd1 _10755_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10710__S1 _10014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19050_ _19500_/CLK _19050_/D vssd1 vssd1 vccd1 vccd1 _19050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16262_ _12854_/X _16261_/Y _16262_/S vssd1 vssd1 vccd1 vccd1 _16262_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_20_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13474_ input20/X _13303_/X _13436_/X vssd1 vssd1 vccd1 vccd1 _13474_/Y sky130_fd_sc_hd__a21oi_1
X_10686_ _11440_/A _10683_/X _10685_/X _10621_/X vssd1 vssd1 vccd1 vccd1 _10686_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18001_ _18001_/A _18001_/B vssd1 vssd1 vccd1 vccd1 _18002_/D sky130_fd_sc_hd__nor2_1
X_15213_ _19134_/Q _15212_/X _15213_/S vssd1 vssd1 vccd1 vccd1 _15214_/A sky130_fd_sc_hd__mux2_1
X_12425_ _18333_/A _12475_/B vssd1 vssd1 vccd1 vccd1 _12425_/X sky130_fd_sc_hd__or2_2
X_16193_ _16193_/A vssd1 vssd1 vccd1 vccd1 _19509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09495__A _18965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15144_ _15144_/A vssd1 vssd1 vccd1 vccd1 _19103_/D sky130_fd_sc_hd__clkbuf_1
X_12356_ _12356_/A vssd1 vssd1 vccd1 vccd1 _18012_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_153_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12633__B _12633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ _10943_/X _11306_/X _11271_/A vssd1 vssd1 vccd1 vccd1 _11307_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15075_ _14592_/X _19071_/Q _15083_/S vssd1 vssd1 vccd1 vccd1 _15076_/A sky130_fd_sc_hd__mux2_1
X_19952_ _19952_/CLK hold7/X vssd1 vssd1 vccd1 vccd1 _19952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12287_ _12395_/S _12287_/B vssd1 vssd1 vccd1 vccd1 _12287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14026_ _14072_/S vssd1 vssd1 vccd1 vccd1 _14035_/S sky130_fd_sc_hd__buf_2
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18903_ _19042_/CLK _18903_/D vssd1 vssd1 vccd1 vccd1 _18903_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output74_A _12117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ _11001_/A _11237_/X _10941_/X vssd1 vssd1 vccd1 vccd1 _11238_/X sky130_fd_sc_hd__a21o_1
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19883_ _20052_/CLK _19883_/D vssd1 vssd1 vccd1 vccd1 _19883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18834_ _19389_/CLK _18834_/D vssd1 vssd1 vccd1 vccd1 _18834_/Q sky130_fd_sc_hd__dfxtp_1
X_11169_ _11164_/X _11166_/Y _11168_/Y _11295_/A vssd1 vssd1 vccd1 vccd1 _11169_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18765_ _19484_/CLK _18765_/D vssd1 vssd1 vccd1 vccd1 _18765_/Q sky130_fd_sc_hd__dfxtp_1
X_15977_ _15977_/A vssd1 vssd1 vccd1 vccd1 _19413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17716_ _17715_/X _17693_/X _17887_/S vssd1 vssd1 vccd1 vccd1 _17716_/X sky130_fd_sc_hd__mux2_1
X_14928_ _19006_/Q _14385_/X _14928_/S vssd1 vssd1 vccd1 vccd1 _14929_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18696_ _19417_/CLK _18696_/D vssd1 vssd1 vccd1 vccd1 _18696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17647_ _17461_/X _17417_/X _17660_/S vssd1 vssd1 vccd1 vccd1 _17647_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14859_ _14592_/X _18975_/Q _14867_/S vssd1 vssd1 vccd1 vccd1 _14860_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14576__A _14657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17578_ _17567_/X _17576_/X _17810_/S vssd1 vssd1 vccd1 vccd1 _17578_/X sky130_fd_sc_hd__mux2_1
X_19317_ _19317_/CLK _19317_/D vssd1 vssd1 vccd1 vccd1 _19317_/Q sky130_fd_sc_hd__dfxtp_1
X_16529_ _19617_/Q _19616_/Q _19615_/Q _16529_/D vssd1 vssd1 vccd1 vccd1 _16540_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__12096__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10609__A _10609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19248_ _19411_/CLK _19248_/D vssd1 vssd1 vccd1 vccd1 _19248_/Q sky130_fd_sc_hd__dfxtp_1
X_19179_ _19406_/CLK _19179_/D vssd1 vssd1 vccd1 vccd1 _19179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15200__A _15299_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ _10368_/A _09903_/B vssd1 vssd1 vccd1 vccd1 _09903_/X sky130_fd_sc_hd__and2_1
XFILLER_99_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09834_ _10509_/S vssd1 vssd1 vccd1 vccd1 _10559_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_113_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20023_ _20027_/CLK _20023_/D vssd1 vssd1 vccd1 vccd1 _20023_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17127__A _17127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _19126_/Q _18892_/Q _19574_/Q _19222_/Q _09763_/S _09526_/A vssd1 vssd1 vccd1
+ vccd1 _09765_/X sky130_fd_sc_hd__mux4_2
XFILLER_74_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15870__A _15916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09696_ _09696_/A vssd1 vssd1 vccd1 vccd1 _09696_/X sky130_fd_sc_hd__buf_2
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11193__S1 _11260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14486__A _14831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12047__A0 _19967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15784__B2 _18458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10519__A _10519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11114__S _11114_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ _10583_/A _10539_/X _10322_/A vssd1 vssd1 vccd1 vccd1 _10540_/X sky130_fd_sc_hd__o21a_1
XFILLER_22_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ _18588_/Q _18849_/Q _18748_/Q _19083_/Q _10470_/X _10462_/A vssd1 vssd1 vccd1
+ vccd1 _10472_/B sky130_fd_sc_hd__mux4_1
XFILLER_155_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14425__S _14434_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12734__A _15700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16206__A _16206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12210_ _12286_/A vssd1 vssd1 vccd1 vccd1 _12583_/S sky130_fd_sc_hd__buf_2
XFILLER_157_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13190_ _19934_/Q vssd1 vssd1 vccd1 vccd1 _13191_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12141_ _19970_/Q _11406_/A _12198_/S vssd1 vssd1 vccd1 vccd1 _17451_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18421__A input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10208__S0 _10160_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12072_ _12320_/A _17394_/B _12071_/X vssd1 vssd1 vccd1 vccd1 _12072_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15900_ _15900_/A vssd1 vssd1 vccd1 vccd1 _19379_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10759__S1 _10718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ _09611_/A _11012_/X _11022_/X _09619_/A _19899_/Q vssd1 vssd1 vccd1 vccd1
+ _11352_/A sky130_fd_sc_hd__a32o_4
XFILLER_104_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16880_ _19724_/Q _19723_/Q _19722_/Q _16880_/D vssd1 vssd1 vccd1 vccd1 _16888_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15831_ _15831_/A vssd1 vssd1 vccd1 vccd1 _19352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11085__A _11085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11089__A1 _10899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18550_ _19431_/CLK _18550_/D vssd1 vssd1 vccd1 vccd1 _18550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _18460_/Q _12973_/X _11421_/A _12969_/X vssd1 vssd1 vccd1 vccd1 _18460_/D
+ sky130_fd_sc_hd__a22o_1
X_15762_ _15761_/X _19341_/Q _15772_/S vssd1 vssd1 vccd1 vccd1 _15763_/A sky130_fd_sc_hd__mux2_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17501_ _17601_/S vssd1 vssd1 vccd1 vccd1 _17686_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11184__S1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _18910_/Q _14417_/X _14713_/S vssd1 vssd1 vccd1 vccd1 _14714_/A sky130_fd_sc_hd__mux2_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18481_ _19464_/CLK _18481_/D vssd1 vssd1 vccd1 vccd1 _18481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11925_ _11961_/A _12638_/B _11962_/A _12475_/A vssd1 vssd1 vccd1 vccd1 _11926_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16087__S _16095_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output112_A _12648_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15693_ _18443_/Q _15693_/B _15693_/C vssd1 vssd1 vccd1 vccd1 _15693_/X sky130_fd_sc_hd__or3_1
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _17702_/B _12529_/A _17450_/S vssd1 vssd1 vccd1 vccd1 _17432_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14644_ _14644_/A vssd1 vssd1 vccd1 vccd1 _14644_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__15775__A1 _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11856_ _11899_/B _11855_/X _11856_/S vssd1 vssd1 vccd1 vccd1 _17594_/A sky130_fd_sc_hd__mux2_2
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12589__A1 _12421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ _10746_/A _10806_/X _09976_/A vssd1 vssd1 vccd1 vccd1 _10807_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14575_ _16371_/A _15373_/C _16371_/C _15589_/B vssd1 vssd1 vccd1 vccd1 _14657_/A
+ sky130_fd_sc_hd__or4_4
X_17363_ _09202_/Y _18301_/A _17358_/X _19888_/Q vssd1 vssd1 vccd1 vccd1 _17364_/B
+ sky130_fd_sc_hd__a22o_1
X_11787_ _11787_/A vssd1 vssd1 vccd1 vccd1 _12606_/D sky130_fd_sc_hd__clkbuf_2
X_19102_ _19794_/CLK _19102_/D vssd1 vssd1 vccd1 vccd1 _19102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16314_ _16317_/B _16313_/X _12127_/X vssd1 vssd1 vccd1 vccd1 _16314_/X sky130_fd_sc_hd__o21a_1
X_10738_ _10734_/X _10736_/X _10737_/X _11438_/A _09979_/X vssd1 vssd1 vccd1 vccd1
+ _10738_/X sky130_fd_sc_hd__o221a_1
X_13526_ input24/X _13353_/X _13354_/X vssd1 vssd1 vccd1 vccd1 _13539_/A sky130_fd_sc_hd__a21oi_1
X_17294_ _17209_/Y _19870_/Q _17302_/S vssd1 vssd1 vccd1 vccd1 _17295_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19033_ _19129_/CLK _19033_/D vssd1 vssd1 vccd1 vccd1 _19033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16245_ _16213_/X _16244_/Y _15712_/Y vssd1 vssd1 vccd1 vccd1 _16245_/X sky130_fd_sc_hd__a21o_1
X_13457_ input19/X _13318_/X _13436_/X vssd1 vssd1 vccd1 vccd1 _13457_/X sky130_fd_sc_hd__a21o_1
X_10669_ _19907_/Q vssd1 vssd1 vccd1 vccd1 _10669_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14335__S _14341_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12644__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ _12410_/A _18036_/B vssd1 vssd1 vccd1 vccd1 _12521_/A sky130_fd_sc_hd__or2_2
XANTENNA__10447__S0 _10337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16176_ _19502_/Q _14634_/A _16178_/S vssd1 vssd1 vccd1 vccd1 _16177_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13388_ _19663_/Q _12887_/X _12889_/X _19795_/Q _13387_/X vssd1 vssd1 vccd1 vccd1
+ _15782_/B sky130_fd_sc_hd__a221o_4
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput106 _17379_/A vssd1 vssd1 vccd1 vccd1 io_dbus_rd_en sky130_fd_sc_hd__buf_2
XFILLER_126_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput117 _12654_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[17] sky130_fd_sc_hd__buf_2
X_15127_ _14669_/X _19095_/Q _15127_/S vssd1 vssd1 vccd1 vccd1 _15128_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput128 _12666_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[27] sky130_fd_sc_hd__buf_2
XANTENNA__12761__B2 _19531_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12339_ _19595_/Q _12339_/B _12339_/C _12339_/D vssd1 vssd1 vccd1 vccd1 _12340_/B
+ sky130_fd_sc_hd__and4_1
Xoutput139 _12643_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[8] sky130_fd_sc_hd__buf_2
XFILLER_5_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18229__A0 _19970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09953__A _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19935_ _19938_/CLK _19935_/D vssd1 vssd1 vccd1 vccd1 _19935_/Q sky130_fd_sc_hd__dfxtp_1
X_15058_ _15058_/A vssd1 vssd1 vccd1 vccd1 _19064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _18637_/Q _13622_/X _14013_/S vssd1 vssd1 vccd1 vccd1 _14010_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14070__S _14072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19866_ _19881_/CLK _19866_/D vssd1 vssd1 vccd1 vccd1 _19866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18817_ _19058_/CLK _18817_/D vssd1 vssd1 vccd1 vccd1 _18817_/Q sky130_fd_sc_hd__dfxtp_1
X_19797_ _19803_/CLK _19797_/D vssd1 vssd1 vccd1 vccd1 _19797_/Q sky130_fd_sc_hd__dfxtp_1
X_09550_ _10368_/A vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__buf_2
XFILLER_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18748_ _19308_/CLK _18748_/D vssd1 vssd1 vccd1 vccd1 _18748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17204__A1 _12772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10827__A1 _09985_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ _11274_/A vssd1 vssd1 vccd1 vccd1 _11202_/A sky130_fd_sc_hd__clkbuf_2
X_18679_ _19272_/CLK _18679_/D vssd1 vssd1 vccd1 vccd1 _18679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11723__A _18340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12538__B _12538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13529__B1 _12805_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10074__A _10074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20006_ _20020_/CLK _20006_/D vssd1 vssd1 vccd1 vccd1 _20006_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10610__S0 _10608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ _09817_/A vssd1 vssd1 vccd1 vccd1 _09899_/A sky130_fd_sc_hd__buf_4
XFILLER_47_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17994__A2 _17861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _09748_/A vssd1 vssd1 vccd1 vccd1 _09749_/A sky130_fd_sc_hd__buf_4
XANTENNA__12807__A2 _13546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _10039_/A vssd1 vssd1 vccd1 vccd1 _09680_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11710_ _11898_/D vssd1 vssd1 vccd1 vccd1 _17581_/S sky130_fd_sc_hd__buf_2
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12804_/A _12837_/B vssd1 vssd1 vccd1 vccd1 _12991_/A sky130_fd_sc_hd__nor2_2
XANTENNA__15757__A1 _12741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11641_ _18288_/A _11663_/C _11641_/C _11641_/D vssd1 vssd1 vccd1 vccd1 _11641_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__11352__B _12638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14360_ _14360_/A vssd1 vssd1 vccd1 vccd1 _18790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11572_ _11570_/B _11570_/C _11570_/A vssd1 vssd1 vccd1 vccd1 _11572_/X sky130_fd_sc_hd__a21o_1
XFILLER_156_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _13311_/A vssd1 vssd1 vccd1 vccd1 _18485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10523_ _10523_/A _10523_/B vssd1 vssd1 vccd1 vccd1 _10523_/X sky130_fd_sc_hd__or2_1
Xinput19 io_dbus_rdata[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_6
XFILLER_11_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11794__A2 _11665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14291_ _14291_/A vssd1 vssd1 vccd1 vccd1 _18760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14155__S _14163_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16030_ _13321_/X _19437_/Q _16034_/S vssd1 vssd1 vccd1 vccd1 _16031_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10429__S0 _10465_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13242_ _19655_/Q vssd1 vssd1 vccd1 vccd1 _16645_/A sky130_fd_sc_hd__clkbuf_2
X_10454_ _10436_/A _10453_/X _10323_/X vssd1 vssd1 vccd1 vccd1 _10454_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_136_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13994__S _13994_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13173_ _13173_/A _13173_/B _19888_/Q input30/X vssd1 vssd1 vccd1 vccd1 _13174_/B
+ sky130_fd_sc_hd__and4_1
X_10385_ _10378_/A _10381_/X _10384_/X _09826_/A vssd1 vssd1 vccd1 vccd1 _10385_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ _19526_/Q _12122_/X _12123_/X vssd1 vssd1 vccd1 vccd1 _12124_/Y sky130_fd_sc_hd__o21ai_1
X_17981_ _12287_/B _17844_/X _17980_/X _17858_/X vssd1 vssd1 vccd1 vccd1 _17981_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19720_ _19720_/CLK _19720_/D vssd1 vssd1 vccd1 vccd1 _19720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16932_ _16957_/C _16959_/B _16931_/Y vssd1 vssd1 vccd1 vccd1 _19739_/D sky130_fd_sc_hd__o21a_1
X_12055_ _12055_/A _12055_/B vssd1 vssd1 vccd1 vccd1 _12056_/A sky130_fd_sc_hd__xnor2_4
XFILLER_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11006_ _19104_/Q _18870_/Q _19552_/Q _19200_/Q _09530_/A _11236_/A vssd1 vssd1 vccd1
+ vccd1 _11006_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17434__A1 _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19651_ _19789_/CLK _19651_/D vssd1 vssd1 vccd1 vccd1 _19651_/Q sky130_fd_sc_hd__dfxtp_1
X_16863_ _19713_/Q _19712_/Q _16863_/C _16863_/D vssd1 vssd1 vccd1 vccd1 _16864_/D
+ sky130_fd_sc_hd__and4_1
X_18602_ _19480_/CLK _18602_/D vssd1 vssd1 vccd1 vccd1 _18602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15814_ _15814_/A _17228_/A vssd1 vssd1 vccd1 vccd1 _15814_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19582_ _19592_/CLK _19582_/D vssd1 vssd1 vccd1 vccd1 _19582_/Q sky130_fd_sc_hd__dfxtp_1
X_16794_ _19702_/Q _16795_/C _16793_/Y vssd1 vssd1 vccd1 vccd1 _19702_/D sky130_fd_sc_hd__o21a_1
XFILLER_133_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18533_ _19510_/CLK _18533_/D vssd1 vssd1 vccd1 vccd1 _18533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _15814_/A _17191_/A vssd1 vssd1 vccd1 vccd1 _15745_/Y sky130_fd_sc_hd__nor2_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _18449_/Q _12951_/X _10727_/A _12954_/X vssd1 vssd1 vccd1 vccd1 _18449_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18464_ _19985_/CLK _18464_/D vssd1 vssd1 vccd1 vccd1 _18464_/Q sky130_fd_sc_hd__dfxtp_2
X_11908_ _19583_/Q _12218_/A vssd1 vssd1 vccd1 vccd1 _11923_/A sky130_fd_sc_hd__or2_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ _15675_/X _19327_/Q _15684_/S vssd1 vssd1 vccd1 vccd1 _15677_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12888_ _12888_/A vssd1 vssd1 vccd1 vccd1 _12889_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13759__A0 _13758_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17415_ _17586_/S vssd1 vssd1 vccd1 vccd1 _17486_/S sky130_fd_sc_hd__clkbuf_2
X_14627_ _14627_/A vssd1 vssd1 vccd1 vccd1 _18879_/D sky130_fd_sc_hd__clkbuf_1
X_18395_ _18306_/A _12880_/A _14481_/X _18394_/Y vssd1 vssd1 vccd1 vccd1 _18396_/B
+ sky130_fd_sc_hd__o22a_1
X_11839_ _12693_/A _12914_/A _11839_/C _11952_/C vssd1 vssd1 vccd1 vccd1 _11839_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_60_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17230__A _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17346_ _17346_/A _17346_/B vssd1 vssd1 vccd1 vccd1 _17358_/A sky130_fd_sc_hd__and2_1
X_14558_ _14558_/A vssd1 vssd1 vccd1 vccd1 _18856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12982__A1 _18466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13509_ input22/X _13353_/A _13436_/X vssd1 vssd1 vccd1 vccd1 _13509_/X sky130_fd_sc_hd__a21o_1
XFILLER_146_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17277_ _17277_/A vssd1 vssd1 vccd1 vccd1 _19862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14489_ _17041_/B _18409_/B vssd1 vssd1 vccd1 vccd1 _18828_/D sky130_fd_sc_hd__nor2_4
XANTENNA__10993__B1 _10920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19016_ _19495_/CLK _19016_/D vssd1 vssd1 vccd1 vccd1 _19016_/Q sky130_fd_sc_hd__dfxtp_1
X_16228_ _16299_/A vssd1 vssd1 vccd1 vccd1 _16369_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__17884__B _17884_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16159_ _19494_/Q _14608_/A _16167_/S vssd1 vssd1 vccd1 vccd1 _16160_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16476__A2 _16449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15684__A0 _15683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12498__B1 _12429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19918_ _19919_/CLK _19918_/D vssd1 vssd1 vccd1 vccd1 _19918_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11396__S1 _09662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_142_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19849_ _19857_/CLK _19849_/D vssd1 vssd1 vccd1 vccd1 _19849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09602_ _09602_/A vssd1 vssd1 vccd1 vccd1 _09603_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09533_ _10811_/S vssd1 vssd1 vccd1 vccd1 _10678_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_58_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13462__A2 _12992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15739__A1 _15738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _18028_/A vssd1 vssd1 vccd1 vccd1 _09464_/X sky130_fd_sc_hd__buf_4
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16963__B _19744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09395_ _20015_/Q _12688_/A _12688_/B _09389_/A vssd1 vssd1 vccd1 vccd1 _09397_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12422__B1 _12421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10433__C1 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__S1 _11059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12284__A _12287_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_67_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10736__B1 _10746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10170_ _09616_/X _10158_/X _10169_/X _09623_/X _19916_/Q vssd1 vssd1 vccd1 vccd1
+ _11421_/A sky130_fd_sc_hd__a32o_2
XANTENNA__10831__S0 _09532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15675__B1 _13597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14004__A _14072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _13860_/A vssd1 vssd1 vccd1 vccd1 _18571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12811_ _19777_/Q _12888_/A _13341_/A _19709_/Q vssd1 vssd1 vccd1 vccd1 _12811_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10678__S _10678_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13791_ _13790_/X _18551_/Q _13797_/S vssd1 vssd1 vccd1 vccd1 _13792_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _15587_/S vssd1 vssd1 vccd1 vccd1 _15539_/S sky130_fd_sc_hd__buf_2
XFILLER_103_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12742_ input70/X vssd1 vssd1 vccd1 vccd1 _12884_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12673_/A _12673_/B vssd1 vssd1 vccd1 vccd1 _12674_/B sky130_fd_sc_hd__or2_1
X_15461_ _19232_/Q _15219_/X _15467_/S vssd1 vssd1 vccd1 vccd1 _15462_/A sky130_fd_sc_hd__mux2_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17200_ _17319_/A vssd1 vssd1 vccd1 vccd1 _18289_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_169_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14412_ _18807_/Q _14411_/X _14418_/S vssd1 vssd1 vccd1 vccd1 _14413_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11624_/A _17336_/A _11624_/C vssd1 vssd1 vccd1 vccd1 _11625_/A sky130_fd_sc_hd__nor3_1
X_18180_ _18180_/A vssd1 vssd1 vccd1 vccd1 _19948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15392_ _15392_/A vssd1 vssd1 vccd1 vccd1 _19201_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10424__C1 _10519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17131_ _19811_/Q _17141_/A _17245_/S vssd1 vssd1 vccd1 vccd1 _17132_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12964__A1 _18453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14343_ _14354_/A vssd1 vssd1 vccd1 vccd1 _14352_/S sky130_fd_sc_hd__buf_2
X_11555_ _11558_/A _11556_/C _11556_/A vssd1 vssd1 vccd1 vccd1 _11555_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10506_ _19910_/Q vssd1 vssd1 vccd1 vccd1 _10506_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_7_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14274_ _14274_/A vssd1 vssd1 vccd1 vccd1 _18752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17062_ _17062_/A _19782_/Q _17062_/C vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__and3_1
XFILLER_144_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ _11482_/X _11484_/X _11485_/X _11473_/A _09473_/A vssd1 vssd1 vccd1 vccd1
+ _11491_/B sky130_fd_sc_hd__o221a_1
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13225_ _19936_/Q _13225_/B vssd1 vssd1 vccd1 vccd1 _13254_/C sky130_fd_sc_hd__and2_1
X_16013_ _16013_/A vssd1 vssd1 vccd1 vccd1 _19429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10437_ _18685_/Q _19180_/Q _10496_/S vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14613__S _14622_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09593__B1 _09479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12192__A2 _12651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ _19332_/Q _13154_/Y _13155_/Y vssd1 vssd1 vccd1 vccd1 _13156_/X sky130_fd_sc_hd__o21a_1
X_10368_ _10368_/A _10368_/B vssd1 vssd1 vccd1 vccd1 _10368_/X sky130_fd_sc_hd__and2_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15666__A0 _15661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _19969_/Q _10727_/A _12198_/S vssd1 vssd1 vccd1 vccd1 _12145_/A sky130_fd_sc_hd__mux2_2
XFILLER_2_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13073_/X _13085_/X _13147_/S vssd1 vssd1 vccd1 vccd1 _13087_/X sky130_fd_sc_hd__mux2_1
X_17964_ _17960_/B _17964_/B vssd1 vssd1 vccd1 vccd1 _17965_/D sky130_fd_sc_hd__and2b_1
X_10299_ _10428_/A _10292_/X _10294_/X _10298_/X vssd1 vssd1 vccd1 vccd1 _10299_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_2_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13141__A1 _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19703_ _19721_/CLK _19703_/D vssd1 vssd1 vccd1 vccd1 _19703_/Q sky130_fd_sc_hd__dfxtp_1
X_16915_ _19736_/Q _19735_/Q _19734_/Q _16915_/D vssd1 vssd1 vccd1 vccd1 _16930_/D
+ sky130_fd_sc_hd__and4_4
XFILLER_66_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12038_ _12038_/A vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18966__D _18966_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17895_ _17903_/B _17899_/B vssd1 vssd1 vccd1 vccd1 _17902_/B sky130_fd_sc_hd__and2b_1
X_19634_ _19637_/CLK _19634_/D vssd1 vssd1 vccd1 vccd1 _19634_/Q sky130_fd_sc_hd__dfxtp_1
X_16846_ _16864_/C _16853_/D _16845_/Y vssd1 vssd1 vccd1 vccd1 _19714_/D sky130_fd_sc_hd__o21a_1
XANTENNA__09991__S1 _09985_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19565_ _19565_/CLK _19565_/D vssd1 vssd1 vccd1 vccd1 _19565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16777_ _19697_/Q _16781_/C _16768_/X vssd1 vssd1 vccd1 vccd1 _16777_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13989_ _13989_/A vssd1 vssd1 vccd1 vccd1 _18629_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13444__A2 _12992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18516_ _19204_/CLK _18516_/D vssd1 vssd1 vccd1 vccd1 _18516_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ _15726_/X _19334_/Q _15747_/S vssd1 vssd1 vccd1 vccd1 _15729_/A sky130_fd_sc_hd__mux2_1
X_19496_ _19498_/CLK _19496_/D vssd1 vssd1 vccd1 vccd1 _19496_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17879__B _17884_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11704__C _12670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18447_ _19938_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_1
X_15659_ _14675_/X _19321_/Q _15659_/S vssd1 vssd1 vccd1 vccd1 _15660_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09180_ _09191_/B vssd1 vssd1 vccd1 vccd1 _11787_/A sky130_fd_sc_hd__clkbuf_2
X_18378_ input64/X vssd1 vssd1 vccd1 vccd1 _18378_/Y sky130_fd_sc_hd__clkinv_8
X_17329_ _11730_/A _11789_/A _11663_/B vssd1 vssd1 vccd1 vccd1 _17392_/A sky130_fd_sc_hd__a21oi_1
XFILLER_147_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13928__A _18295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__S0 _11000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11391__B1 _10655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11143__B1 _10980_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13663__A _15238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16974__A _17073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ _09813_/A vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__buf_2
XANTENNA__11446__A1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__B2 _19922_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09447_ _18288_/A _11663_/B _11663_/C vssd1 vssd1 vccd1 vccd1 _09448_/C sky130_fd_sc_hd__or3_1
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16185__S _16189_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ _16808_/A _16808_/B _20018_/Q _20017_/Q vssd1 vssd1 vccd1 vccd1 _12797_/B
+ sky130_fd_sc_hd__or4bb_2
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18126__A2 _17558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09811__A1 _10161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11340_ _10986_/A _11339_/X _10988_/A vssd1 vssd1 vccd1 vccd1 _11340_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_137_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11271_ _11271_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11271_/X sky130_fd_sc_hd__or2_1
XANTENNA__12742__A input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _14074_/A vssd1 vssd1 vccd1 vccd1 _15061_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10222_ _09860_/A _10221_/X _09696_/A vssd1 vssd1 vccd1 vccd1 _10222_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10804__S0 _10073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _10207_/A _10153_/B vssd1 vssd1 vccd1 vccd1 _10153_/X sky130_fd_sc_hd__or2_1
XFILLER_121_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10084_ _10084_/A vssd1 vssd1 vccd1 vccd1 _10618_/A sky130_fd_sc_hd__clkbuf_2
X_14961_ _19021_/Q _14433_/X _14961_/S vssd1 vssd1 vccd1 vccd1 _14962_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input36_A io_ibus_inst[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09878__A1 _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_16700_ _19787_/Q _19789_/Q _19788_/Q _17074_/A vssd1 vssd1 vccd1 vccd1 _17082_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13912_ _13912_/A vssd1 vssd1 vccd1 vccd1 _18595_/D sky130_fd_sc_hd__clkbuf_1
X_17680_ _17676_/Y _17679_/Y _17741_/S vssd1 vssd1 vccd1 vccd1 _17681_/A sky130_fd_sc_hd__mux2_1
X_14892_ _14640_/X _18990_/Q _14900_/S vssd1 vssd1 vccd1 vccd1 _14893_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16631_ _16631_/A _16636_/C vssd1 vssd1 vccd1 vccd1 _16631_/Y sky130_fd_sc_hd__nor2_1
X_13843_ _13843_/A vssd1 vssd1 vccd1 vccd1 _18567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11093__A _11170_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19350_ _19844_/CLK _19350_/D vssd1 vssd1 vccd1 vccd1 _19350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16562_ _19627_/Q _16564_/C _16561_/Y vssd1 vssd1 vccd1 vccd1 _19627_/D sky130_fd_sc_hd__o21a_1
X_10986_ _10986_/A vssd1 vssd1 vccd1 vccd1 _11216_/A sky130_fd_sc_hd__clkbuf_2
X_13774_ _14599_/A vssd1 vssd1 vccd1 vccd1 _13774_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18301_ _18301_/A vssd1 vssd1 vccd1 vccd1 _18302_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15513_ _19256_/Q _15295_/X _15515_/S vssd1 vssd1 vccd1 vccd1 _15514_/A sky130_fd_sc_hd__mux2_1
X_19281_ _19411_/CLK _19281_/D vssd1 vssd1 vccd1 vccd1 _19281_/Q sky130_fd_sc_hd__dfxtp_1
X_12725_ _19658_/Q vssd1 vssd1 vccd1 vccd1 _16653_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16095__S _16095_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16493_ _19608_/Q _16487_/X _12585_/X _12589_/X _12749_/X vssd1 vssd1 vccd1 vccd1
+ _19608_/D sky130_fd_sc_hd__o221a_1
XFILLER_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18232_ _18232_/A vssd1 vssd1 vccd1 vccd1 _19971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15444_ _15444_/A vssd1 vssd1 vccd1 vccd1 _19225_/D sky130_fd_sc_hd__clkbuf_1
X_12656_ _12657_/A _12656_/B vssd1 vssd1 vccd1 vccd1 _12656_/Y sky130_fd_sc_hd__nor2_8
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18117__A2 _17558_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18163_ _18163_/A vssd1 vssd1 vccd1 vccd1 _19940_/D sky130_fd_sc_hd__clkbuf_1
X_11607_ _13066_/A vssd1 vssd1 vccd1 vccd1 _11607_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11296__S0 _10977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12587_ _17240_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _12587_/X sky130_fd_sc_hd__or2_1
X_15375_ _15443_/S vssd1 vssd1 vccd1 vccd1 _15384_/S sky130_fd_sc_hd__buf_2
XFILLER_168_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17114_ _17122_/A _17114_/B _17114_/C vssd1 vssd1 vccd1 vccd1 _19800_/D sky130_fd_sc_hd__nor3_1
X_14326_ _18775_/Q _13664_/X _14330_/S vssd1 vssd1 vccd1 vccd1 _14327_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17876__A1 _10772_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11538_ _11538_/A _11538_/B _11584_/B _11425_/Y vssd1 vssd1 vccd1 vccd1 _11538_/X
+ sky130_fd_sc_hd__or4b_1
X_18094_ _18054_/X _17696_/Y _18093_/X _18072_/X vssd1 vssd1 vccd1 vccd1 _18094_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15439__S _15439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13748__A _19887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17045_ _17044_/A _17044_/B _19776_/Q vssd1 vssd1 vccd1 vccd1 _17046_/C sky130_fd_sc_hd__a21oi_1
X_14257_ _13796_/X _18745_/Q _14257_/S vssd1 vssd1 vccd1 vccd1 _14258_/A sky130_fd_sc_hd__mux2_1
X_11469_ _09748_/A _11458_/X _11467_/X _09755_/A _11468_/Y vssd1 vssd1 vccd1 vccd1
+ _12668_/B sky130_fd_sc_hd__o32a_4
XFILLER_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12652__A _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13208_ _19748_/Q _12692_/A _13207_/X _12714_/A vssd1 vssd1 vccd1 vccd1 _13208_/X
+ sky130_fd_sc_hd__a211o_1
X_14188_ _13799_/X _18714_/Q _14196_/S vssd1 vssd1 vccd1 vccd1 _14189_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10172__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13139_ _19521_/Q _12799_/Y _13245_/A _19331_/Q vssd1 vssd1 vccd1 vccd1 _13139_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18996_ _19092_/CLK _18996_/D vssd1 vssd1 vccd1 vccd1 _18996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15682__B _17160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17947_ _17945_/B _17949_/A vssd1 vssd1 vccd1 vccd1 _17947_/X sky130_fd_sc_hd__and2b_1
XFILLER_85_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_15_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11220__S0 _11083_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17878_ _17919_/A vssd1 vssd1 vccd1 vccd1 _18002_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19617_ _19620_/CLK _19617_/D vssd1 vssd1 vccd1 vccd1 _19617_/Q sky130_fd_sc_hd__dfxtp_1
X_16829_ _16845_/A _16829_/B vssd1 vssd1 vccd1 vccd1 _16829_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10884__C1 _09975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12099__A _18349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19548_ _19671_/CLK _19548_/D vssd1 vssd1 vccd1 vccd1 _19548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ _09301_/A vssd1 vssd1 vccd1 vccd1 _12664_/A sky130_fd_sc_hd__buf_4
XFILLER_62_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19479_ _19573_/CLK _19479_/D vssd1 vssd1 vccd1 vccd1 _19479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14518__S _14524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09232_ _09271_/C _09271_/B _20025_/Q vssd1 vssd1 vccd1 vccd1 _11648_/C sky130_fd_sc_hd__or3b_4
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15203__A _15203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12928__A1 _11324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14253__S _14257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11364__B1 _09475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10082__A _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09996_ _09996_/A vssd1 vssd1 vccd1 vccd1 _09996_/X sky130_fd_sc_hd__buf_2
XFILLER_103_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14489__A _17041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13393__A _15267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11211__S0 _11083_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11625__B _11625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10840_ _10840_/A _10840_/B vssd1 vssd1 vccd1 vccd1 _10840_/X sky130_fd_sc_hd__or2_1
XANTENNA__12616__B1 _17542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09810__S _10195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18408__B _18408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ _10764_/Y _10766_/Y _10768_/Y _10770_/Y _09717_/A vssd1 vssd1 vccd1 vccd1
+ _10771_/X sky130_fd_sc_hd__o221a_2
XANTENNA__14428__S _14434_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17555__B1 _09419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13332__S _13358_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11641__A _18288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12510_ _19604_/Q _12511_/C _19605_/Q vssd1 vssd1 vccd1 vccd1 _12512_/A sky130_fd_sc_hd__a21oi_1
XFILLER_13_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13490_ input21/X _13318_/X _13436_/X vssd1 vssd1 vccd1 vccd1 _13490_/X sky130_fd_sc_hd__a21o_1
X_12441_ _12538_/A _12436_/Y _12440_/X vssd1 vssd1 vccd1 vccd1 _12441_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11278__S0 _10977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14952__A _14974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15160_ _15160_/A vssd1 vssd1 vccd1 vccd1 _19111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12372_ _17210_/A _12373_/C _19838_/Q vssd1 vssd1 vccd1 vccd1 _12372_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14111_ _14133_/A vssd1 vssd1 vccd1 vccd1 _14120_/S sky130_fd_sc_hd__buf_2
X_11323_ _11199_/A _11322_/X _09609_/B _09617_/A vssd1 vssd1 vccd1 vccd1 _11323_/X
+ sky130_fd_sc_hd__a211o_1
X_15091_ _15091_/A vssd1 vssd1 vccd1 vccd1 _19078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14163__S _14163_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14042_ _18652_/Q _13685_/X _14046_/S vssd1 vssd1 vccd1 vccd1 _14043_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11254_ _09611_/A _11244_/X _11253_/X _09619_/A _19896_/Q vssd1 vssd1 vccd1 vccd1
+ _11254_/Y sky130_fd_sc_hd__a32oi_1
XFILLER_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10205_ _10205_/A _10205_/B _10205_/C vssd1 vssd1 vccd1 vccd1 _10205_/X sky130_fd_sc_hd__or3_2
X_18850_ _19564_/CLK _18850_/D vssd1 vssd1 vccd1 vccd1 _18850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10253__S1 _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11185_ _11178_/A _11184_/X _10920_/A vssd1 vssd1 vccd1 vccd1 _11185_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17801_ _17799_/X _17800_/X _17887_/S vssd1 vssd1 vccd1 vccd1 _17801_/X sky130_fd_sc_hd__mux2_1
X_10136_ _10137_/A _12666_/B vssd1 vssd1 vccd1 vccd1 _11544_/A sky130_fd_sc_hd__or2_1
XFILLER_67_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18781_ _19406_/CLK _18781_/D vssd1 vssd1 vccd1 vccd1 _18781_/Q sky130_fd_sc_hd__dfxtp_1
X_15993_ _13009_/X _19420_/Q _16001_/S vssd1 vssd1 vccd1 vccd1 _15994_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13507__S _13524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11816__A _11816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17732_ _17524_/X _18083_/B _17731_/Y _17667_/A vssd1 vssd1 vccd1 vccd1 _17732_/X
+ sky130_fd_sc_hd__a211o_1
X_14944_ _19013_/Q _14408_/X _14950_/S vssd1 vssd1 vccd1 vccd1 _14945_/A sky130_fd_sc_hd__mux2_1
X_10067_ _09998_/X _10046_/X _10064_/X _10065_/X _10066_/Y vssd1 vssd1 vccd1 vccd1
+ _12665_/B sky130_fd_sc_hd__o32a_4
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_189_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17663_ _17845_/B _17661_/X _17922_/S vssd1 vssd1 vccd1 vccd1 _17664_/A sky130_fd_sc_hd__mux2_1
X_14875_ _14875_/A vssd1 vssd1 vccd1 vccd1 _18982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19402_ _19402_/CLK _19402_/D vssd1 vssd1 vccd1 vccd1 _19402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16614_ _19645_/Q _16611_/B _16613_/Y vssd1 vssd1 vccd1 vccd1 _19645_/D sky130_fd_sc_hd__o21a_1
X_13826_ _13825_/X _18562_/Q _13829_/S vssd1 vssd1 vccd1 vccd1 _13827_/A sky130_fd_sc_hd__mux2_1
X_17594_ _17594_/A vssd1 vssd1 vccd1 vccd1 _17805_/S sky130_fd_sc_hd__buf_2
XFILLER_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11505__S1 _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19333_ _19859_/CLK _19333_/D vssd1 vssd1 vccd1 vccd1 _19333_/Q sky130_fd_sc_hd__dfxtp_1
X_16545_ _16547_/B _16547_/C _16544_/Y vssd1 vssd1 vccd1 vccd1 _19621_/D sky130_fd_sc_hd__o21a_1
X_13757_ _13757_/A vssd1 vssd1 vccd1 vccd1 _18540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10969_ _10969_/A _10969_/B vssd1 vssd1 vccd1 vccd1 _10969_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12647__A _12647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16119__A _16119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12708_ _19814_/Q _17140_/C _12707_/X _19340_/Q vssd1 vssd1 vccd1 vccd1 _12708_/X
+ sky130_fd_sc_hd__a22o_1
X_19264_ _19395_/CLK _19264_/D vssd1 vssd1 vccd1 vccd1 _19264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16476_ _12263_/A _16449_/X _12265_/X _12268_/Y _16468_/X vssd1 vssd1 vccd1 vccd1
+ _19595_/D sky130_fd_sc_hd__o221a_1
X_13688_ _15257_/A vssd1 vssd1 vccd1 vccd1 _14634_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18215_ _18215_/A vssd1 vssd1 vccd1 vccd1 _19963_/D sky130_fd_sc_hd__clkbuf_1
X_15427_ _15427_/A vssd1 vssd1 vccd1 vccd1 _19217_/D sky130_fd_sc_hd__clkbuf_1
X_19195_ _19727_/CLK _19195_/D vssd1 vssd1 vccd1 vccd1 _19195_/Q sky130_fd_sc_hd__dfxtp_1
X_12639_ _12639_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _12639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09956__A _10074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18146_ _16248_/A _19965_/Q _18148_/S vssd1 vssd1 vccd1 vccd1 _18147_/A sky130_fd_sc_hd__mux2_1
X_15358_ _15358_/A vssd1 vssd1 vccd1 vccd1 _15367_/S sky130_fd_sc_hd__buf_4
XFILLER_156_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09882__S0 _09881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14309_ _14309_/A vssd1 vssd1 vccd1 vccd1 _18767_/D sky130_fd_sc_hd__clkbuf_1
X_18077_ _18079_/A _18079_/B _18077_/S vssd1 vssd1 vccd1 vccd1 _18077_/X sky130_fd_sc_hd__mux2_1
X_15289_ _15289_/A vssd1 vssd1 vccd1 vccd1 _15289_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17028_ _17066_/A _17033_/C vssd1 vssd1 vccd1 vccd1 _17028_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11346__B1 _09752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09850_ _10337_/A vssd1 vssd1 vccd1 vccd1 _10392_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_124_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11441__S0 _10625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__A _10988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _09616_/X _09771_/X _09780_/X _09623_/X _19921_/Q vssd1 vssd1 vccd1 vccd1
+ _11537_/A sky130_fd_sc_hd__a32o_2
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _19203_/CLK _18979_/D vssd1 vssd1 vccd1 vccd1 _18979_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10321__B2 _19913_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13941__A _13998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_12_0_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_12_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09215_ _09215_/A _09215_/B vssd1 vssd1 vccd1 vccd1 _17379_/A sky130_fd_sc_hd__nand2_8
XFILLER_167_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10077__A _10817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18244__A _18255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10805__A _10805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11432__S0 _10625_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14711__S _14713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16276__A0 _19527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09979_ _09979_/A vssd1 vssd1 vccd1 vccd1 _09979_/X sky130_fd_sc_hd__buf_2
XFILLER_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18017__A1 _12362_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_190_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _13342_/A vssd1 vssd1 vccd1 vccd1 _12990_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11355__B _12643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11941_ _19584_/Q vssd1 vssd1 vccd1 vccd1 _11974_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _14660_/A vssd1 vssd1 vccd1 vccd1 _14660_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _12366_/A _11864_/Y _11870_/X _11871_/X vssd1 vssd1 vccd1 vccd1 _11872_/Y
+ sky130_fd_sc_hd__a211oi_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _16371_/A vssd1 vssd1 vccd1 vccd1 _15373_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10823_ _11574_/A _10823_/B vssd1 vssd1 vccd1 vccd1 _11575_/A sky130_fd_sc_hd__nor2_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14591_ _14591_/A vssd1 vssd1 vccd1 vccd1 _18868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11371__A _11371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ _19537_/Q _16328_/X _16365_/S vssd1 vssd1 vccd1 vccd1 _16331_/A sky130_fd_sc_hd__mux2_1
X_13542_ _13542_/A vssd1 vssd1 vccd1 vccd1 _18499_/D sky130_fd_sc_hd__clkbuf_1
X_10754_ _10754_/A _10754_/B vssd1 vssd1 vccd1 vccd1 _10754_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10171__S0 _09881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _16265_/A _16265_/C vssd1 vssd1 vccd1 vccd1 _16261_/Y sky130_fd_sc_hd__xnor2_1
X_10685_ _10805_/A _10685_/B vssd1 vssd1 vccd1 vccd1 _10685_/X sky130_fd_sc_hd__or2_1
X_13473_ _13473_/A vssd1 vssd1 vccd1 vccd1 _18495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14682__A _14750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18000_ _18000_/A _18000_/B vssd1 vssd1 vccd1 vccd1 _18002_/C sky130_fd_sc_hd__nor2_1
XFILLER_40_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15212_ _15212_/A vssd1 vssd1 vccd1 vccd1 _15212_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_172_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19837_/CLK sky130_fd_sc_hd__clkbuf_16
X_12424_ _12416_/A _12363_/X _12418_/X _12423_/Y vssd1 vssd1 vccd1 vccd1 _12424_/X
+ sky130_fd_sc_hd__o22a_4
X_16192_ _19509_/Q _14656_/A _16200_/S vssd1 vssd1 vccd1 vccd1 _16193_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15143_ _19103_/Q vssd1 vssd1 vccd1 vccd1 _15144_/A sky130_fd_sc_hd__clkbuf_1
X_12355_ _19978_/Q _11418_/A _17464_/S vssd1 vssd1 vccd1 vccd1 _12356_/A sky130_fd_sc_hd__mux2_4
XFILLER_154_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ _18795_/Q _19130_/Q _11306_/S vssd1 vssd1 vccd1 vccd1 _11306_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15074_ _15131_/S vssd1 vssd1 vccd1 vccd1 _15083_/S sky130_fd_sc_hd__buf_2
X_12286_ _12286_/A vssd1 vssd1 vccd1 vccd1 _12395_/S sky130_fd_sc_hd__buf_2
X_19951_ _19985_/CLK _19951_/D vssd1 vssd1 vccd1 vccd1 _19951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_187_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19859_/CLK sky130_fd_sc_hd__clkbuf_16
X_11237_ _18670_/Q _19165_/Q _11237_/S vssd1 vssd1 vccd1 vccd1 _11237_/X sky130_fd_sc_hd__mux2_1
X_18902_ _19490_/CLK _18902_/D vssd1 vssd1 vccd1 vccd1 _18902_/Q sky130_fd_sc_hd__dfxtp_1
X_14025_ _14025_/A vssd1 vssd1 vccd1 vccd1 _18644_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19882_ _19892_/CLK _19882_/D vssd1 vssd1 vccd1 vccd1 _19882_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12930__A _18127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18833_ _19734_/CLK _18833_/D vssd1 vssd1 vccd1 vccd1 _18833_/Q sky130_fd_sc_hd__dfxtp_1
X_11168_ _11168_/A _11168_/B vssd1 vssd1 vccd1 vccd1 _11168_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10119_ _10909_/S vssd1 vssd1 vccd1 vccd1 _10119_/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_110_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19482_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18764_ _19258_/CLK _18764_/D vssd1 vssd1 vccd1 vccd1 _18764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15976_ _19413_/Q _15279_/X _15984_/S vssd1 vssd1 vccd1 vccd1 _15977_/A sky130_fd_sc_hd__mux2_1
X_11099_ _11153_/A _11099_/B vssd1 vssd1 vccd1 vccd1 _11099_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17715_ _17483_/X _17502_/X _17799_/S vssd1 vssd1 vccd1 vccd1 _17715_/X sky130_fd_sc_hd__mux2_1
X_14927_ _14927_/A vssd1 vssd1 vccd1 vccd1 _19005_/D sky130_fd_sc_hd__clkbuf_1
X_18695_ _19416_/CLK _18695_/D vssd1 vssd1 vccd1 vccd1 _18695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18329__A _18341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15452__S _15456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17646_ _17646_/A vssd1 vssd1 vccd1 vccd1 _17667_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14858_ _14915_/S vssd1 vssd1 vccd1 vccd1 _14867_/S sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_125_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19074_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13809_ _14634_/A vssd1 vssd1 vccd1 vccd1 _13809_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__14068__S _14068_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17577_ _17688_/A vssd1 vssd1 vccd1 vccd1 _17810_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_91_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14789_ _18948_/Q _14420_/X _14797_/S vssd1 vssd1 vccd1 vccd1 _14790_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19316_ _19401_/CLK _19316_/D vssd1 vssd1 vccd1 vccd1 _19316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16528_ _16528_/A _16528_/B _16528_/C vssd1 vssd1 vccd1 vccd1 _19616_/D sky130_fd_sc_hd__nor3_1
XANTENNA__18192__A0 _16361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19247_ _19412_/CLK _19247_/D vssd1 vssd1 vccd1 vccd1 _19247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16459_ _16459_/A vssd1 vssd1 vccd1 vccd1 _19584_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14592__A _14592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19178_ _19405_/CLK _19178_/D vssd1 vssd1 vccd1 vccd1 _19178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18129_ _18129_/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10625__A _10826_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13308__A1 _13060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15627__S _15633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09902_ _18691_/Q _19186_/Q _09902_/S vssd1 vssd1 vccd1 vccd1 _09903_/B sky130_fd_sc_hd__mux2_1
XFILLER_132_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14531__S _14535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20022_ _20027_/CLK _20022_/D vssd1 vssd1 vccd1 vccd1 _20022_/Q sky130_fd_sc_hd__dfxtp_1
X_09833_ _09833_/A _09833_/B vssd1 vssd1 vccd1 vccd1 _09833_/X sky130_fd_sc_hd__or2_1
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12819__A0 _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _10161_/A _09763_/X _09567_/A vssd1 vssd1 vccd1 vccd1 _09764_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10360__A _19913_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09695_ _09695_/A vssd1 vssd1 vccd1 vccd1 _09696_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13492__B1 _19953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13671__A _15244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10845__A2 _19555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12047__A1 _10821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12287__A _12395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_137_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11007__C1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10470_ _11428_/S vssd1 vssd1 vccd1 vccd1 _10470_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13547__B2 _19545_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ _17903_/B _12140_/B vssd1 vssd1 vccd1 vccd1 _12143_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__15839__A3 _15819_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15537__S _15539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12071_ _18349_/A _17381_/A _12099_/B _12070_/X vssd1 vssd1 vccd1 vccd1 _12071_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10208__S1 _09809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11022_ _09473_/A _11014_/X _11016_/X _11021_/X _09601_/A vssd1 vssd1 vccd1 vccd1
+ _11022_/X sky130_fd_sc_hd__a311o_2
XFILLER_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13057__S _13090_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11366__A _11440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15830_ _15829_/X _19352_/Q _15835_/S vssd1 vssd1 vccd1 vccd1 _15831_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _19910_/Q _12772_/B _15800_/S vssd1 vssd1 vccd1 vccd1 _15761_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12973_ _17861_/A vssd1 vssd1 vccd1 vccd1 _12973_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_42_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19311_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _17498_/X _17499_/X _17500_/S vssd1 vssd1 vccd1 vccd1 _17500_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _14712_/A vssd1 vssd1 vccd1 vccd1 _18909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _19431_/CLK _18480_/D vssd1 vssd1 vccd1 vccd1 _18480_/Q sky130_fd_sc_hd__dfxtp_1
X_11924_ _11924_/A vssd1 vssd1 vccd1 vccd1 _11924_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _15692_/A vssd1 vssd1 vccd1 vccd1 _19329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17431_ _17431_/A vssd1 vssd1 vccd1 vccd1 _17702_/B sky130_fd_sc_hd__clkbuf_2
X_14643_ _14643_/A vssd1 vssd1 vccd1 vccd1 _18884_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17988__A _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _11704_/X _11853_/X _11854_/X _12320_/B vssd1 vssd1 vccd1 vccd1 _11855_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output105_A _11673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15775__A2 _13370_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11305__S _11305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10806_ _18645_/Q _19236_/Q _19398_/Q _18613_/Q _10081_/X _10691_/A vssd1 vssd1 vccd1
+ vccd1 _10806_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17362_ _17362_/A vssd1 vssd1 vccd1 vccd1 _19887_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_57_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19952_/CLK sky130_fd_sc_hd__clkbuf_16
X_14574_ _14574_/A vssd1 vssd1 vccd1 vccd1 _14574_/X sky130_fd_sc_hd__clkbuf_2
X_11786_ _11786_/A vssd1 vssd1 vccd1 vccd1 _18283_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19101_ _19455_/CLK _19101_/D vssd1 vssd1 vccd1 vccd1 _19101_/Q sky130_fd_sc_hd__dfxtp_1
X_16313_ _16313_/A _16321_/D vssd1 vssd1 vccd1 vccd1 _16313_/X sky130_fd_sc_hd__and2_1
X_13525_ _13525_/A vssd1 vssd1 vccd1 vccd1 _18498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10737_ _19109_/Q _18875_/Q _19557_/Q _19205_/Q _10614_/X _10682_/X vssd1 vssd1 vccd1
+ vccd1 _10737_/X sky130_fd_sc_hd__mux4_2
X_17293_ _17304_/A vssd1 vssd1 vccd1 vccd1 _17302_/S sky130_fd_sc_hd__buf_2
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14616__S _14622_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19032_ _19288_/CLK _19032_/D vssd1 vssd1 vccd1 vccd1 _19032_/Q sky130_fd_sc_hd__dfxtp_1
X_16244_ _16248_/A _16248_/C vssd1 vssd1 vccd1 vccd1 _16244_/Y sky130_fd_sc_hd__xnor2_2
X_13456_ _13456_/A vssd1 vssd1 vccd1 vccd1 _18494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10668_ _10660_/Y _10662_/Y _10664_/Y _10667_/Y _09717_/A vssd1 vssd1 vccd1 vccd1
+ _10668_/X sky130_fd_sc_hd__o221a_1
XFILLER_12_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12644__B _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12407_ _12407_/A vssd1 vssd1 vccd1 vccd1 _18036_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__10447__S1 _10326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16175_ _16175_/A vssd1 vssd1 vccd1 vccd1 _19501_/D sky130_fd_sc_hd__clkbuf_1
X_10599_ _19908_/Q vssd1 vssd1 vccd1 vccd1 _10599_/Y sky130_fd_sc_hd__inv_2
X_13387_ _19727_/Q _13341_/X _13342_/X _19695_/Q _13386_/X vssd1 vssd1 vccd1 vccd1
+ _13387_/X sky130_fd_sc_hd__a221o_2
XFILLER_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput107 _09188_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_st_type[0] sky130_fd_sc_hd__buf_2
X_15126_ _15126_/A vssd1 vssd1 vccd1 vccd1 _19094_/D sky130_fd_sc_hd__clkbuf_1
Xoutput118 _12655_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[18] sky130_fd_sc_hd__buf_2
XANTENNA__12761__A2 _13560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput129 _12667_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[28] sky130_fd_sc_hd__buf_2
X_12338_ _12338_/A _16474_/A _12338_/C vssd1 vssd1 vccd1 vccd1 _12339_/D sky130_fd_sc_hd__and3_1
XFILLER_142_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18969__D _18969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19934_ _19938_/CLK _19934_/D vssd1 vssd1 vccd1 vccd1 _19934_/Q sky130_fd_sc_hd__dfxtp_1
X_15057_ _19064_/Q _14468_/X _15059_/S vssd1 vssd1 vccd1 vccd1 _15058_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12660__A _12663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ _12263_/A _12115_/X _12265_/X _12268_/Y vssd1 vssd1 vccd1 vccd1 _12269_/X
+ sky130_fd_sc_hd__o22a_4
X_14008_ _14008_/A vssd1 vssd1 vccd1 vccd1 _18636_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19865_ _19865_/CLK _19865_/D vssd1 vssd1 vccd1 vccd1 _19865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18816_ _19504_/CLK _18816_/D vssd1 vssd1 vccd1 vccd1 _18816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19796_ _19803_/CLK _19796_/D vssd1 vssd1 vccd1 vccd1 _19796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18747_ _19306_/CLK _18747_/D vssd1 vssd1 vccd1 vccd1 _18747_/Q sky130_fd_sc_hd__dfxtp_1
X_15959_ _15959_/A vssd1 vssd1 vccd1 vccd1 _19405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18678_ _18845_/CLK _18678_/D vssd1 vssd1 vccd1 vccd1 _18678_/Q sky130_fd_sc_hd__dfxtp_1
X_09480_ _18967_/Q vssd1 vssd1 vccd1 vccd1 _11274_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10383__S0 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13226__A0 _19904_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17629_ _17604_/B _17628_/Y _17649_/A vssd1 vssd1 vccd1 vccd1 _17629_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15910__S _15912_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17138__A input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20005_ _20048_/CLK _20005_/D vssd1 vssd1 vccd1 vccd1 _20005_/Q sky130_fd_sc_hd__dfxtp_1
X_09816_ _10312_/A vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__buf_2
XANTENNA__15881__A _15903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10090__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10610__S1 _10609_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16651__B1 _16624_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09747_ _09998_/A vssd1 vssd1 vccd1 vccd1 _09748_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15092__S _15094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09678_ _10051_/A vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__buf_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10374__S0 _10416_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11640_ _11640_/A _11723_/B _11640_/C vssd1 vssd1 vccd1 vccd1 _11641_/D sky130_fd_sc_hd__or3_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10126__S0 _11449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11779__B1 _12492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11571_ _10728_/A _11570_/Y _11408_/Y vssd1 vssd1 vccd1 vccd1 _11571_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_156_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13310_ _18485_/Q _13309_/X _13358_/S vssd1 vssd1 vccd1 vccd1 _13311_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10522_ _19500_/Q _18912_/Q _18949_/Q _18523_/Q _10470_/X _10462_/A vssd1 vssd1 vccd1
+ vccd1 _10523_/B sky130_fd_sc_hd__mux4_1
X_14290_ _13844_/X _18760_/Q _14290_/S vssd1 vssd1 vccd1 vccd1 _14291_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13241_ _13241_/A vssd1 vssd1 vccd1 vccd1 _18481_/D sky130_fd_sc_hd__clkbuf_1
X_10453_ _19470_/Q _19308_/Q _18717_/Q _18487_/Q _10325_/X _10497_/A vssd1 vssd1 vccd1
+ vccd1 _10453_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17747__S _18109_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10429__S1 _10291_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input66_A io_ibus_valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ _10428_/A _10384_/B vssd1 vssd1 vccd1 vccd1 _10384_/X sky130_fd_sc_hd__or2_1
XFILLER_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13172_ _13172_/A vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17131__A1 _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17048__A _17066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13576__A _16268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ _12492_/A vssd1 vssd1 vccd1 vccd1 _12123_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17980_ _17619_/X _17894_/X _17979_/X vssd1 vssd1 vccd1 vccd1 _17980_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12480__A _12480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16931_ _16946_/A _16965_/C vssd1 vssd1 vccd1 vccd1 _16931_/Y sky130_fd_sc_hd__nor2_1
X_12054_ _12002_/A _12002_/B _12021_/A _12021_/B _12053_/Y vssd1 vssd1 vccd1 vccd1
+ _12055_/B sky130_fd_sc_hd__a41o_2
XFILLER_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15791__A _15806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11005_ _10084_/A _11004_/X _11204_/A vssd1 vssd1 vccd1 vccd1 _11005_/X sky130_fd_sc_hd__a21o_1
X_16862_ _16865_/A _16870_/D _16861_/Y vssd1 vssd1 vccd1 vccd1 _19719_/D sky130_fd_sc_hd__o21a_1
X_19650_ _19782_/CLK _19650_/D vssd1 vssd1 vccd1 vccd1 _19650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15813_ _18463_/Q _13577_/X _15812_/X vssd1 vssd1 vccd1 vccd1 _17228_/A sky130_fd_sc_hd__a21oi_2
X_18601_ _19203_/CLK _18601_/D vssd1 vssd1 vccd1 vccd1 _18601_/Q sky130_fd_sc_hd__dfxtp_1
X_19581_ _20000_/CLK _19581_/D vssd1 vssd1 vccd1 vccd1 _19581_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16098__S _16106_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16793_ _16818_/A _16793_/B vssd1 vssd1 vccd1 vccd1 _16793_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18532_ _19027_/CLK _18532_/D vssd1 vssd1 vccd1 vccd1 _18532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11467__C1 _09717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15744_ _18451_/Q _13577_/X _15743_/X vssd1 vssd1 vccd1 vccd1 _17191_/A sky130_fd_sc_hd__a21oi_4
X_12956_ _18448_/Q _12951_/X _12076_/A _12954_/X vssd1 vssd1 vccd1 vccd1 _18448_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12639__B _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _19952_/CLK _18463_/D vssd1 vssd1 vccd1 vccd1 _18463_/Q sky130_fd_sc_hd__dfxtp_2
X_11907_ _11933_/C _11907_/B vssd1 vssd1 vccd1 vccd1 _11907_/X sky130_fd_sc_hd__xor2_4
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _19896_/Q _15668_/X _13597_/B vssd1 vssd1 vccd1 vccd1 _15675_/X sky130_fd_sc_hd__a21o_1
X_12887_ _12887_/A vssd1 vssd1 vccd1 vccd1 _12887_/X sky130_fd_sc_hd__buf_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15730__S _15757_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17414_ _17414_/A vssd1 vssd1 vccd1 vccd1 _17586_/S sky130_fd_sc_hd__buf_2
X_14626_ _14624_/X _18879_/Q _14638_/S vssd1 vssd1 vccd1 vccd1 _14627_/A sky130_fd_sc_hd__mux2_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11838_ _19771_/Q vssd1 vssd1 vccd1 vccd1 _12914_/A sky130_fd_sc_hd__clkbuf_2
X_18394_ input38/X vssd1 vssd1 vccd1 vccd1 _18394_/Y sky130_fd_sc_hd__inv_6
XFILLER_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18326__B _18326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17345_ _17345_/A vssd1 vssd1 vccd1 vccd1 _19883_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _13828_/X _18856_/Q _14557_/S vssd1 vssd1 vccd1 vccd1 _14558_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11769_ _12066_/B vssd1 vssd1 vccd1 vccd1 _16487_/A sky130_fd_sc_hd__buf_2
XANTENNA__12655__A _12657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13508_ _13508_/A vssd1 vssd1 vccd1 vccd1 _18497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17276_ _12874_/X _19862_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17277_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14488_ _17339_/A _14485_/X _14486_/X _14487_/Y vssd1 vssd1 vccd1 vccd1 _18409_/B
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__10993__A1 _11216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19015_ _19366_/CLK _19015_/D vssd1 vssd1 vccd1 vccd1 _19015_/Q sky130_fd_sc_hd__dfxtp_1
X_16227_ _15688_/X _16225_/Y _16262_/S vssd1 vssd1 vccd1 vccd1 _16227_/X sky130_fd_sc_hd__mux2_1
X_13439_ _13428_/A _13438_/C _19950_/Q vssd1 vssd1 vccd1 vccd1 _13439_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_162_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16158_ _16204_/S vssd1 vssd1 vccd1 vccd1 _16167_/S sky130_fd_sc_hd__buf_2
XANTENNA__11942__B1 _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15109_ _15109_/A vssd1 vssd1 vccd1 vccd1 _19086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16089_ _13230_/X _19463_/Q _16095_/S vssd1 vssd1 vccd1 vccd1 _16090_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19917_ _19986_/CLK _19917_/D vssd1 vssd1 vccd1 vccd1 _19917_/Q sky130_fd_sc_hd__dfxtp_4
X_19848_ _19881_/CLK _19848_/D vssd1 vssd1 vccd1 vccd1 _19848_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09601_ _09601_/A vssd1 vssd1 vccd1 vccd1 _09602_/A sky130_fd_sc_hd__buf_2
XANTENNA__16633__B1 _16624_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19779_ _19783_/CLK _19779_/D vssd1 vssd1 vccd1 vccd1 _19779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19323__D _19323_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ _09532_/A vssd1 vssd1 vccd1 vccd1 _10811_/S sky130_fd_sc_hd__buf_4
XFILLER_37_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15206__A _15206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18386__B1 _18374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ _12933_/A vssd1 vssd1 vccd1 vccd1 _18028_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17421__A _17421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09394_ _09394_/A _13136_/B vssd1 vssd1 vccd1 vccd1 _09394_/X sky130_fd_sc_hd__or2_1
XFILLER_40_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10659__S1 _10014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09874__A _09887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10736__A1 _09813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10813__A _10813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15675__A1 _19896_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12489__A1 _19540_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ _17247_/B _12810_/B vssd1 vssd1 vccd1 vccd1 _12810_/Y sky130_fd_sc_hd__nor2_4
XFILLER_47_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11644__A _11704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13790_ _14615_/A vssd1 vssd1 vccd1 vccd1 _13790_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12741_ _12732_/X _12735_/X _12738_/Y _13577_/A _18453_/Q vssd1 vssd1 vccd1 vccd1
+ _12741_/X sky130_fd_sc_hd__a32o_4
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18427__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15460_ _15460_/A vssd1 vssd1 vccd1 vccd1 _19231_/D sky130_fd_sc_hd__clkbuf_1
X_12672_ _12672_/A vssd1 vssd1 vccd1 vccd1 _12673_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14615_/A vssd1 vssd1 vccd1 vccd1 _14411_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _17392_/B _17391_/A vssd1 vssd1 vccd1 vccd1 _11623_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14166__S _14174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15391_ _14599_/X _19201_/Q _15395_/S vssd1 vssd1 vccd1 vccd1 _15392_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12475__A _12475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13070__S _13090_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17130_ _17130_/A vssd1 vssd1 vccd1 vccd1 _19810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14342_ _14342_/A vssd1 vssd1 vccd1 vccd1 _18782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11554_ _11554_/A _11554_/B vssd1 vssd1 vccd1 vccd1 _11554_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17985__B _17985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10505_ _09709_/A _10498_/X _10500_/Y _10504_/Y _09740_/A vssd1 vssd1 vccd1 vccd1
+ _10505_/X sky130_fd_sc_hd__o311a_1
XFILLER_128_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17061_ _17062_/A _17062_/C _17060_/Y vssd1 vssd1 vccd1 vccd1 _19781_/D sky130_fd_sc_hd__o21a_1
X_14273_ _13819_/X _18752_/Q _14279_/S vssd1 vssd1 vccd1 vccd1 _14274_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11485_ _19128_/Q _18894_/Q _19576_/Q _19224_/Q _10812_/S _09514_/A vssd1 vssd1 vccd1
+ vccd1 _11485_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _13195_/X _19429_/Q _16012_/S vssd1 vssd1 vccd1 vccd1 _16013_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12716__A2 _13142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13224_ _16265_/A _13225_/B _13066_/A vssd1 vssd1 vccd1 vccd1 _13224_/Y sky130_fd_sc_hd__o21ai_1
X_10436_ _10436_/A _10436_/B vssd1 vssd1 vccd1 vccd1 _10436_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output172_A _16461_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12922__B _18461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13155_ _12837_/A _12818_/B _13154_/Y vssd1 vssd1 vccd1 vccd1 _13155_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10367_ _18686_/Q _19181_/Q _10367_/S vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__mux2_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12106_ _17884_/A _12106_/B vssd1 vssd1 vccd1 vccd1 _12108_/A sky130_fd_sc_hd__xnor2_2
XFILLER_151_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11538__B _11538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10298_ _09520_/A _10295_/X _10478_/A vssd1 vssd1 vccd1 vccd1 _10298_/X sky130_fd_sc_hd__a21o_1
XFILLER_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13147_/S sky130_fd_sc_hd__buf_2
XFILLER_88_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17963_ _17976_/A _17963_/B vssd1 vssd1 vccd1 vccd1 _17965_/C sky130_fd_sc_hd__nor2_1
XFILLER_78_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19702_ _19721_/CLK _19702_/D vssd1 vssd1 vccd1 vccd1 _19702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16914_ _16925_/B _16918_/D _19736_/Q vssd1 vssd1 vccd1 vccd1 _16916_/B sky130_fd_sc_hd__a21oi_1
X_12037_ _12037_/A _12037_/B vssd1 vssd1 vccd1 vccd1 _12038_/A sky130_fd_sc_hd__and2_2
X_17894_ _17600_/X _17664_/Y _17530_/A vssd1 vssd1 vccd1 vccd1 _17894_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16615__B1 _16577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19633_ _19637_/CLK _19633_/D vssd1 vssd1 vccd1 vccd1 _19633_/Q sky130_fd_sc_hd__dfxtp_1
X_16845_ _16845_/A _16845_/B vssd1 vssd1 vccd1 vccd1 _16845_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19564_ _19564_/CLK _19564_/D vssd1 vssd1 vccd1 vccd1 _19564_/Q sky130_fd_sc_hd__dfxtp_1
X_16776_ _19696_/Q _16774_/B _16775_/Y vssd1 vssd1 vccd1 vccd1 _19696_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10338__S0 _10337_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13988_ _18629_/Q _13723_/X _13994_/S vssd1 vssd1 vccd1 vccd1 _13989_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15727_ _15844_/S vssd1 vssd1 vccd1 vccd1 _15747_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_18_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18515_ _19493_/CLK _18515_/D vssd1 vssd1 vccd1 vccd1 _18515_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _18319_/A _11808_/X _12942_/S vssd1 vssd1 vccd1 vccd1 _12939_/X sky130_fd_sc_hd__mux2_1
X_19495_ _19495_/CLK _19495_/D vssd1 vssd1 vccd1 vccd1 _19495_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15658_ _15658_/A vssd1 vssd1 vccd1 vccd1 _19320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18446_ _19930_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09959__A _11204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14609_ _14676_/S vssd1 vssd1 vccd1 vccd1 _14622_/S sky130_fd_sc_hd__buf_6
XFILLER_61_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18377_ _18380_/A _18377_/B vssd1 vssd1 vccd1 vccd1 _20028_/D sky130_fd_sc_hd__nor2_1
X_15589_ _16062_/B _15589_/B vssd1 vssd1 vccd1 vccd1 _15646_/A sky130_fd_sc_hd__or2_4
XANTENNA__12385__A _12385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17328_ _17323_/A _17327_/A _12594_/C _17327_/Y vssd1 vssd1 vccd1 vccd1 _17335_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_119_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_11_clock_A _19998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17343__A1 _18301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17895__B _17899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17259_ _17259_/A vssd1 vssd1 vccd1 vccd1 _19854_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14804__S _14808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09694__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11066__S1 _11065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11143__A1 _10899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18071__A2 _17743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11464__A _11464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09515_ _09515_/A vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__buf_8
XFILLER_71_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _17331_/B _11789_/C vssd1 vssd1 vccd1 vccd1 _11663_/C sky130_fd_sc_hd__or2_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09377_ _13527_/B _13077_/B _12888_/A _12989_/A vssd1 vssd1 vccd1 vccd1 _09377_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10501__S0 _10392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09808__S _10195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11270_ _19485_/Q _18897_/Q _18934_/Q _18508_/Q _11262_/X _11059_/A vssd1 vssd1 vccd1
+ vccd1 _11271_/B sky130_fd_sc_hd__mux4_2
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10221_ _19120_/Q _18886_/Q _19568_/Q _19216_/Q _09653_/A _09927_/A vssd1 vssd1 vccd1
+ vccd1 _10221_/X sky130_fd_sc_hd__mux4_2
XFILLER_152_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10804__S1 _10609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14015__A _14072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10152_ _19379_/Q _18993_/Q _19443_/Q _18562_/Q _10162_/S _10196_/A vssd1 vssd1 vccd1
+ vccd1 _10153_/B sky130_fd_sc_hd__mux4_1
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14960_ _14960_/A vssd1 vssd1 vccd1 vccd1 _19020_/D sky130_fd_sc_hd__clkbuf_1
X_10083_ _10083_/A vssd1 vssd1 vccd1 vccd1 _10084_/A sky130_fd_sc_hd__buf_4
XFILLER_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11134__A1 _10875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__buf_2
XFILLER_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13911_ _13828_/X _18595_/Q _13911_/S vssd1 vssd1 vccd1 vccd1 _13912_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input29_A io_dbus_rdata[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ _14902_/A vssd1 vssd1 vccd1 vccd1 _14900_/S sky130_fd_sc_hd__buf_2
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16630_ _16630_/A vssd1 vssd1 vccd1 vccd1 _16636_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13842_ _13841_/X _18567_/Q _13845_/S vssd1 vssd1 vccd1 vccd1 _13843_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16561_ _19627_/Q _16564_/C _16533_/X vssd1 vssd1 vccd1 vccd1 _16561_/Y sky130_fd_sc_hd__a21oi_1
X_13773_ _13773_/A vssd1 vssd1 vccd1 vccd1 _18545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16376__S _16382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10985_ _11025_/A _10985_/B vssd1 vssd1 vccd1 vccd1 _10985_/Y sky130_fd_sc_hd__nor2_1
X_15512_ _15512_/A vssd1 vssd1 vccd1 vccd1 _19255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17022__B1 _17021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18300_ _20032_/Q _18291_/X _18299_/Y _18289_/X vssd1 vssd1 vccd1 vccd1 _20000_/D
+ sky130_fd_sc_hd__o211a_1
X_19280_ _19906_/CLK _19280_/D vssd1 vssd1 vccd1 vccd1 _19280_/Q sky130_fd_sc_hd__dfxtp_1
X_12724_ _16921_/C _12719_/X _12723_/X _19690_/Q vssd1 vssd1 vccd1 vccd1 _13301_/C
+ sky130_fd_sc_hd__a22o_2
XFILLER_16_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16492_ _12561_/A _16487_/X _12563_/X _12566_/Y _12749_/X vssd1 vssd1 vccd1 vccd1
+ _19607_/D sky130_fd_sc_hd__o221a_1
XFILLER_71_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10740__S0 _10608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18231_ _19971_/Q hold18/X _18231_/S vssd1 vssd1 vccd1 vccd1 _18232_/A sky130_fd_sc_hd__mux2_1
X_15443_ _14675_/X _19225_/Q _15443_/S vssd1 vssd1 vccd1 vccd1 _15444_/A sky130_fd_sc_hd__mux2_1
X_12655_ _12657_/A _12655_/B vssd1 vssd1 vccd1 vccd1 _12655_/Y sky130_fd_sc_hd__nor2_4
XFILLER_169_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10718__A _10718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11606_ _18929_/Q vssd1 vssd1 vccd1 vccd1 _13066_/A sky130_fd_sc_hd__clkbuf_2
X_18162_ _13282_/A _19972_/Q _18170_/S vssd1 vssd1 vccd1 vccd1 _18163_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15374_ _15430_/A vssd1 vssd1 vccd1 vccd1 _15443_/S sky130_fd_sc_hd__buf_4
XFILLER_12_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12586_ _19847_/Q vssd1 vssd1 vccd1 vccd1 _17240_/A sky130_fd_sc_hd__buf_2
XANTENNA__11296__S1 _10006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_185_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17113_ _17112_/A _17112_/C _19800_/Q vssd1 vssd1 vccd1 vccd1 _17114_/C sky130_fd_sc_hd__a21oi_1
X_14325_ _14325_/A vssd1 vssd1 vccd1 vccd1 _18774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11537_ _11537_/A _12667_/B _11538_/A vssd1 vssd1 vccd1 vccd1 _11537_/X sky130_fd_sc_hd__or3_1
X_18093_ _17781_/X _17691_/X _18092_/X _17796_/X vssd1 vssd1 vccd1 vccd1 _18093_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17876__A2 _17861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12933__A _12933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17044_ _17044_/A _17044_/B _19776_/Q vssd1 vssd1 vccd1 vccd1 _17046_/B sky130_fd_sc_hd__and3_1
XANTENNA_output97_A _11864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14256_ _14256_/A vssd1 vssd1 vccd1 vccd1 _18744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11468_ _19922_/Q vssd1 vssd1 vccd1 vccd1 _11468_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13748__B _13748_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13207_ _19334_/Q _12759_/X _12758_/A _19524_/Q _13206_/X vssd1 vssd1 vccd1 vccd1
+ _13207_/X sky130_fd_sc_hd__a221o_1
X_10419_ _09899_/A _10416_/X _10418_/X vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__a21o_1
X_14187_ _14209_/A vssd1 vssd1 vccd1 vccd1 _14196_/S sky130_fd_sc_hd__buf_2
X_11399_ _11399_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11399_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13138_ _19857_/Q _12992_/A _12893_/B _19810_/Q _13137_/X vssd1 vssd1 vccd1 vccd1
+ _13138_/X sky130_fd_sc_hd__a221o_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _19571_/CLK _18995_/D vssd1 vssd1 vccd1 vccd1 _18995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13764__A _14589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17236__A _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _15209_/A vssd1 vssd1 vccd1 vccd1 _13069_/X sky130_fd_sc_hd__clkbuf_1
X_17946_ _17945_/A _17949_/A _17814_/X _17945_/Y vssd1 vssd1 vccd1 vccd1 _17946_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13483__B _13483_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11676__A2 _12606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__S1 _11164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17877_ _17627_/X _17681_/A _17719_/X vssd1 vssd1 vccd1 vccd1 _17877_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17261__A0 _15688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19616_ _19620_/CLK _19616_/D vssd1 vssd1 vccd1 vccd1 _19616_/Q sky130_fd_sc_hd__dfxtp_1
X_16828_ _19710_/Q _16863_/C vssd1 vssd1 vccd1 vccd1 _16829_/B sky130_fd_sc_hd__and2_1
XFILLER_65_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19547_ _19726_/CLK _19547_/D vssd1 vssd1 vccd1 vccd1 _19547_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12625__A1 _12621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16759_ _19690_/Q _16757_/B _16758_/Y vssd1 vssd1 vccd1 vccd1 _19690_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13703__S _13715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09300_ _09426_/A _09329_/A _12594_/B vssd1 vssd1 vccd1 vccd1 _17381_/A sky130_fd_sc_hd__or3_4
XFILLER_62_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10636__B1 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19478_ _19478_/CLK _19478_/D vssd1 vssd1 vccd1 vccd1 _19478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10731__S0 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09231_ _20033_/Q vssd1 vssd1 vccd1 vccd1 _11523_/A sky130_fd_sc_hd__inv_2
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18429_ _18435_/A _18429_/B vssd1 vssd1 vccd1 vccd1 _20050_/D sky130_fd_sc_hd__nor2_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13050__A1 _13588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16315__A _16315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18277__C1 _17243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11364__A1 _10730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09995_ _09979_/X _09987_/X _09989_/X _09994_/X _09602_/A vssd1 vssd1 vccd1 vccd1
+ _09995_/X sky130_fd_sc_hd__a311o_1
XANTENNA__15365__S _15367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17146__A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11211__S1 _11164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16196__S _16200_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14709__S _14713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10770_ _10757_/A _10769_/X _10655_/X vssd1 vssd1 vccd1 vccd1 _10770_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17555__A1 _12675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09429_ _12099_/B vssd1 vssd1 vccd1 vccd1 _12942_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12440_ _11818_/X _11819_/X _12439_/Y _11977_/X vssd1 vssd1 vccd1 vccd1 _12440_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_100_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11278__S1 _10006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__B1 _11352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12371_ _12366_/X _12367_/Y _12370_/Y vssd1 vssd1 vccd1 vccd1 _12371_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14110_ _14110_/A vssd1 vssd1 vccd1 vccd1 _18681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11322_ _09470_/A _11315_/Y _11317_/Y _11319_/Y _11321_/Y vssd1 vssd1 vccd1 vccd1
+ _11322_/X sky130_fd_sc_hd__o32a_2
XFILLER_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15090_ _14615_/X _19078_/Q _15094_/S vssd1 vssd1 vccd1 vccd1 _15091_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14041_ _14041_/A vssd1 vssd1 vccd1 vccd1 _18651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11253_ _11246_/X _11248_/X _11250_/X _11252_/X _09600_/A vssd1 vssd1 vccd1 vccd1
+ _11253_/X sky130_fd_sc_hd__a221o_2
XFILLER_107_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10789__S0 _10751_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ _10209_/A _10201_/X _10203_/X _09826_/X vssd1 vssd1 vccd1 vccd1 _10205_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15783__B _18458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ _19454_/Q _19292_/Q _18701_/Q _18471_/Q _11161_/X _10974_/A vssd1 vssd1 vccd1
+ vccd1 _11184_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17800_ _17673_/X _17686_/X _17800_/S vssd1 vssd1 vccd1 vccd1 _17800_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10135_ _09998_/X _10123_/X _10133_/X _10065_/X _10134_/Y vssd1 vssd1 vccd1 vccd1
+ _12666_/B sky130_fd_sc_hd__o32a_4
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18780_ _19406_/CLK _18780_/D vssd1 vssd1 vccd1 vccd1 _18780_/Q sky130_fd_sc_hd__dfxtp_1
X_15992_ _16060_/S vssd1 vssd1 vccd1 vccd1 _16001_/S sky130_fd_sc_hd__clkbuf_4
X_14943_ _14943_/A vssd1 vssd1 vccd1 vccd1 _19012_/D sky130_fd_sc_hd__clkbuf_1
X_10066_ _19919_/Q vssd1 vssd1 vccd1 vccd1 _10066_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17731_ _17723_/X _17728_/Y _17730_/X vssd1 vssd1 vccd1 vccd1 _17731_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_85_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output135_A _12636_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14874_ _14615_/X _18982_/Q _14878_/S vssd1 vssd1 vccd1 vccd1 _14875_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17662_ _17662_/A vssd1 vssd1 vccd1 vccd1 _17922_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19401_ _19401_/CLK _19401_/D vssd1 vssd1 vccd1 vccd1 _19401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13825_ _14650_/A vssd1 vssd1 vccd1 vccd1 _13825_/X sky130_fd_sc_hd__clkbuf_1
X_16613_ _16631_/A _16617_/C vssd1 vssd1 vccd1 vccd1 _16613_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12607__A1 _11601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17593_ _17585_/X _17592_/X _17810_/S vssd1 vssd1 vccd1 vccd1 _17593_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14619__S _14622_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11832__A _19819_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19332_ _19620_/CLK _19332_/D vssd1 vssd1 vccd1 vccd1 _19332_/Q sky130_fd_sc_hd__dfxtp_1
X_16544_ _16547_/B _16547_/C _16533_/X vssd1 vssd1 vccd1 vccd1 _16544_/Y sky130_fd_sc_hd__a21oi_1
X_13756_ _13755_/X _18540_/Q _13765_/S vssd1 vssd1 vccd1 vccd1 _13757_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10968_ _18802_/Q _19137_/Q _10968_/S vssd1 vssd1 vccd1 vccd1 _10969_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13280__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12647__B _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ _13245_/A vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__clkbuf_2
X_19263_ _19391_/CLK _19263_/D vssd1 vssd1 vccd1 vccd1 _19263_/Q sky130_fd_sc_hd__dfxtp_1
X_16475_ _16474_/Y _12494_/A _12243_/X _12248_/Y _12908_/X vssd1 vssd1 vccd1 vccd1
+ _19594_/D sky130_fd_sc_hd__a221oi_1
X_13687_ _13687_/A vssd1 vssd1 vccd1 vccd1 _18524_/D sky130_fd_sc_hd__clkbuf_1
X_10899_ _10899_/A vssd1 vssd1 vccd1 vccd1 _10929_/A sky130_fd_sc_hd__clkbuf_2
X_15426_ _14650_/X _19217_/Q _15428_/S vssd1 vssd1 vccd1 vccd1 _15427_/A sky130_fd_sc_hd__mux2_1
X_18214_ _19963_/Q _11974_/A _18220_/S vssd1 vssd1 vccd1 vccd1 _18215_/A sky130_fd_sc_hd__mux2_1
X_19194_ _19196_/CLK _19194_/D vssd1 vssd1 vccd1 vccd1 _19194_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13032__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12638_ _12639_/A _12638_/B vssd1 vssd1 vccd1 vccd1 _12638_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__13032__B2 _13007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15357_ _15357_/A vssd1 vssd1 vccd1 vccd1 _19186_/D sky130_fd_sc_hd__clkbuf_1
X_18145_ _18145_/A vssd1 vssd1 vccd1 vccd1 _19932_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12663__A _12663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ _12473_/X _12669_/B _12474_/X _12568_/X vssd1 vssd1 vccd1 vccd1 _18111_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16135__A _16191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09882__S1 _09874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14308_ _18767_/Q _13630_/X _14308_/S vssd1 vssd1 vccd1 vccd1 _14309_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18076_ _18079_/A _18079_/B vssd1 vssd1 vccd1 vccd1 _18076_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15288_ _15288_/A vssd1 vssd1 vccd1 vccd1 _19157_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17027_ _19765_/Q _19764_/Q _17027_/C _17027_/D vssd1 vssd1 vccd1 vccd1 _17033_/C
+ sky130_fd_sc_hd__and4_1
X_14239_ _14239_/A vssd1 vssd1 vccd1 vccd1 _18736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11346__A1 _09745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11346__B2 _09342_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11441__S1 _10604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11897__A2 _12633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _09773_/X _09775_/X _09777_/X _09779_/X _09605_/X vssd1 vssd1 vccd1 vccd1
+ _09780_/X sky130_fd_sc_hd__a221o_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _19299_/CLK _18978_/D vssd1 vssd1 vccd1 vccd1 _18978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _17929_/A vssd1 vssd1 vccd1 vccd1 _17929_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10952__S0 _09530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14529__S _14535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11742__A _11910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09214_ _09275_/B _09275_/D _09214_/C vssd1 vssd1 vccd1 vccd1 _09215_/B sky130_fd_sc_hd__or3_4
XFILLER_10_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14264__S _14268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11432__S1 _10604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_opt_1_0_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09978_ _10834_/A _09978_/B _09978_/C vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__or3_2
XFILLER_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_133_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11940_ _11940_/A vssd1 vssd1 vccd1 vccd1 _11940_/Y sky130_fd_sc_hd__inv_6
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11871_ _11977_/A vssd1 vssd1 vccd1 vccd1 _11871_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _14844_/C vssd1 vssd1 vccd1 vccd1 _16371_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10822_ _10821_/B _12645_/B vssd1 vssd1 vccd1 vccd1 _10823_/B sky130_fd_sc_hd__and2b_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14590_ _14589_/X _18868_/Q _14590_/S vssd1 vssd1 vccd1 vccd1 _14591_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13262__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09466__B1 _09465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13541_ _18499_/Q _13540_/X _13558_/S vssd1 vssd1 vccd1 vccd1 _13542_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_1_clock clkbuf_1_1_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_10753_ _18806_/Q _19141_/Q _10753_/S vssd1 vssd1 vccd1 vccd1 _10754_/B sky130_fd_sc_hd__mux2_1
XANTENNA__14963__A _14974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10171__S1 _10219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16260_ _16260_/A vssd1 vssd1 vccd1 vccd1 _19524_/D sky130_fd_sc_hd__clkbuf_1
X_13472_ _18495_/Q _13471_/X _13524_/S vssd1 vssd1 vccd1 vccd1 _13473_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ _18583_/Q _18844_/Q _18743_/Q _19078_/Q _10617_/X _10682_/A vssd1 vssd1 vccd1
+ vccd1 _10685_/B sky130_fd_sc_hd__mux4_2
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _15211_/A vssd1 vssd1 vccd1 vccd1 _19133_/D sky130_fd_sc_hd__clkbuf_1
X_12423_ _12470_/C _12422_/Y _12628_/A vssd1 vssd1 vccd1 vccd1 _12423_/Y sky130_fd_sc_hd__o21ai_2
X_16191_ _16191_/A vssd1 vssd1 vccd1 vccd1 _16200_/S sky130_fd_sc_hd__buf_4
XANTENNA__14174__S _14174_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11120__S0 _10999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15142_ _15142_/A vssd1 vssd1 vccd1 vccd1 _19102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12354_ _12573_/S vssd1 vssd1 vccd1 vccd1 _17464_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_127_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17700__A1 _17702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17485__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ _18667_/Q _19162_/Q _11305_/S vssd1 vssd1 vccd1 vccd1 _11305_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13317__A2 _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19950_ _19985_/CLK _19950_/D vssd1 vssd1 vccd1 vccd1 _19950_/Q sky130_fd_sc_hd__dfxtp_2
X_15073_ _15073_/A vssd1 vssd1 vccd1 vccd1 _19070_/D sky130_fd_sc_hd__clkbuf_1
X_12285_ _19596_/Q vssd1 vssd1 vccd1 vccd1 _12339_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18901_ _19487_/CLK _18901_/D vssd1 vssd1 vccd1 vccd1 _18901_/Q sky130_fd_sc_hd__dfxtp_1
X_14024_ _18644_/Q _13651_/X _14024_/S vssd1 vssd1 vccd1 vccd1 _14025_/A sky130_fd_sc_hd__mux2_1
X_11236_ _11236_/A _11236_/B vssd1 vssd1 vccd1 vccd1 _11236_/X sky130_fd_sc_hd__and2_1
XFILLER_171_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19881_ _19881_/CLK _19881_/D vssd1 vssd1 vccd1 vccd1 _19881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11879__A2 _09345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17464__A0 _19968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18832_ _19389_/CLK _18832_/D vssd1 vssd1 vccd1 vccd1 _18832_/Q sky130_fd_sc_hd__dfxtp_1
X_11167_ _18797_/Q _19132_/Q _11222_/S vssd1 vssd1 vccd1 vccd1 _11168_/B sky130_fd_sc_hd__mux2_1
XFILLER_132_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10118_ _18598_/Q _18859_/Q _18758_/Q _19093_/Q _10753_/S _10014_/A vssd1 vssd1 vccd1
+ vccd1 _10118_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18763_ _19258_/CLK _18763_/D vssd1 vssd1 vccd1 vccd1 _18763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15975_ _15975_/A vssd1 vssd1 vccd1 vccd1 _15984_/S sky130_fd_sc_hd__buf_4
X_11098_ _19361_/Q _18975_/Q _19425_/Q _18544_/Q _11035_/X _11330_/A vssd1 vssd1 vccd1
+ vccd1 _11099_/B sky130_fd_sc_hd__mux4_1
XFILLER_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15733__S _15757_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17714_ _17711_/X _17712_/X _17887_/S vssd1 vssd1 vccd1 vccd1 _17714_/X sky130_fd_sc_hd__mux2_1
X_10049_ _19382_/Q _18996_/Q _19446_/Q _18565_/Q _11451_/S _10037_/X vssd1 vssd1 vccd1
+ vccd1 _10050_/B sky130_fd_sc_hd__mux4_1
X_14926_ _19005_/Q _14382_/X _14928_/S vssd1 vssd1 vccd1 vccd1 _14927_/A sky130_fd_sc_hd__mux2_1
X_18694_ _19285_/CLK _18694_/D vssd1 vssd1 vccd1 vccd1 _18694_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15778__B1 _16315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17645_ _17626_/X _17633_/Y _17644_/X vssd1 vssd1 vccd1 vccd1 _17645_/X sky130_fd_sc_hd__a21o_1
X_14857_ _14857_/A vssd1 vssd1 vccd1 vccd1 _18974_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12658__A _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11562__A _11562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13808_ _13808_/A vssd1 vssd1 vccd1 vccd1 _18556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14788_ _14810_/A vssd1 vssd1 vccd1 vccd1 _14797_/S sky130_fd_sc_hd__clkbuf_4
X_17576_ _17571_/X _17574_/X _17759_/S vssd1 vssd1 vccd1 vccd1 _17576_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19315_ _19571_/CLK _19315_/D vssd1 vssd1 vccd1 vccd1 _19315_/Q sky130_fd_sc_hd__dfxtp_1
X_16527_ _19616_/Q _16527_/B _16527_/C vssd1 vssd1 vccd1 vccd1 _16528_/C sky130_fd_sc_hd__and3_1
XFILLER_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13739_ _14672_/A vssd1 vssd1 vccd1 vccd1 _13739_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19246_ _19409_/CLK _19246_/D vssd1 vssd1 vccd1 vccd1 _19246_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09967__A _09967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16458_ _18404_/A _16458_/B vssd1 vssd1 vccd1 vccd1 _16459_/A sky130_fd_sc_hd__or2_1
XFILLER_31_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15409_ _14624_/X _19209_/Q _15417_/S vssd1 vssd1 vccd1 vccd1 _15410_/A sky130_fd_sc_hd__mux2_1
X_19177_ _19405_/CLK _19177_/D vssd1 vssd1 vccd1 vccd1 _19177_/Q sky130_fd_sc_hd__dfxtp_1
X_16389_ _13149_/X _19553_/Q _16393_/S vssd1 vssd1 vccd1 vccd1 _16390_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18128_ _19925_/Q _19957_/Q _18136_/S vssd1 vssd1 vccd1 vccd1 _18129_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15908__S _15912_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18059_ _17771_/X _18055_/Y _18058_/Y vssd1 vssd1 vccd1 vccd1 _18059_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_144_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09901_ _09901_/A vssd1 vssd1 vccd1 vccd1 _09902_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10527__C1 _10307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20021_ _20027_/CLK _20021_/D vssd1 vssd1 vccd1 vccd1 _20021_/Q sky130_fd_sc_hd__dfxtp_1
X_09832_ _19509_/Q _18921_/Q _18958_/Q _18532_/Q _09812_/X _09822_/X vssd1 vssd1 vccd1
+ vccd1 _09833_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09393__C1 _12677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15209__A _15209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _18695_/Q _19190_/Q _09763_/S vssd1 vssd1 vccd1 vccd1 _09763_/X sky130_fd_sc_hd__mux2_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13952__A _13998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09694_ _09694_/A vssd1 vssd1 vccd1 vccd1 _09695_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13492__A1 _16347_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12568__A _18347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12287__B _12287_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11255__B1 _12634_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A _10817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18255__A _18255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11102__S0 _11035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14722__S _14724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12070_ _20028_/Q _11901_/A _17394_/B vssd1 vssd1 vccd1 vccd1 _12070_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__10518__C1 _10307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17446__A0 _17914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ _11016_/A _11017_/X _11020_/X _09975_/A vssd1 vssd1 vccd1 vccd1 _11021_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15553__S _15561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15760_ _15760_/A vssd1 vssd1 vccd1 vccd1 _15800_/S sky130_fd_sc_hd__buf_2
XANTENNA__17334__A _18118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _18459_/Q _12966_/X _10240_/A _12969_/X vssd1 vssd1 vccd1 vccd1 _18459_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09551__S _09763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A io_dbus_rdata[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14711_ _18909_/Q _14414_/X _14713_/S vssd1 vssd1 vccd1 vccd1 _14712_/A sky130_fd_sc_hd__mux2_1
X_11923_ _11923_/A _11923_/B vssd1 vssd1 vccd1 vccd1 _11924_/A sky130_fd_sc_hd__and2_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _15689_/X _19329_/Q _15720_/S vssd1 vssd1 vccd1 vccd1 _15692_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _14640_/X _18884_/Q _14654_/S vssd1 vssd1 vccd1 vccd1 _14643_/A sky130_fd_sc_hd__mux2_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17430_ _17642_/B _12553_/A _17450_/S vssd1 vssd1 vccd1 vccd1 _17430_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11854_ _20032_/Q _11854_/B vssd1 vssd1 vccd1 vccd1 _11854_/X sky130_fd_sc_hd__or2_1
XFILLER_73_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _10805_/A _10805_/B vssd1 vssd1 vccd1 vccd1 _10805_/X sky130_fd_sc_hd__or2_1
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14573_ _14573_/A vssd1 vssd1 vccd1 vccd1 _18863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17361_ _17373_/A _17361_/B vssd1 vssd1 vccd1 vccd1 _17362_/A sky130_fd_sc_hd__and2_1
XFILLER_60_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14693__A _14750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ _11785_/A vssd1 vssd1 vccd1 vccd1 _18286_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13801__S _13813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11341__S0 _11161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19100_ _19196_/CLK _19100_/D vssd1 vssd1 vccd1 vccd1 _19100_/Q sky130_fd_sc_hd__dfxtp_1
X_13524_ _18498_/Q _13523_/X _13524_/S vssd1 vssd1 vccd1 vccd1 _13525_/A sky130_fd_sc_hd__mux2_1
X_16312_ _16313_/A _16321_/D vssd1 vssd1 vccd1 vccd1 _16317_/B sky130_fd_sc_hd__nor2_1
X_10736_ _09813_/A _10735_/X _10746_/A vssd1 vssd1 vccd1 vccd1 _10736_/X sky130_fd_sc_hd__a21o_1
X_17292_ _17292_/A vssd1 vssd1 vccd1 vccd1 _19869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19031_ _19063_/CLK _19031_/D vssd1 vssd1 vccd1 vccd1 _19031_/Q sky130_fd_sc_hd__dfxtp_1
X_16243_ _16243_/A vssd1 vssd1 vccd1 vccd1 _19521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13455_ _18494_/Q _13453_/X _13524_/S vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ _10768_/A _10666_/X _10655_/X vssd1 vssd1 vccd1 vccd1 _10667_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12417__S _12562_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10726__A _10727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12406_ _19980_/Q _11421_/A _12528_/S vssd1 vssd1 vccd1 vccd1 _12407_/A sky130_fd_sc_hd__mux2_4
XFILLER_12_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16174_ _19501_/Q _14631_/A _16178_/S vssd1 vssd1 vccd1 vccd1 _16175_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13386_ hold14/A _12891_/X _13385_/X vssd1 vssd1 vccd1 vccd1 _13386_/X sky130_fd_sc_hd__o21a_1
X_10598_ _10322_/A _10588_/Y _10593_/X _10597_/Y _09740_/A vssd1 vssd1 vccd1 vccd1
+ _10598_/X sky130_fd_sc_hd__o311a_2
X_15125_ _14666_/X _19094_/Q _15127_/S vssd1 vssd1 vccd1 vccd1 _15126_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15728__S _15747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 _11704_/A vssd1 vssd1 vccd1 vccd1 io_dbus_st_type[1] sky130_fd_sc_hd__buf_2
XFILLER_127_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12337_ _19598_/Q vssd1 vssd1 vccd1 vccd1 _12340_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14632__S _14638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput119 _12656_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[19] sky130_fd_sc_hd__buf_2
XFILLER_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09726__S _09726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15056_ _15056_/A vssd1 vssd1 vccd1 vccd1 _19063_/D sky130_fd_sc_hd__clkbuf_1
X_19933_ _19938_/CLK _19933_/D vssd1 vssd1 vccd1 vccd1 _19933_/Q sky130_fd_sc_hd__dfxtp_1
X_12268_ _12215_/X _12266_/Y _12316_/C _12218_/X vssd1 vssd1 vccd1 vccd1 _12268_/Y
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__12660__B _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ _18636_/Q _13618_/X _14013_/S vssd1 vssd1 vccd1 vccd1 _14008_/A sky130_fd_sc_hd__mux2_1
X_11219_ _11212_/Y _11214_/Y _11216_/Y _11218_/Y _10994_/X vssd1 vssd1 vccd1 vccd1
+ _11219_/X sky130_fd_sc_hd__o221a_2
X_19864_ _19865_/CLK _19864_/D vssd1 vssd1 vccd1 vccd1 _19864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12199_ _12229_/A _17447_/A vssd1 vssd1 vccd1 vccd1 _12201_/A sky130_fd_sc_hd__nand2_1
XFILLER_95_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput90 _12509_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[27] sky130_fd_sc_hd__buf_2
X_18815_ _19504_/CLK _18815_/D vssd1 vssd1 vccd1 vccd1 _18815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19795_ _19803_/CLK _19795_/D vssd1 vssd1 vccd1 vccd1 _19795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18746_ _19305_/CLK _18746_/D vssd1 vssd1 vccd1 vccd1 _18746_/Q sky130_fd_sc_hd__dfxtp_1
X_15958_ _19405_/Q _15254_/X _15962_/S vssd1 vssd1 vccd1 vccd1 _15959_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13474__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ _14666_/X _18998_/Q _14911_/S vssd1 vssd1 vccd1 vccd1 _14910_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13491__B _19953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18677_ _19268_/CLK _18677_/D vssd1 vssd1 vccd1 vccd1 _18677_/Q sky130_fd_sc_hd__dfxtp_1
X_15889_ _15889_/A vssd1 vssd1 vccd1 vccd1 _19374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10383__S1 _09841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17628_ _17628_/A vssd1 vssd1 vccd1 vccd1 _17628_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13226__A1 _12851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17559_ _17798_/A vssd1 vssd1 vccd1 vccd1 _17560_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13711__S _13715_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__S0 _11026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19229_ _19391_/CLK _19229_/D vssd1 vssd1 vccd1 vccd1 _19229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10748__C1 _09603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14542__S _14546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09905__A1 _09822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09815_ _09815_/A vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__buf_2
X_20004_ _20048_/CLK _20004_/D vssd1 vssd1 vccd1 vccd1 _20004_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input3_A io_dbus_rdata[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09746_ _09746_/A vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_171_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19540_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09677_ _11141_/A vssd1 vssd1 vccd1 vccd1 _10051_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10374__S1 _09520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13217__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_186_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19881_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10126__S1 _10718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11779__A1 _19819_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11930__A _17772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11570_ _11570_/A _11570_/B _11570_/C vssd1 vssd1 vccd1 vccd1 _11570_/Y sky130_fd_sc_hd__nand3_2
XFILLER_35_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12745__B _18281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ _10521_/A _10521_/B vssd1 vssd1 vccd1 vccd1 _10521_/X sky130_fd_sc_hd__or2_1
XFILLER_155_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09819__S1 _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _18481_/Q _13239_/X _13278_/S vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10452_ _10490_/A _10452_/B vssd1 vssd1 vccd1 vccd1 _10452_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13857__A _13913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ _13214_/C _13299_/C _13171_/C vssd1 vssd1 vccd1 vccd1 _13171_/X sky130_fd_sc_hd__and3b_1
XFILLER_163_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10383_ _19471_/Q _19309_/Q _18718_/Q _18488_/Q _10382_/X _09841_/A vssd1 vssd1 vccd1
+ vccd1 _10384_/B sky130_fd_sc_hd__mux4_1
XFILLER_124_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12122_ _12584_/B vssd1 vssd1 vccd1 vccd1 _12122_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input59_A io_ibus_inst[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_124_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19200_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16930_ _19739_/Q _19738_/Q _19737_/Q _16930_/D vssd1 vssd1 vccd1 vccd1 _16965_/C
+ sky130_fd_sc_hd__and4_1
X_12053_ _12052_/Y _12021_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12053_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_81_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11004_ _18801_/Q _19136_/Q _11004_/S vssd1 vssd1 vccd1 vccd1 _11004_/X sky130_fd_sc_hd__mux2_1
X_16861_ _16865_/A _16870_/D _16860_/X vssd1 vssd1 vccd1 vccd1 _16861_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18600_ _19063_/CLK _18600_/D vssd1 vssd1 vccd1 vccd1 _18600_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_139_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19484_/CLK sky130_fd_sc_hd__clkbuf_16
X_15812_ _18463_/Q _13467_/X _15811_/Y _15700_/X vssd1 vssd1 vccd1 vccd1 _15812_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19580_ _19592_/CLK _19580_/D vssd1 vssd1 vccd1 vccd1 _19580_/Q sky130_fd_sc_hd__dfxtp_1
X_16792_ _19702_/Q _16795_/C vssd1 vssd1 vccd1 vccd1 _16793_/B sky130_fd_sc_hd__and2_1
XFILLER_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18531_ _19377_/CLK _18531_/D vssd1 vssd1 vccd1 vccd1 _18531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15743_ _18451_/Q _13269_/X _15742_/Y _13580_/X vssd1 vssd1 vccd1 vccd1 _15743_/X
+ sky130_fd_sc_hd__o211a_1
X_12955_ _18447_/Q _12951_/X _10821_/B _12954_/X vssd1 vssd1 vccd1 vccd1 _18447_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18395__B2 _18394_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11906_ _11933_/A _11933_/B _11861_/A vssd1 vssd1 vccd1 vccd1 _11907_/B sky130_fd_sc_hd__a21o_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _19952_/CLK _18462_/D vssd1 vssd1 vccd1 vccd1 _18462_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13208__A1 _19748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15674_/A vssd1 vssd1 vccd1 vccd1 _19326_/D sky130_fd_sc_hd__clkbuf_1
X_12886_ _13527_/B vssd1 vssd1 vccd1 vccd1 _12887_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17792_/B _12432_/A _17419_/A vssd1 vssd1 vccd1 vccd1 _17413_/X sky130_fd_sc_hd__mux2_1
X_14625_ _14657_/A vssd1 vssd1 vccd1 vccd1 _14638_/S sky130_fd_sc_hd__buf_2
X_11837_ _11837_/A _11952_/B vssd1 vssd1 vccd1 vccd1 _11950_/B sky130_fd_sc_hd__nor2_2
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18393_ _18396_/A _18393_/B vssd1 vssd1 vccd1 vccd1 _20033_/D sky130_fd_sc_hd__nor2_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11314__S0 _10999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12967__B1 _10459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _14556_/A vssd1 vssd1 vccd1 vccd1 _18855_/D sky130_fd_sc_hd__clkbuf_1
X_17344_ _17355_/A _17344_/B vssd1 vssd1 vccd1 vccd1 _17345_/A sky130_fd_sc_hd__and2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11768_ _11920_/A vssd1 vssd1 vccd1 vccd1 _12066_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12655__B _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ _18647_/Q _19238_/Q _19400_/Q _18615_/Q _10649_/X _10754_/A vssd1 vssd1 vccd1
+ vccd1 _10720_/B sky130_fd_sc_hd__mux4_1
X_13507_ _18497_/Q _13506_/X _13524_/S vssd1 vssd1 vccd1 vccd1 _13508_/A sky130_fd_sc_hd__mux2_1
X_17275_ _17275_/A vssd1 vssd1 vccd1 vccd1 _19861_/D sky130_fd_sc_hd__clkbuf_1
X_14487_ input47/X vssd1 vssd1 vccd1 vccd1 _14487_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_174_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10456__A _19911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11699_ _11699_/A _11699_/B vssd1 vssd1 vccd1 vccd1 _11699_/X sky130_fd_sc_hd__and2_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19014_ _19495_/CLK _19014_/D vssd1 vssd1 vccd1 vccd1 _19014_/Q sky130_fd_sc_hd__dfxtp_1
X_16226_ _16226_/A vssd1 vssd1 vccd1 vccd1 _16262_/S sky130_fd_sc_hd__clkbuf_2
X_13438_ _19949_/Q _19950_/Q _13438_/C vssd1 vssd1 vccd1 vccd1 _13460_/B sky130_fd_sc_hd__and3_1
XFILLER_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13767__A _14592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16157_ _16157_/A vssd1 vssd1 vccd1 vccd1 _19493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13369_ _16922_/B _13341_/X _13342_/X _19694_/Q _13368_/X vssd1 vssd1 vccd1 vccd1
+ _13369_/X sky130_fd_sc_hd__a221o_2
XFILLER_155_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12671__A _12671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15108_ _14640_/X _19086_/Q _15116_/S vssd1 vssd1 vccd1 vccd1 _15109_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16330__A0 _19537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16088_ _16088_/A vssd1 vssd1 vccd1 vccd1 _19462_/D sky130_fd_sc_hd__clkbuf_1
X_15039_ _15039_/A vssd1 vssd1 vccd1 vccd1 _19055_/D sky130_fd_sc_hd__clkbuf_1
X_19916_ _19919_/CLK _19916_/D vssd1 vssd1 vccd1 vccd1 _19916_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19847_ _19876_/CLK _19847_/D vssd1 vssd1 vccd1 vccd1 _19847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17830__A0 _17832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ _09600_/A vssd1 vssd1 vccd1 vccd1 _09601_/A sky130_fd_sc_hd__buf_2
XFILLER_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19778_ _19877_/CLK _19778_/D vssd1 vssd1 vccd1 vccd1 _19778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09531_ _09967_/A vssd1 vssd1 vccd1 vccd1 _09532_/A sky130_fd_sc_hd__buf_2
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18729_ _19482_/CLK _18729_/D vssd1 vssd1 vccd1 vccd1 _18729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15921__S _15929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18386__B2 _18385_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09462_ _12747_/A _17322_/A vssd1 vssd1 vccd1 vccd1 _12933_/A sky130_fd_sc_hd__nand2_4
XFILLER_58_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10681__A1 _09814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09393_ _13136_/D _12693_/C _12914_/B _12677_/A _12697_/A vssd1 vssd1 vccd1 vccd1
+ _09401_/B sky130_fd_sc_hd__a2111oi_1
XFILLER_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15222__A _15222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12186__A1 _16226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19565_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13677__A _13719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10292__S0 _10465_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15892__A _15903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19985_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_120_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09729_ _18602_/Q _18863_/Q _18762_/Q _19097_/Q _09655_/X _09727_/A vssd1 vssd1 vccd1
+ vccd1 _09729_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ _12853_/A vssd1 vssd1 vccd1 vccd1 _13577_/A sky130_fd_sc_hd__buf_2
XFILLER_28_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12671_/A vssd1 vssd1 vccd1 vccd1 _12671_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17331__B _17331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12756__A _12756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16228__A _16299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14410_ _14410_/A vssd1 vssd1 vccd1 vccd1 _18806_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11660__A _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12949__B1 _11352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11622_ _11622_/A vssd1 vssd1 vccd1 vccd1 _17392_/B sky130_fd_sc_hd__inv_2
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15390_/A vssd1 vssd1 vccd1 vccd1 _19200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14341_ _18782_/Q _13693_/X _14341_/S vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _11556_/A _11558_/A _11556_/C _10364_/A vssd1 vssd1 vccd1 vccd1 _11553_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10504_ _10500_/A _10501_/X _10503_/X vssd1 vssd1 vccd1 vccd1 _10504_/Y sky130_fd_sc_hd__o21ai_1
X_17060_ _17062_/A _17062_/C _17059_/X vssd1 vssd1 vccd1 vccd1 _17060_/Y sky130_fd_sc_hd__a21oi_1
X_14272_ _14272_/A vssd1 vssd1 vccd1 vccd1 _18751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11484_ _09957_/A _11483_/X _11478_/A vssd1 vssd1 vccd1 vccd1 _11484_/X sky130_fd_sc_hd__a21o_1
X_16011_ _16011_/A vssd1 vssd1 vccd1 vccd1 _19428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13223_ _19936_/Q vssd1 vssd1 vccd1 vccd1 _16265_/A sky130_fd_sc_hd__clkbuf_2
X_10435_ _19116_/Q _18882_/Q _19564_/Q _19212_/Q _10325_/X _10497_/A vssd1 vssd1 vccd1
+ vccd1 _10436_/B sky130_fd_sc_hd__mux4_1
XFILLER_137_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12491__A _19843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13154_ _13154_/A vssd1 vssd1 vccd1 vccd1 _13154_/Y sky130_fd_sc_hd__inv_2
X_10366_ _19117_/Q _18883_/Q _19565_/Q _19213_/Q _09505_/A _10312_/X vssd1 vssd1 vccd1
+ vccd1 _10366_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output165_A _12590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12194_/A _12195_/B vssd1 vssd1 vccd1 vccd1 _12106_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _19897_/Q _15679_/B _13430_/S vssd1 vssd1 vccd1 vccd1 _13085_/X sky130_fd_sc_hd__mux2_1
X_17962_ _18078_/S _17963_/B _17961_/X _17723_/A vssd1 vssd1 vccd1 vccd1 _17965_/B
+ sky130_fd_sc_hd__o211a_1
X_10297_ _10571_/A vssd1 vssd1 vccd1 vccd1 _10478_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19701_ _19737_/CLK _19701_/D vssd1 vssd1 vccd1 vccd1 _19701_/Q sky130_fd_sc_hd__dfxtp_1
X_16913_ _16925_/B _16918_/D _16912_/X vssd1 vssd1 vccd1 vccd1 _19735_/D sky130_fd_sc_hd__o21ba_1
X_12036_ _12026_/X _12030_/X _12031_/X _12035_/Y vssd1 vssd1 vccd1 vccd1 _12037_/B
+ sky130_fd_sc_hd__a31o_1
X_17893_ _17893_/A vssd1 vssd1 vccd1 vccd1 _19905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19632_ _19637_/CLK _19632_/D vssd1 vssd1 vccd1 vccd1 _19632_/Q sky130_fd_sc_hd__dfxtp_1
X_16844_ _16864_/C _16848_/C _16848_/D vssd1 vssd1 vccd1 vccd1 _16845_/B sky130_fd_sc_hd__and3_1
XFILLER_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19563_ _19563_/CLK _19563_/D vssd1 vssd1 vccd1 vccd1 _19563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16775_ _16775_/A _16781_/C vssd1 vssd1 vccd1 vccd1 _16775_/Y sky130_fd_sc_hd__nor2_1
X_13987_ _13987_/A vssd1 vssd1 vccd1 vccd1 _18628_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12101__A1 _12606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10338__S1 _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18368__B2 _18367_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18514_ _19491_/CLK _18514_/D vssd1 vssd1 vccd1 vccd1 _18514_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ _19903_/Q _15724_/X _15757_/S vssd1 vssd1 vccd1 vccd1 _15726_/X sky130_fd_sc_hd__mux2_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19494_ _19559_/CLK _19494_/D vssd1 vssd1 vccd1 vccd1 _19494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12938_ _18439_/Q _09464_/X _11348_/A _12947_/A _12937_/X vssd1 vssd1 vccd1 vccd1
+ _18439_/D sky130_fd_sc_hd__a221o_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18445_ _19938_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__14357__S _14363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ _14672_/X _19320_/Q _15659_/S vssd1 vssd1 vccd1 vccd1 _15658_/A sky130_fd_sc_hd__mux2_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12666__A _12669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ _19622_/Q _12861_/X _12868_/X vssd1 vssd1 vccd1 vccd1 _12869_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14608_ _14608_/A vssd1 vssd1 vccd1 vccd1 _14608_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18376_ _18288_/A _18373_/X _18374_/X _18375_/Y vssd1 vssd1 vccd1 vccd1 _18377_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15588_ _15588_/A vssd1 vssd1 vccd1 vccd1 _19289_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17327_ _17327_/A _17327_/B vssd1 vssd1 vccd1 vccd1 _17327_/Y sky130_fd_sc_hd__nor2_1
X_14539_ _14539_/A vssd1 vssd1 vccd1 vccd1 _18847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09975__A _09975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17258_ _17160_/Y _19854_/Q _17258_/S vssd1 vssd1 vccd1 vccd1 _17259_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15696__B _17166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16209_ _18198_/A _16315_/C vssd1 vssd1 vccd1 vccd1 _16299_/A sky130_fd_sc_hd__nor2_2
XFILLER_128_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14092__S _14098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17189_ _19830_/Q _17195_/B vssd1 vssd1 vccd1 vccd1 _17189_/X sky130_fd_sc_hd__or2_1
XANTENNA__10914__A _11026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15916__S _15916_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16601__A _16631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15651__S _15655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ _09514_/A vssd1 vssd1 vccd1 vccd1 _09515_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_140_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _20031_/Q _20030_/Q _20029_/Q _11639_/B vssd1 vssd1 vccd1 vccd1 _11789_/C
+ sky130_fd_sc_hd__or4_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11851__B1 _10065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09376_ _12689_/B _16809_/A _12804_/A vssd1 vssd1 vccd1 vccd1 _12989_/A sky130_fd_sc_hd__nor3_4
XFILLER_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10501__S1 _10397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12159__A1 _12026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ _09868_/A _10217_/Y _10219_/Y _09936_/A vssd1 vssd1 vccd1 vccd1 _10220_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _10151_/A vssd1 vssd1 vccd1 vccd1 _10196_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17607__A _17607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10082_ _10082_/A vssd1 vssd1 vccd1 vccd1 _10083_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13910_ _13910_/A vssd1 vssd1 vccd1 vccd1 _18594_/D sky130_fd_sc_hd__clkbuf_1
X_14890_ _14890_/A vssd1 vssd1 vccd1 vccd1 _18989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13841_ _14666_/A vssd1 vssd1 vccd1 vccd1 _13841_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15561__S _15561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16560_ _19626_/Q _16558_/B _16559_/Y vssd1 vssd1 vccd1 vccd1 _19626_/D sky130_fd_sc_hd__o21a_1
XFILLER_56_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13772_ _13771_/X _18545_/Q _13781_/S vssd1 vssd1 vccd1 vccd1 _13773_/A sky130_fd_sc_hd__mux2_1
X_10984_ _19363_/Q _18977_/Q _19427_/Q _18546_/Q _10018_/A _11225_/A vssd1 vssd1 vccd1
+ vccd1 _10985_/B sky130_fd_sc_hd__mux4_1
XFILLER_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15511_ _19255_/Q _15292_/X _15511_/S vssd1 vssd1 vccd1 vccd1 _15512_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12723_ _12723_/A vssd1 vssd1 vccd1 vccd1 _12723_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14177__S _14185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16491_ _19606_/Q _16487_/X _12543_/Y _12546_/Y _12749_/X vssd1 vssd1 vccd1 vccd1
+ _19606_/D sky130_fd_sc_hd__o221a_1
XFILLER_43_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18230_ _18230_/A vssd1 vssd1 vccd1 vccd1 _19970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12654_ _12657_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _12654_/Y sky130_fd_sc_hd__nor2_2
X_15442_ _15442_/A vssd1 vssd1 vccd1 vccd1 _19224_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17488__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11605_ _11911_/A vssd1 vssd1 vccd1 vccd1 _19323_/D sky130_fd_sc_hd__clkinv_2
XFILLER_8_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18161_ _18183_/A vssd1 vssd1 vccd1 vccd1 _18170_/S sky130_fd_sc_hd__clkbuf_2
X_15373_ _15373_/A _15373_/B _15373_/C vssd1 vssd1 vccd1 vccd1 _15430_/A sky130_fd_sc_hd__or3_4
X_12585_ _12208_/X _12583_/X _12584_/X _12212_/X vssd1 vssd1 vccd1 vccd1 _12585_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14905__S _14911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_128_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17112_ _17112_/A _19800_/Q _17112_/C vssd1 vssd1 vccd1 vccd1 _17114_/B sky130_fd_sc_hd__and3_1
X_14324_ _18774_/Q _13660_/X _14330_/S vssd1 vssd1 vccd1 vccd1 _14325_/A sky130_fd_sc_hd__mux2_1
X_11536_ _11536_/A _11536_/B vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__nand2_1
X_18092_ _17785_/X _18089_/X _18091_/Y _17705_/A vssd1 vssd1 vccd1 vccd1 _18092_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12933__B _12937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14255_ _13793_/X _18744_/Q _14257_/S vssd1 vssd1 vccd1 vccd1 _14256_/A sky130_fd_sc_hd__mux2_1
X_17043_ _17044_/A _17044_/B _17042_/Y vssd1 vssd1 vccd1 vccd1 _19775_/D sky130_fd_sc_hd__o21a_1
X_11467_ _11460_/Y _11462_/Y _11464_/Y _11466_/Y _09717_/A vssd1 vssd1 vccd1 vccd1
+ _11467_/X sky130_fd_sc_hd__o221a_1
XANTENNA__10734__A _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13206_ _19860_/Q _12699_/A _13205_/X _17180_/A vssd1 vssd1 vccd1 vccd1 _13206_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13110__A _13558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10418_ _10368_/A _10417_/X _10478_/A vssd1 vssd1 vccd1 vccd1 _10418_/X sky130_fd_sc_hd__a21o_1
X_14186_ _14186_/A vssd1 vssd1 vccd1 vccd1 _18713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11398_ _18648_/Q _19239_/Q _19401_/Q _18616_/Q _10640_/S _10637_/A vssd1 vssd1 vccd1
+ vccd1 _11399_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _19815_/Q _12677_/A _12804_/Y _19745_/Q _12805_/Y vssd1 vssd1 vccd1 vccd1
+ _13137_/X sky130_fd_sc_hd__a221o_1
X_10349_ _10448_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10349_/Y sky130_fd_sc_hd__nor2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18994_ _19476_/CLK _18994_/D vssd1 vssd1 vccd1 vccd1 _18994_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10581__B1 _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _13060_/X _13067_/X _12988_/A input26/X vssd1 vssd1 vccd1 vccd1 _15209_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_79_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17945_ _17945_/A _17945_/B vssd1 vssd1 vccd1 vccd1 _17945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12019_ _12020_/A _17459_/A vssd1 vssd1 vccd1 vccd1 _12021_/A sky130_fd_sc_hd__nand2_1
X_17876_ _10772_/Y _17861_/X _17875_/X vssd1 vssd1 vccd1 vccd1 _19904_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19615_ _19620_/CLK _19615_/D vssd1 vssd1 vccd1 vccd1 _19615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16827_ _19709_/Q _16823_/B _16826_/Y vssd1 vssd1 vccd1 vccd1 _19709_/D sky130_fd_sc_hd__o21a_1
XFILLER_94_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13780__A _14605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19546_ _19671_/CLK _19546_/D vssd1 vssd1 vccd1 vccd1 _19546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16758_ _16775_/A _16763_/C vssd1 vssd1 vccd1 vccd1 _16758_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10636__A1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15709_ _18445_/Q _15709_/B _15709_/C vssd1 vssd1 vccd1 vccd1 _15709_/X sky130_fd_sc_hd__or3_1
X_19477_ _19481_/CLK _19477_/D vssd1 vssd1 vccd1 vccd1 _19477_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10636__B2 _19907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16689_ _19671_/Q _16689_/B _16689_/C vssd1 vssd1 vccd1 vccd1 _16691_/B sky130_fd_sc_hd__and3_1
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10731__S1 _10609_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09230_ _11601_/A _09238_/A _11730_/C vssd1 vssd1 vccd1 vccd1 _09303_/A sky130_fd_sc_hd__or3_1
X_18428_ _17338_/A _18413_/X _18414_/X _18427_/Y vssd1 vssd1 vccd1 vccd1 _18429_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_22_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12389__B2 _12356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18359_ _18359_/A _18359_/B vssd1 vssd1 vccd1 vccd1 _20023_/D sky130_fd_sc_hd__nor2_1
XFILLER_147_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14815__S _14819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16524__B1 _12908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16315__B _16315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10363__B _12657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09994_ _10730_/A _09991_/X _09993_/X _09976_/X vssd1 vssd1 vccd1 vccd1 _09994_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12313__A1 _19533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18201__A0 _19957_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09428_ _17327_/B _11895_/C vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__and2_1
XFILLER_138_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09359_ _20012_/Q vssd1 vssd1 vccd1 vccd1 _09398_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11052__A1 _10961_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12370_ _19535_/Q _12122_/X _16303_/A vssd1 vssd1 vccd1 vccd1 _12370_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11052__B2 _12638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16515__B1 _12908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11321_ _11271_/A _11320_/X _09470_/A vssd1 vssd1 vccd1 vccd1 _11321_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10554__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14026__A _14072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14040_ _18651_/Q _13681_/X _14046_/S vssd1 vssd1 vccd1 vccd1 _14041_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18268__A0 _19988_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11252_ _11117_/X _11251_/X _10949_/X vssd1 vssd1 vccd1 vccd1 _11252_/X sky130_fd_sc_hd__o21a_1
XFILLER_153_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10203_ _10243_/A _10203_/B vssd1 vssd1 vccd1 vccd1 _10203_/X sky130_fd_sc_hd__or2_1
XANTENNA__10789__S1 _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12552__A1 _11470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14460__S _14466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11183_ _11183_/A _11183_/B vssd1 vssd1 vccd1 vccd1 _11183_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input41_A io_ibus_inst[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _19920_/Q vssd1 vssd1 vccd1 vccd1 _10134_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_122_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15991_ _16047_/A vssd1 vssd1 vccd1 vccd1 _16060_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17730_ _17616_/A _17724_/Y _17729_/Y _17995_/A vssd1 vssd1 vccd1 vccd1 _17730_/X
+ sky130_fd_sc_hd__a211o_1
X_14942_ _19012_/Q _14404_/X _14950_/S vssd1 vssd1 vccd1 vccd1 _14943_/A sky130_fd_sc_hd__mux2_1
X_10065_ _10065_/A vssd1 vssd1 vccd1 vccd1 _10065_/X sky130_fd_sc_hd__buf_2
XFILLER_85_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_54_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17661_ _17601_/X _17660_/X _17800_/S vssd1 vssd1 vccd1 vccd1 _17661_/X sky130_fd_sc_hd__mux2_1
X_14873_ _14873_/A vssd1 vssd1 vccd1 vccd1 _18981_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19400_ _19560_/CLK _19400_/D vssd1 vssd1 vccd1 vccd1 _19400_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output128_A _12666_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13804__S _13813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16612_ _16612_/A vssd1 vssd1 vccd1 vccd1 _16617_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13824_ _13824_/A vssd1 vssd1 vccd1 vccd1 _18561_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12068__B1 _12137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17592_ _17628_/A _17591_/X _17602_/S vssd1 vssd1 vccd1 vccd1 _17592_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19331_ _19881_/CLK _19331_/D vssd1 vssd1 vccd1 vccd1 _19331_/Q sky130_fd_sc_hd__dfxtp_1
X_16543_ _19620_/Q _16539_/C _16542_/Y vssd1 vssd1 vccd1 vccd1 _19620_/D sky130_fd_sc_hd__o21a_1
XFILLER_16_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13755_ _14580_/A vssd1 vssd1 vccd1 vccd1 _13755_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10967_ _10967_/A vssd1 vssd1 vccd1 vccd1 _10967_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13280__A2 _13172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ _12864_/A vssd1 vssd1 vccd1 vccd1 _13245_/A sky130_fd_sc_hd__clkbuf_2
X_19262_ _19391_/CLK _19262_/D vssd1 vssd1 vccd1 vccd1 _19262_/Q sky130_fd_sc_hd__dfxtp_1
X_16474_ _16474_/A vssd1 vssd1 vccd1 vccd1 _16474_/Y sky130_fd_sc_hd__inv_2
X_13686_ _18524_/Q _13685_/X _13694_/S vssd1 vssd1 vccd1 vccd1 _13687_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10898_ _09612_/A _10885_/X _10897_/X _09996_/A _19901_/Q vssd1 vssd1 vccd1 vccd1
+ _11355_/A sky130_fd_sc_hd__a32o_4
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18213_ _18213_/A vssd1 vssd1 vccd1 vccd1 _19962_/D sky130_fd_sc_hd__clkbuf_1
X_15425_ _15425_/A vssd1 vssd1 vccd1 vccd1 _19216_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19193_ _19416_/CLK _19193_/D vssd1 vssd1 vccd1 vccd1 _19193_/Q sky130_fd_sc_hd__dfxtp_1
X_12637_ _12637_/A _12637_/B vssd1 vssd1 vccd1 vccd1 _12637_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14635__S _14638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10477__S0 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18144_ _19932_/Q _19964_/Q _18148_/S vssd1 vssd1 vccd1 vccd1 _18145_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15356_ _19186_/Q _15276_/X _15356_/S vssd1 vssd1 vccd1 vccd1 _15357_/A sky130_fd_sc_hd__mux2_1
X_12568_ _18347_/A _12568_/B vssd1 vssd1 vccd1 vccd1 _12568_/X sky130_fd_sc_hd__or2_1
XFILLER_79_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12663__B _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14307_ _14307_/A vssd1 vssd1 vccd1 vccd1 _18766_/D sky130_fd_sc_hd__clkbuf_1
X_11519_ _11534_/A _11519_/B vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__and2_4
X_18075_ _19919_/Q _18019_/X _18074_/X vssd1 vssd1 vccd1 vccd1 _19919_/D sky130_fd_sc_hd__o21a_1
X_12499_ _18079_/A _12499_/B vssd1 vssd1 vccd1 vccd1 _12503_/A sky130_fd_sc_hd__xor2_1
X_15287_ _19157_/Q _15286_/X hold9/A vssd1 vssd1 vccd1 vccd1 _15288_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17026_ _17046_/A _17026_/B _17026_/C vssd1 vssd1 vccd1 vccd1 _19764_/D sky130_fd_sc_hd__nor3_1
X_14238_ _13767_/X _18736_/Q _14246_/S vssd1 vssd1 vccd1 vccd1 _14239_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11346__A2 _11336_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14169_ _14169_/A vssd1 vssd1 vccd1 vccd1 _18705_/D sky130_fd_sc_hd__clkbuf_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15693__C _15693_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18977_ _19553_/CLK _18977_/D vssd1 vssd1 vccd1 vccd1 _18977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _18054_/A vssd1 vssd1 vccd1 vccd1 _17928_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17859_ _12056_/A _17844_/X _17857_/Y _17858_/X vssd1 vssd1 vccd1 vccd1 _17859_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10952__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15796__A1 _19916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19529_ _19988_/CLK _19529_/D vssd1 vssd1 vccd1 vccd1 _19529_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13015__A _19887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ _09264_/B _09425_/B vssd1 vssd1 vccd1 vccd1 _09214_/C sky130_fd_sc_hd__or2b_1
XFILLER_167_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12782__B2 _19532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13685__A _14631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15376__S _15384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09977_ _09989_/A _09971_/X _09974_/X _09976_/X vssd1 vssd1 vccd1 vccd1 _09978_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10821__B _10821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_opt_5_0_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_clock clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_29_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11870_ _11912_/B _12088_/B _11870_/C _11870_/D vssd1 vssd1 vccd1 vccd1 _11870_/X
+ sky130_fd_sc_hd__and4b_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10821_ _12645_/B _10821_/B vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__and2b_1
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13262__A2 _13172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10752_ _10752_/A vssd1 vssd1 vccd1 vccd1 _10752_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13540_ _15295_/A vssd1 vssd1 vccd1 vccd1 _13540_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _15283_/A vssd1 vssd1 vccd1 vccd1 _13471_/X sky130_fd_sc_hd__clkbuf_2
X_10683_ _18775_/Q _19046_/Q _19270_/Q _19014_/Q _10608_/X _10682_/X vssd1 vssd1 vccd1
+ vccd1 _10683_/X sky130_fd_sc_hd__mux4_2
X_12422_ _19840_/Q _12399_/X _12421_/X vssd1 vssd1 vccd1 vccd1 _12422_/Y sky130_fd_sc_hd__o21ai_1
X_15210_ _19133_/Q _15209_/X _15213_/S vssd1 vssd1 vccd1 vccd1 _15211_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16190_ _16190_/A vssd1 vssd1 vccd1 vccd1 _19508_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11120__S1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12353_ _18012_/A _12353_/B vssd1 vssd1 vccd1 vccd1 _12358_/A sky130_fd_sc_hd__xnor2_1
X_15141_ _19102_/Q vssd1 vssd1 vccd1 vccd1 _15142_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11304_ _11304_/A _11304_/B vssd1 vssd1 vccd1 vccd1 _11304_/Y sky130_fd_sc_hd__nor2_1
X_15072_ _14589_/X _19070_/Q _15072_/S vssd1 vssd1 vccd1 vccd1 _15073_/A sky130_fd_sc_hd__mux2_1
X_12284_ _12287_/B vssd1 vssd1 vccd1 vccd1 _12284_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18900_ _19488_/CLK _18900_/D vssd1 vssd1 vccd1 vccd1 _18900_/Q sky130_fd_sc_hd__dfxtp_1
X_14023_ _14023_/A vssd1 vssd1 vccd1 vccd1 _18643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13595__A _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11235_ _18798_/Q _19133_/Q _11306_/S vssd1 vssd1 vccd1 vccd1 _11236_/B sky130_fd_sc_hd__mux2_1
XANTENNA__14190__S _14196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19880_ _19881_/CLK _19880_/D vssd1 vssd1 vccd1 vccd1 _19880_/Q sky130_fd_sc_hd__dfxtp_1
X_18831_ _19666_/CLK _18831_/D vssd1 vssd1 vccd1 vccd1 _18831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17464__A1 _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10631__S0 _10678_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11166_ _11166_/A vssd1 vssd1 vccd1 vccd1 _11166_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10117_ _10847_/S vssd1 vssd1 vccd1 vccd1 _10753_/S sky130_fd_sc_hd__buf_4
X_18762_ _19285_/CLK _18762_/D vssd1 vssd1 vccd1 vccd1 _18762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15974_ _15974_/A vssd1 vssd1 vccd1 vccd1 _19412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11097_ _11295_/A vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17216__A1 _15784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17713_ _17741_/S vssd1 vssd1 vccd1 vccd1 _17887_/S sky130_fd_sc_hd__clkbuf_2
X_10048_ _10048_/A vssd1 vssd1 vccd1 vccd1 _11451_/S sky130_fd_sc_hd__buf_4
X_14925_ _14925_/A vssd1 vssd1 vccd1 vccd1 _19004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18693_ _19510_/CLK _18693_/D vssd1 vssd1 vccd1 vccd1 _18693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17644_ _17634_/X _17640_/X _17643_/Y _17940_/A vssd1 vssd1 vccd1 vccd1 _17644_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__15778__A1 _19913_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14856_ _14589_/X _18974_/Q _14856_/S vssd1 vssd1 vccd1 vccd1 _14857_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13807_ _13806_/X _18556_/Q _13813_/S vssd1 vssd1 vccd1 vccd1 _13808_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11562__B _12654_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17575_ _17602_/S vssd1 vssd1 vccd1 vccd1 _17759_/S sky130_fd_sc_hd__clkbuf_2
X_14787_ _14787_/A vssd1 vssd1 vccd1 vccd1 _18947_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10459__A _10459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11999_ _11968_/A _17412_/A _11998_/X vssd1 vssd1 vccd1 vccd1 _11999_/X sky130_fd_sc_hd__o21a_1
X_19314_ _19314_/CLK _19314_/D vssd1 vssd1 vccd1 vccd1 _19314_/Q sky130_fd_sc_hd__dfxtp_1
X_16526_ _16527_/B _16527_/C _19616_/Q vssd1 vssd1 vccd1 vccd1 _16528_/B sky130_fd_sc_hd__a21oi_1
XFILLER_90_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13738_ _15295_/A vssd1 vssd1 vccd1 vccd1 _14672_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19245_ _19503_/CLK _19245_/D vssd1 vssd1 vccd1 vccd1 _19245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16457_ _11923_/A _11923_/B _16455_/X vssd1 vssd1 vccd1 vccd1 _19583_/D sky130_fd_sc_hd__a21o_1
X_13669_ _18520_/Q _13668_/X _13673_/S vssd1 vssd1 vccd1 vccd1 _13670_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14365__S _14367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15408_ _15430_/A vssd1 vssd1 vccd1 vccd1 _15417_/S sky130_fd_sc_hd__buf_2
X_19176_ _19401_/CLK _19176_/D vssd1 vssd1 vccd1 vccd1 _19176_/Q sky130_fd_sc_hd__dfxtp_1
X_16388_ _16388_/A vssd1 vssd1 vccd1 vccd1 _19552_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18127_ _18127_/A vssd1 vssd1 vccd1 vccd1 _18136_/S sky130_fd_sc_hd__clkbuf_2
X_15339_ _19178_/Q _15251_/X _15345_/S vssd1 vssd1 vccd1 vccd1 _15340_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18361__A input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09983__A _09983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18058_ _18058_/A _18058_/B vssd1 vssd1 vccd1 vccd1 _18058_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _19122_/Q _18888_/Q _19570_/Q _19218_/Q _10197_/S _09899_/X vssd1 vssd1 vccd1
+ vccd1 _09900_/X sky130_fd_sc_hd__mux4_1
X_17009_ _19760_/Q vssd1 vssd1 vccd1 vccd1 _17016_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_99_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20020_ _20020_/CLK _20020_/D vssd1 vssd1 vccd1 vccd1 _20020_/Q sky130_fd_sc_hd__dfxtp_1
X_09831_ _10207_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _09831_/X sky130_fd_sc_hd__or2_1
XFILLER_86_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _09762_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09762_/X sky130_fd_sc_hd__and2_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _09693_/A vssd1 vssd1 vccd1 vccd1 _09694_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15225__A _15225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__B1 _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14275__S _14279_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12584__A _19544_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11007__B2 _11014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11102__S1 _11168_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10766__B1 _10056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18271__A _18352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10861__S0 _10777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13619__S _13631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17446__A1 _17960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _11125_/A _11020_/B vssd1 vssd1 vccd1 vccd1 _11020_/X sky130_fd_sc_hd__or2_1
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _18458_/Q _12966_/X _11418_/A _12969_/X vssd1 vssd1 vccd1 vccd1 _18458_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12759__A _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _14710_/A vssd1 vssd1 vccd1 vccd1 _18908_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11663__A _20028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11890_/X _11914_/X _11916_/X _11921_/Y vssd1 vssd1 vccd1 vccd1 _11923_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_85_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _15844_/S vssd1 vssd1 vccd1 vccd1 _15720_/S sky130_fd_sc_hd__buf_2
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _14657_/A vssd1 vssd1 vccd1 vccd1 _14654_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _18333_/A _18321_/A _11853_/S vssd1 vssd1 vccd1 vccd1 _11853_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14974__A _14974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _19462_/Q _19300_/Q _18709_/Q _18479_/Q _10073_/X _10609_/A vssd1 vssd1 vccd1
+ vccd1 _10805_/B sky130_fd_sc_hd__mux4_2
XFILLER_26_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17360_ _19887_/Q _17358_/X _17359_/X vssd1 vssd1 vccd1 vccd1 _17361_/B sky130_fd_sc_hd__a21bo_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14572_ _13850_/X _18863_/Q _14572_/S vssd1 vssd1 vccd1 vccd1 _14573_/A sky130_fd_sc_hd__mux2_1
X_11784_ _19516_/Q _11782_/X _13591_/A vssd1 vssd1 vccd1 vccd1 _11784_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11341__S1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16311_ _19533_/Q _16300_/X _16309_/Y _16310_/X vssd1 vssd1 vccd1 vccd1 _19533_/D
+ sky130_fd_sc_hd__o22a_1
X_13523_ _15292_/A vssd1 vssd1 vccd1 vccd1 _13523_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14185__S _14185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10735_ _18806_/Q _19141_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _10735_/X sky130_fd_sc_hd__mux2_1
X_17291_ _15770_/X _19869_/Q _17291_/S vssd1 vssd1 vccd1 vccd1 _17292_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12494__A _12494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19030_ _19286_/CLK _19030_/D vssd1 vssd1 vccd1 vccd1 _19030_/Q sky130_fd_sc_hd__dfxtp_1
X_16242_ _19521_/Q _16241_/X _16252_/S vssd1 vssd1 vccd1 vccd1 _16243_/A sky130_fd_sc_hd__mux2_1
X_13454_ _13454_/A vssd1 vssd1 vccd1 vccd1 _13524_/S sky130_fd_sc_hd__buf_4
X_10666_ _18649_/Q _19240_/Q _19402_/Q _18617_/Q _10653_/X _10665_/X vssd1 vssd1 vccd1
+ vccd1 _10666_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10726__B _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ _18033_/B _12405_/B vssd1 vssd1 vccd1 vccd1 _12410_/A sky130_fd_sc_hd__xnor2_1
X_16173_ _16173_/A vssd1 vssd1 vccd1 vccd1 _19500_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10218__S _10218_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13385_ _19759_/Q _12892_/X _13384_/X _12896_/X vssd1 vssd1 vccd1 vccd1 _13385_/X
+ sky130_fd_sc_hd__a211o_1
X_10597_ _10588_/A _10594_/X _10596_/X vssd1 vssd1 vccd1 vccd1 _10597_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__14913__S _14915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15124_ _15124_/A vssd1 vssd1 vccd1 vccd1 _19093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput109 _12631_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[0] sky130_fd_sc_hd__buf_2
XFILLER_127_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10852__S0 _10053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12336_ _12336_/A vssd1 vssd1 vccd1 vccd1 _12336_/Y sky130_fd_sc_hd__inv_6
XFILLER_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14499__B2 _14498_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15055_ _19063_/Q _14465_/X _15055_/S vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12267_ _19834_/Q _19833_/Q _12267_/C vssd1 vssd1 vccd1 vccd1 _12316_/C sky130_fd_sc_hd__and3_2
X_19932_ _19938_/CLK _19932_/D vssd1 vssd1 vccd1 vccd1 _19932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14006_ _14006_/A vssd1 vssd1 vccd1 vccd1 _18635_/D sky130_fd_sc_hd__clkbuf_1
X_11218_ _11153_/A _11217_/X _09703_/A vssd1 vssd1 vccd1 vccd1 _11218_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09308__A _20044_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19863_ _19865_/CLK _19863_/D vssd1 vssd1 vccd1 vccd1 _19863_/Q sky130_fd_sc_hd__dfxtp_1
X_12198_ _19972_/Q _11411_/A _12198_/S vssd1 vssd1 vccd1 vccd1 _17447_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput80 _12284_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[18] sky130_fd_sc_hd__buf_2
Xoutput91 _12538_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[28] sky130_fd_sc_hd__buf_2
XFILLER_96_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18814_ _19053_/CLK _18814_/D vssd1 vssd1 vccd1 vccd1 _18814_/Q sky130_fd_sc_hd__dfxtp_1
X_11149_ _18799_/Q _19134_/Q _11222_/S vssd1 vssd1 vccd1 vccd1 _11149_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17525__A _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19794_ _19794_/CLK _19794_/D vssd1 vssd1 vccd1 vccd1 _19794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18745_ _19560_/CLK _18745_/D vssd1 vssd1 vccd1 vccd1 _18745_/Q sky130_fd_sc_hd__dfxtp_1
X_15957_ _15957_/A vssd1 vssd1 vccd1 vccd1 _19404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12669__A _12669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11573__A _12076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ _14908_/A vssd1 vssd1 vccd1 vccd1 _18997_/D sky130_fd_sc_hd__clkbuf_1
X_18676_ _19204_/CLK _18676_/D vssd1 vssd1 vccd1 vccd1 _18676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15888_ _13331_/X _19374_/Q _15890_/S vssd1 vssd1 vccd1 vccd1 _15889_/A sky130_fd_sc_hd__mux2_1
X_17627_ _17923_/S vssd1 vssd1 vccd1 vccd1 _17627_/X sky130_fd_sc_hd__clkbuf_2
X_14839_ _18319_/A _16315_/A _14825_/X _14838_/Y vssd1 vssd1 vccd1 vccd1 _18406_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17558_ _18019_/A vssd1 vssd1 vccd1 vccd1 _17558_/X sky130_fd_sc_hd__buf_2
XANTENNA__11332__S1 _11179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16509_ _16820_/A vssd1 vssd1 vccd1 vccd1 _17101_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16176__A1 _14634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17489_ _17586_/S vssd1 vssd1 vccd1 vccd1 _17590_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_149_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10917__A _10917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19228_ _19392_/CLK _19228_/D vssd1 vssd1 vccd1 vccd1 _19228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_176_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19159_ _19511_/CLK _19159_/D vssd1 vssd1 vccd1 vccd1 _19159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14823__S _14823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17125__B1 _17101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12851__B _12851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09218__A _19890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_1_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_143_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20003_ _20048_/CLK _20003_/D vssd1 vssd1 vccd1 vccd1 _20003_/Q sky130_fd_sc_hd__dfxtp_1
X_09814_ _09814_/A vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13963__A _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ _09745_/A vssd1 vssd1 vccd1 vccd1 _09746_/A sky130_fd_sc_hd__buf_2
XFILLER_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _10986_/A vssd1 vssd1 vccd1 vccd1 _11141_/A sky130_fd_sc_hd__buf_2
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17170__A _19823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16167__A1 _14621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12440__A3 _12439_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10520_ _19372_/Q _18986_/Q _19436_/Q _18555_/Q _10470_/X _10510_/A vssd1 vssd1 vccd1
+ vccd1 _10521_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12745__C _17245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _18653_/Q _19244_/Q _19406_/Q _18621_/Q _10337_/X _09667_/A vssd1 vssd1 vccd1
+ vccd1 _10452_/B sky130_fd_sc_hd__mux4_1
XFILLER_108_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14733__S _14735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10739__B1 _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ _16248_/A _13170_/B vssd1 vssd1 vccd1 vccd1 _13171_/C sky130_fd_sc_hd__or2_1
X_10382_ _10382_/A vssd1 vssd1 vccd1 vccd1 _10382_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ _11745_/X _12118_/Y _12178_/C _12120_/X vssd1 vssd1 vccd1 vccd1 _12121_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_151_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ _12052_/A vssd1 vssd1 vccd1 vccd1 _12052_/Y sky130_fd_sc_hd__inv_2
X_11003_ _11003_/A vssd1 vssd1 vccd1 vccd1 _11004_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16860_ _16860_/A vssd1 vssd1 vccd1 vccd1 _16860_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15811_ _15811_/A _18463_/Q vssd1 vssd1 vccd1 vccd1 _15811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13592__B _13592_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16791_ _16874_/A _16791_/B _16795_/C vssd1 vssd1 vccd1 vccd1 _19701_/D sky130_fd_sc_hd__nor3_1
XFILLER_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18530_ _19507_/CLK _18530_/D vssd1 vssd1 vccd1 vccd1 _18530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15742_ _15818_/A _18451_/Q vssd1 vssd1 vccd1 vccd1 _15742_/Y sky130_fd_sc_hd__nand2_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12954_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _19985_/CLK _18461_/D vssd1 vssd1 vccd1 vccd1 _18461_/Q sky130_fd_sc_hd__dfxtp_2
X_11905_ _11905_/A _17421_/A vssd1 vssd1 vccd1 vccd1 _11933_/C sky130_fd_sc_hd__xor2_4
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15673_ _15672_/Y _19326_/Q _15684_/S vssd1 vssd1 vccd1 vccd1 _15674_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12893_/A _16678_/A _12829_/X vssd1 vssd1 vccd1 vccd1 _12885_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _17412_/A vssd1 vssd1 vccd1 vccd1 _17792_/B sky130_fd_sc_hd__clkbuf_2
X_14624_ _14624_/A vssd1 vssd1 vccd1 vccd1 _14624_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _13604_/A _11773_/X _11835_/X vssd1 vssd1 vccd1 vccd1 _11843_/B sky130_fd_sc_hd__a21oi_1
X_18392_ _18302_/A _12880_/A _14481_/X _18391_/Y vssd1 vssd1 vccd1 vccd1 _18393_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12967__A1 _18455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11314__S1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _18301_/A _17324_/X _17326_/X _17342_/X _19883_/Q vssd1 vssd1 vccd1 vccd1
+ _17344_/B sky130_fd_sc_hd__a41o_1
X_14555_ _13825_/X _18855_/Q _14557_/S vssd1 vssd1 vccd1 vccd1 _14556_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11767_ _11767_/A vssd1 vssd1 vccd1 vccd1 _11767_/Y sky130_fd_sc_hd__inv_6
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14209__A _14209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13506_ _15289_/A vssd1 vssd1 vccd1 vccd1 _13506_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10718_ _10718_/A vssd1 vssd1 vccd1 vccd1 _10754_/A sky130_fd_sc_hd__clkbuf_4
X_17274_ _12854_/X _19861_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17275_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14486_ _14831_/A vssd1 vssd1 vccd1 vccd1 _14486_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11698_ _20028_/Q _12639_/A vssd1 vssd1 vccd1 vccd1 _11699_/B sky130_fd_sc_hd__or2_1
XFILLER_174_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19013_ _19369_/CLK _19013_/D vssd1 vssd1 vccd1 vccd1 _19013_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15739__S _15757_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16225_ _16232_/A _16232_/C vssd1 vssd1 vccd1 vccd1 _16225_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11078__S0 _10999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13437_ input18/X _13318_/X _13436_/X vssd1 vssd1 vccd1 vccd1 _13437_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10649_ _10700_/S vssd1 vssd1 vccd1 vccd1 _10649_/X sky130_fd_sc_hd__clkbuf_4
X_16156_ _19493_/Q _14605_/A _16156_/S vssd1 vssd1 vccd1 vccd1 _16157_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13368_ _19630_/Q _13204_/X _13367_/X vssd1 vssd1 vccd1 vccd1 _13368_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15107_ _15118_/A vssd1 vssd1 vccd1 vccd1 _15116_/S sky130_fd_sc_hd__buf_2
XFILLER_5_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12319_ _12378_/B _12319_/B vssd1 vssd1 vccd1 vccd1 _12377_/A sky130_fd_sc_hd__nand2_1
X_16087_ _13219_/X _19462_/Q _16095_/S vssd1 vssd1 vccd1 vccd1 _16088_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13299_ _13312_/B _13299_/B _13299_/C vssd1 vssd1 vccd1 vccd1 _13299_/X sky130_fd_sc_hd__and3b_1
XFILLER_142_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15038_ _19055_/Q _14440_/X _15044_/S vssd1 vssd1 vccd1 vccd1 _15039_/A sky130_fd_sc_hd__mux2_1
X_19915_ _19919_/CLK _19915_/D vssd1 vssd1 vccd1 vccd1 _19915_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11155__B1 _09703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15474__S _15478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19846_ _19879_/CLK _19846_/D vssd1 vssd1 vccd1 vccd1 _19846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17830__A1 _17832_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16989_ _16994_/C _16992_/C _16860_/X vssd1 vssd1 vccd1 vccd1 _16989_/Y sky130_fd_sc_hd__a21oi_1
X_19777_ _19877_/CLK _19777_/D vssd1 vssd1 vccd1 vccd1 _19777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11458__A1 _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09530_ _09530_/A vssd1 vssd1 vccd1 vccd1 _09967_/A sky130_fd_sc_hd__clkbuf_4
X_18728_ _19481_/CLK _18728_/D vssd1 vssd1 vccd1 vccd1 _18728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09461_ _14479_/C _12420_/A vssd1 vssd1 vccd1 vccd1 _17322_/A sky130_fd_sc_hd__nor2_4
X_18659_ _19412_/CLK _18659_/D vssd1 vssd1 vccd1 vccd1 _18659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17702__B _17702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09392_ _12700_/A _12700_/B _09392_/C vssd1 vssd1 vccd1 vccd1 _12697_/A sky130_fd_sc_hd__and3_1
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09501__A _11429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15649__S _15655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14553__S _14557_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10816__S0 _11483_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17149__B _17346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17864__S _18109_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10292__S1 _10291_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15384__S _15384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13693__A _14637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18074__A1 _12485_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17821__A1 _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15832__A0 _13519_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09728_ _09727_/A _09725_/Y _09727_/Y _09722_/A vssd1 vssd1 vccd1 vccd1 _09728_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09659_ _09659_/A vssd1 vssd1 vccd1 vccd1 _09660_/A sky130_fd_sc_hd__buf_2
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12670_ _12670_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__and2_2
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11660__B _17346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _17379_/A _17391_/C vssd1 vssd1 vccd1 vccd1 _11621_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10822__A_N _10821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14340_ _14340_/A vssd1 vssd1 vccd1 vccd1 _18781_/D sky130_fd_sc_hd__clkbuf_1
X_11552_ _11552_/A _11554_/A _11552_/C vssd1 vssd1 vccd1 vccd1 _11552_/Y sky130_fd_sc_hd__nand3_1
X_10503_ _10548_/A _10502_/X _10323_/A vssd1 vssd1 vccd1 vccd1 _10503_/X sky130_fd_sc_hd__o21a_1
XANTENNA__15559__S _15561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14271_ _13815_/X _18751_/Q _14279_/S vssd1 vssd1 vccd1 vccd1 _14272_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14463__S _14466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11483_ _18825_/Q _19160_/Q _11483_/S vssd1 vssd1 vccd1 vccd1 _11483_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12772__A _17245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ _13178_/X _19428_/Q _16012_/S vssd1 vssd1 vccd1 vccd1 _16011_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13374__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ _09615_/A _10424_/X _10433_/X _09622_/A _19911_/Q vssd1 vssd1 vccd1 vccd1
+ _10459_/A sky130_fd_sc_hd__a32o_4
X_13222_ _13222_/A vssd1 vssd1 vccd1 vccd1 _18479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10365_ _10365_/A vssd1 vssd1 vccd1 vccd1 _11556_/A sky130_fd_sc_hd__inv_2
X_13153_ _19682_/Q vssd1 vssd1 vccd1 vccd1 _16737_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _12104_/A _17853_/A _12104_/C _17866_/A vssd1 vssd1 vccd1 vccd1 _12195_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13084_ _13163_/A vssd1 vssd1 vccd1 vccd1 _13430_/S sky130_fd_sc_hd__clkbuf_2
X_17961_ _18033_/A _17964_/B _17607_/A _17960_/Y vssd1 vssd1 vccd1 vccd1 _17961_/X
+ sky130_fd_sc_hd__a211o_1
X_10296_ _10296_/A vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output158_A _12448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13807__S _13813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19700_ _19737_/CLK _19700_/D vssd1 vssd1 vccd1 vccd1 _19700_/Q sky130_fd_sc_hd__dfxtp_1
X_16912_ _16925_/B _16925_/C _16915_/D _16875_/X vssd1 vssd1 vccd1 vccd1 _16912_/X
+ sky130_fd_sc_hd__a31o_1
X_12035_ _12855_/A _12033_/Y _12092_/C _11920_/X vssd1 vssd1 vccd1 vccd1 _12035_/Y
+ sky130_fd_sc_hd__o31ai_1
X_17892_ _19905_/Q _17891_/X _18085_/S vssd1 vssd1 vccd1 vccd1 _17893_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16843_ _19713_/Q _16838_/A _16842_/Y vssd1 vssd1 vccd1 vccd1 _19713_/D sky130_fd_sc_hd__o21a_1
X_19631_ _19768_/CLK _19631_/D vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_124_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10896__C1 _09975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15823__A0 _19920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19562_ _19563_/CLK _19562_/D vssd1 vssd1 vccd1 vccd1 _19562_/Q sky130_fd_sc_hd__dfxtp_1
X_16774_ _19696_/Q _16774_/B vssd1 vssd1 vccd1 vccd1 _16781_/C sky130_fd_sc_hd__and2_1
XANTENNA__12012__A _17176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13986_ _18628_/Q _13718_/X _13994_/S vssd1 vssd1 vccd1 vccd1 _13987_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18513_ _19490_/CLK _18513_/D vssd1 vssd1 vccd1 vccd1 _18513_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15725_ _15760_/A vssd1 vssd1 vccd1 vccd1 _15757_/S sky130_fd_sc_hd__buf_2
XFILLER_46_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12937_ _18316_/A _18196_/S _12937_/C vssd1 vssd1 vccd1 vccd1 _12937_/X sky130_fd_sc_hd__and3_1
X_19493_ _19493_/CLK _19493_/D vssd1 vssd1 vccd1 vccd1 _19493_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14638__S _14638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18444_ _19938_/CLK _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_1
X_15656_ _15656_/A vssd1 vssd1 vccd1 vccd1 _19319_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12868_ _19750_/Q _12840_/X _12867_/X _12846_/X vssd1 vssd1 vccd1 vccd1 _12868_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12666__B _12666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14607_/A vssd1 vssd1 vccd1 vccd1 _18873_/D sky130_fd_sc_hd__clkbuf_1
X_18375_ input63/X vssd1 vssd1 vccd1 vccd1 _18375_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_61_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ _11976_/B vssd1 vssd1 vccd1 vccd1 _11819_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15587_ _19289_/Q _15298_/X _15587_/S vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__mux2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12837_/A _17247_/A vssd1 vssd1 vccd1 vccd1 _12799_/Y sky130_fd_sc_hd__nor2_2
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17326_ _09304_/A _09266_/X _11643_/A _12651_/B _17325_/X vssd1 vssd1 vccd1 vccd1
+ _17326_/X sky130_fd_sc_hd__o2111a_1
X_14538_ _13799_/X _18847_/Q _14546_/S vssd1 vssd1 vccd1 vccd1 _14539_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257_ _17257_/A vssd1 vssd1 vccd1 vccd1 _19853_/D sky130_fd_sc_hd__clkbuf_1
X_14469_ _18825_/Q _14468_/X _14472_/S vssd1 vssd1 vccd1 vccd1 _14470_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_49_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16208_ _18932_/Q _13562_/Y _16208_/S vssd1 vssd1 vccd1 vccd1 _16315_/C sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_170_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19542_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17188_ _12874_/X _17182_/X _17187_/X _17185_/X vssd1 vssd1 vccd1 vccd1 _19829_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16139_ _19485_/Q _14580_/A _16145_/S vssd1 vssd1 vccd1 vccd1 _16140_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10274__S1 _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_185_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19852_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19829_ _19831_/CLK _19829_/D vssd1 vssd1 vccd1 vccd1 _19829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11237__S _11237_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13018__A _13454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09513_ _09513_/A vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10103__B2 _19920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__B1 _09752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _18311_/A _20032_/Q vssd1 vssd1 vccd1 vccd1 _11639_/B sky130_fd_sc_hd__or2_1
XANTENNA__11851__A1 _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_123_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19201_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09375_ _09375_/A vssd1 vssd1 vccd1 vccd1 _16809_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13688__A _15257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_138_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19486_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16064__A _16132_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13108__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__A _11001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10150_ _10209_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _10150_/X sky130_fd_sc_hd__or2_1
XANTENNA__13108__B2 _13007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13627__S _13631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15408__A _15430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _11483_/S vssd1 vssd1 vccd1 vccd1 _10081_/X sky130_fd_sc_hd__buf_4
XFILLER_0_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10840__A _10840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13840_ _13840_/A vssd1 vssd1 vccd1 vccd1 _18566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17342__B _17342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13771_ _14596_/A vssd1 vssd1 vccd1 vccd1 _13771_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10983_ _09999_/A _10965_/Y _10972_/X _10982_/Y _09736_/A vssd1 vssd1 vccd1 vccd1
+ _10983_/X sky130_fd_sc_hd__o311a_1
XFILLER_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11671__A _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15510_ _15510_/A vssd1 vssd1 vccd1 vccd1 _19254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12722_ _12776_/A vssd1 vssd1 vccd1 vccd1 _12723_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16490_ _19605_/Q _16487_/X _12514_/X _12518_/X _16482_/X vssd1 vssd1 vccd1 vccd1
+ _19605_/D sky130_fd_sc_hd__o221a_1
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16230__A0 _19519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17769__S _18109_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15441_ _14672_/X _19224_/Q _15443_/S vssd1 vssd1 vccd1 vccd1 _15442_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12653_ _12657_/A _12653_/B vssd1 vssd1 vccd1 vccd1 _12653_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__10287__A _19914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11604_ _11604_/A _11604_/B _11603_/X vssd1 vssd1 vccd1 vccd1 _11911_/A sky130_fd_sc_hd__nor3b_2
X_18160_ _18160_/A vssd1 vssd1 vccd1 vccd1 _19939_/D sky130_fd_sc_hd__clkbuf_1
X_15372_ _15372_/A vssd1 vssd1 vccd1 vccd1 _19193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12584_ _19544_/Q _12584_/B vssd1 vssd1 vccd1 vccd1 _12584_/X sky130_fd_sc_hd__or2_1
X_17111_ _17112_/A _17112_/C _17110_/Y vssd1 vssd1 vccd1 vccd1 _19799_/D sky130_fd_sc_hd__o21a_1
X_14323_ _14323_/A vssd1 vssd1 vccd1 vccd1 _18773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18091_ _17791_/X _18087_/Y _18090_/Y vssd1 vssd1 vccd1 vccd1 _18091_/Y sky130_fd_sc_hd__a21oi_1
X_11535_ _11535_/A vssd1 vssd1 vccd1 vccd1 _11535_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_50_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17042_ _17044_/A _17044_/B _17021_/X vssd1 vssd1 vccd1 vccd1 _17042_/Y sky130_fd_sc_hd__a21oi_1
X_14254_ _14254_/A vssd1 vssd1 vccd1 vccd1 _18743_/D sky130_fd_sc_hd__clkbuf_1
X_11466_ _11460_/A _11465_/X _09707_/A vssd1 vssd1 vccd1 vccd1 _11466_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_109_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13205_ _13205_/A vssd1 vssd1 vccd1 vccd1 _13205_/X sky130_fd_sc_hd__buf_2
X_10417_ _18685_/Q _19180_/Q _10417_/S vssd1 vssd1 vccd1 vccd1 _10417_/X sky130_fd_sc_hd__mux2_1
X_14185_ _13796_/X _18713_/Q _14185_/S vssd1 vssd1 vccd1 vccd1 _14186_/A sky130_fd_sc_hd__mux2_1
X_11397_ _10052_/X _11396_/X _10056_/X vssd1 vssd1 vccd1 vccd1 _11397_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16297__A0 _19531_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13136_ _09394_/A _13136_/B _18326_/A _13136_/D vssd1 vssd1 vccd1 vccd1 _17146_/B
+ sky130_fd_sc_hd__and4b_1
X_10348_ _19376_/Q _18990_/Q _19440_/Q _18559_/Q _09651_/A _09667_/A vssd1 vssd1 vccd1
+ vccd1 _10349_/B sky130_fd_sc_hd__mux4_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _19313_/CLK _18993_/D vssd1 vssd1 vccd1 vccd1 _18993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18038__A1 _17533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11205__S0 _10937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ _10279_/A _10279_/B vssd1 vssd1 vccd1 vccd1 _10279_/Y sky130_fd_sc_hd__nor2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13094_/C _13063_/Y _13065_/X _13066_/X vssd1 vssd1 vccd1 vccd1 _13067_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10750__A _11359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17944_ _19908_/Q _17758_/X _17943_/X vssd1 vssd1 vccd1 vccd1 _19908_/D sky130_fd_sc_hd__o21a_1
XFILLER_79_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12018_ _19966_/Q _10869_/A _12077_/S vssd1 vssd1 vccd1 vccd1 _17459_/A sky130_fd_sc_hd__mux2_2
XFILLER_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17875_ _12084_/A _17966_/B _17870_/X _17874_/Y _11657_/S vssd1 vssd1 vccd1 vccd1
+ _17875_/X sky130_fd_sc_hd__o221a_2
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11057__S _11057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19614_ _19620_/CLK _19614_/D vssd1 vssd1 vccd1 vccd1 _19614_/Q sky130_fd_sc_hd__dfxtp_1
X_16826_ _16845_/A _16863_/C vssd1 vssd1 vccd1 vccd1 _16826_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16757_ _19690_/Q _16757_/B vssd1 vssd1 vccd1 vccd1 _16763_/C sky130_fd_sc_hd__and2_1
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19545_ _19836_/CLK _19545_/D vssd1 vssd1 vccd1 vccd1 _19545_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19566_/CLK sky130_fd_sc_hd__clkbuf_16
X_13969_ _13969_/A vssd1 vssd1 vccd1 vccd1 _18620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12677__A _12677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15708_ _16213_/A vssd1 vssd1 vccd1 vccd1 _15708_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19476_ _19476_/CLK _19476_/D vssd1 vssd1 vccd1 vccd1 _19476_/Q sky130_fd_sc_hd__dfxtp_1
X_16688_ _16689_/B _16689_/C _16687_/Y vssd1 vssd1 vccd1 vccd1 _19670_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_0_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16221__B1 _12492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15639_ _15639_/A vssd1 vssd1 vccd1 vccd1 _19311_/D sky130_fd_sc_hd__clkbuf_1
X_18427_ input55/X vssd1 vssd1 vccd1 vccd1 _18427_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_55_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19906_/CLK sky130_fd_sc_hd__clkbuf_16
X_18358_ _18276_/A _12795_/X _14831_/X _18357_/Y vssd1 vssd1 vccd1 vccd1 _18359_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09885__S0 _10175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17309_ _15822_/X _19877_/Q _17313_/S vssd1 vssd1 vccd1 vccd1 _17310_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18289_ _18289_/A vssd1 vssd1 vccd1 vccd1 _18289_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15927__S _15929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09993_ _11378_/A _09993_/B vssd1 vssd1 vccd1 vccd1 _09993_/X sky130_fd_sc_hd__or2_1
XFILLER_142_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18029__A1 _12391_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15228__A _15228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09226__A _20050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17788__A0 _17792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16460__B1 _16455_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17162__B _17197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12587__A _17240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11491__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ _11690_/D vssd1 vssd1 vccd1 vccd1 _11895_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18274__A _18352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09358_ _16808_/D _09357_/Y _19771_/Q _18345_/A vssd1 vssd1 vccd1 vccd1 _09358_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11052__A2 _12639_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09289_ _19997_/Q vssd1 vssd1 vccd1 vccd1 _14148_/A sky130_fd_sc_hd__buf_4
XANTENNA__13329__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11320_ _19484_/Q _18896_/Q _18933_/Q _18507_/Q _11003_/A _11059_/A vssd1 vssd1 vccd1
+ vccd1 _11320_/X sky130_fd_sc_hd__mux4_2
XFILLER_153_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_clock clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__10554__B _12653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11251_ _18638_/Q _19229_/Q _19391_/Q _18606_/Q _11057_/S _10943_/X vssd1 vssd1 vccd1
+ vccd1 _11251_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10202_ _18593_/Q _18854_/Q _18753_/Q _19088_/Q _09902_/S _09822_/A vssd1 vssd1 vccd1
+ vccd1 _10203_/B sky130_fd_sc_hd__mux4_1
X_11182_ _18637_/Q _19228_/Q _19390_/Q _18605_/Q _10017_/A _10917_/A vssd1 vssd1 vccd1
+ vccd1 _11183_/B sky130_fd_sc_hd__mux4_1
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18428__A1_N _17338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__A0 _19959_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10133_ _10125_/Y _10127_/Y _10130_/Y _10132_/Y _10063_/X vssd1 vssd1 vccd1 vccd1
+ _10133_/X sky130_fd_sc_hd__o221a_2
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15990_ _16371_/D _15990_/B vssd1 vssd1 vccd1 vccd1 _16047_/A sky130_fd_sc_hd__or2_4
XFILLER_0_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10064_ _10050_/Y _10057_/Y _10060_/Y _10062_/Y _10063_/X vssd1 vssd1 vccd1 vccd1
+ _10064_/X sky130_fd_sc_hd__o221a_1
X_14941_ _14987_/S vssd1 vssd1 vccd1 vccd1 _14950_/S sky130_fd_sc_hd__buf_2
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input34_A io_ibus_inst[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11512__B1 _10655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17660_ _17508_/X _17500_/X _17660_/S vssd1 vssd1 vccd1 vccd1 _17660_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17353__A _18273_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14872_ _14612_/X _18981_/Q _14878_/S vssd1 vssd1 vccd1 vccd1 _14873_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16611_ _16629_/A _16611_/B _16611_/C vssd1 vssd1 vccd1 vccd1 _19644_/D sky130_fd_sc_hd__nor3_1
X_13823_ _13822_/X _18561_/Q _13829_/S vssd1 vssd1 vccd1 vccd1 _13824_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17591_ _17589_/X _17590_/X _17674_/S vssd1 vssd1 vccd1 vccd1 _17591_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14188__S _14196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16542_ _16550_/A _16547_/C vssd1 vssd1 vccd1 vccd1 _16542_/Y sky130_fd_sc_hd__nor2_1
X_19330_ _19873_/CLK _19330_/D vssd1 vssd1 vccd1 vccd1 _19330_/Q sky130_fd_sc_hd__dfxtp_1
X_13754_ _13754_/A vssd1 vssd1 vccd1 vccd1 _18539_/D sky130_fd_sc_hd__clkbuf_1
X_10966_ _18674_/Q _19169_/Q _11026_/S vssd1 vssd1 vccd1 vccd1 _10967_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12705_ _18326_/A _15662_/A vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__nor2_2
X_19261_ _19391_/CLK _19261_/D vssd1 vssd1 vccd1 vccd1 _19261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16473_ _12338_/A _16449_/X _12213_/X _12219_/Y _16468_/X vssd1 vssd1 vccd1 vccd1
+ _19593_/D sky130_fd_sc_hd__o221a_1
X_13685_ _14631_/A vssd1 vssd1 vccd1 vccd1 _13685_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09302__C _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10897_ _09473_/A _10887_/X _10889_/X _10896_/X _09601_/A vssd1 vssd1 vccd1 vccd1
+ _10897_/X sky130_fd_sc_hd__a311o_1
XANTENNA__13820__S _13829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18212_ _19962_/Q _19583_/Q _18220_/S vssd1 vssd1 vccd1 vccd1 _18213_/A sky130_fd_sc_hd__mux2_1
X_15424_ _14647_/X _19216_/Q _15428_/S vssd1 vssd1 vccd1 vccd1 _15425_/A sky130_fd_sc_hd__mux2_1
X_19192_ _19418_/CLK _19192_/D vssd1 vssd1 vccd1 vccd1 _19192_/Q sky130_fd_sc_hd__dfxtp_1
X_12636_ _12637_/A _12636_/B vssd1 vssd1 vccd1 vccd1 _12636_/Y sky130_fd_sc_hd__nor2_8
XFILLER_141_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18143_ _18143_/A vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__clkbuf_1
X_15355_ _15355_/A vssd1 vssd1 vccd1 vccd1 _19185_/D sky130_fd_sc_hd__clkbuf_1
X_12567_ _12561_/A _12537_/X _12563_/X _12566_/Y vssd1 vssd1 vccd1 vccd1 _12567_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14306_ _18766_/Q _13626_/X _14308_/S vssd1 vssd1 vccd1 vccd1 _14307_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11518_ _12593_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _11519_/B sky130_fd_sc_hd__nand2_1
X_18074_ _12485_/Y _18007_/X _18073_/X _18028_/X vssd1 vssd1 vccd1 vccd1 _18074_/X
+ sky130_fd_sc_hd__a211o_1
X_15286_ _15286_/A vssd1 vssd1 vccd1 vccd1 _15286_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12498_ _12427_/A _12429_/B _12451_/A _18068_/A _12429_/A vssd1 vssd1 vccd1 vccd1
+ _12499_/B sky130_fd_sc_hd__o41a_1
XFILLER_116_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17025_ _19764_/Q _17027_/C _17025_/C vssd1 vssd1 vccd1 vccd1 _17026_/C sky130_fd_sc_hd__and3_1
XANTENNA__15747__S _15747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14237_ _14294_/S vssd1 vssd1 vccd1 vccd1 _14246_/S sky130_fd_sc_hd__buf_2
XANTENNA__14651__S _14654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11426__S0 _10690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11449_ _18696_/Q _19191_/Q _11449_/S vssd1 vssd1 vccd1 vccd1 _11450_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11346__A3 _11345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17247__B _17247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14168_ _13771_/X _18705_/Q _14174_/S vssd1 vssd1 vccd1 vccd1 _14169_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _19856_/Q _12755_/A _12696_/A _19823_/Q vssd1 vssd1 vccd1 vccd1 _13119_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _14099_/A vssd1 vssd1 vccd1 vccd1 _18676_/D sky130_fd_sc_hd__clkbuf_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _19552_/CLK _18976_/D vssd1 vssd1 vccd1 vccd1 _18976_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _17927_/A vssd1 vssd1 vccd1 vccd1 _19907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17858_ _18127_/A vssd1 vssd1 vccd1 vccd1 _17858_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15245__A1 _15244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16809_ _16809_/A _16809_/B _16809_/C _16809_/D vssd1 vssd1 vccd1 vccd1 _16809_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__14098__S _14098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17789_ _17958_/A vssd1 vssd1 vccd1 vccd1 _18089_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_47_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11267__C1 _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19528_ _19540_/CLK _19528_/D vssd1 vssd1 vccd1 vccd1 _19528_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10165__S0 _09508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13015__B _13748_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19459_ _19553_/CLK _19459_/D vssd1 vssd1 vccd1 vccd1 _19459_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09880__C1 _09741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09212_ _09272_/C vssd1 vssd1 vccd1 vccd1 _09425_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10655__A _10655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15657__S _15659_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09976_ _09976_/A vssd1 vssd1 vccd1 vccd1 _09976_/X sky130_fd_sc_hd__buf_2
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12298__A1 _18321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13905__S _13911_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _09612_/A _10808_/X _10819_/X _09996_/A _19903_/Q vssd1 vssd1 vccd1 vccd1
+ _10821_/B sky130_fd_sc_hd__a32o_4
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18186__A0 _16347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09466__A2 _09419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10751_ _18678_/Q _19173_/Q _10751_/S vssd1 vssd1 vccd1 vccd1 _10752_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13640__S _13652_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13470_ _13324_/X _13457_/X _13461_/Y _13469_/X vssd1 vssd1 vccd1 vccd1 _15283_/A
+ sky130_fd_sc_hd__a22o_2
X_10682_ _10682_/A vssd1 vssd1 vccd1 vccd1 _10682_/X sky130_fd_sc_hd__buf_2
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12421_ _15806_/A vssd1 vssd1 vccd1 vccd1 _12421_/X sky130_fd_sc_hd__buf_2
XANTENNA__17989__A_N _17985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10565__A _10574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14037__A _14059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12773__A2 _12749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ _15140_/A vssd1 vssd1 vccd1 vccd1 _19101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12352_ _17525_/A _18001_/A _12324_/B vssd1 vssd1 vccd1 vccd1 _12353_/B sky130_fd_sc_hd__a21oi_1
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11303_ _19098_/Q _18864_/Q _19546_/Q _19194_/Q _11004_/S _11061_/A vssd1 vssd1 vccd1
+ vccd1 _11304_/B sky130_fd_sc_hd__mux4_1
XFILLER_4_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15071_ _15071_/A vssd1 vssd1 vccd1 vccd1 _19069_/D sky130_fd_sc_hd__clkbuf_1
X_12283_ _12283_/A _12283_/B vssd1 vssd1 vccd1 vccd1 _12287_/B sky130_fd_sc_hd__xnor2_4
XFILLER_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14022_ _18643_/Q _13647_/X _14024_/S vssd1 vssd1 vccd1 vccd1 _14023_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11234_ _19101_/Q _18867_/Q _19549_/Q _19197_/Q _11129_/X _11061_/A vssd1 vssd1 vccd1
+ vccd1 _11234_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18830_ _19671_/CLK _18830_/D vssd1 vssd1 vccd1 vccd1 _18830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ _18669_/Q _19164_/Q _11327_/S vssd1 vssd1 vccd1 vccd1 _11166_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10631__S1 _10604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10116_ _10116_/A vssd1 vssd1 vccd1 vccd1 _10846_/A sky130_fd_sc_hd__buf_2
XANTENNA_output140_A _12644_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15973_ _19412_/Q _15276_/X _15973_/S vssd1 vssd1 vccd1 vccd1 _15974_/A sky130_fd_sc_hd__mux2_1
X_11096_ _11096_/A vssd1 vssd1 vccd1 vccd1 _11295_/A sky130_fd_sc_hd__clkbuf_2
X_18761_ _19299_/CLK _18761_/D vssd1 vssd1 vccd1 vccd1 _18761_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16398__S _16404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17712_ _17456_/X _17491_/X _17799_/S vssd1 vssd1 vccd1 vccd1 _17712_/X sky130_fd_sc_hd__mux2_1
X_10047_ _11495_/S vssd1 vssd1 vccd1 vccd1 _10048_/A sky130_fd_sc_hd__clkbuf_4
X_14924_ _19004_/Q _14379_/X _14928_/S vssd1 vssd1 vccd1 vccd1 _14925_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18692_ _19287_/CLK _18692_/D vssd1 vssd1 vccd1 vccd1 _18692_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10395__S0 _10268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14855_ _14855_/A vssd1 vssd1 vccd1 vccd1 _18973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17643_ _18121_/B _17637_/Y _17642_/Y vssd1 vssd1 vccd1 vccd1 _17643_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13806_ _14631_/A vssd1 vssd1 vccd1 vccd1 _13806_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17574_ _17572_/X _17573_/X _17608_/A vssd1 vssd1 vccd1 vccd1 _17574_/X sky130_fd_sc_hd__mux2_1
X_14786_ _18947_/Q _14417_/X _14786_/S vssd1 vssd1 vccd1 vccd1 _14787_/A sky130_fd_sc_hd__mux2_1
X_11998_ _11932_/A _11969_/A _11968_/A _17412_/A vssd1 vssd1 vccd1 vccd1 _11998_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10459__B _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19313_ _19313_/CLK _19313_/D vssd1 vssd1 vccd1 vccd1 _19313_/Q sky130_fd_sc_hd__dfxtp_1
X_16525_ _16527_/B _16527_/C _16524_/Y vssd1 vssd1 vccd1 vccd1 _19615_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13737_ _13737_/A vssd1 vssd1 vccd1 vccd1 _18536_/D sky130_fd_sc_hd__clkbuf_1
X_10949_ _18968_/Q vssd1 vssd1 vccd1 vccd1 _10949_/X sky130_fd_sc_hd__buf_2
XFILLER_149_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19244_ _19406_/CLK _19244_/D vssd1 vssd1 vccd1 vccd1 _19244_/Q sky130_fd_sc_hd__dfxtp_1
X_16456_ _11892_/A _11892_/B _16455_/X vssd1 vssd1 vccd1 vccd1 _19582_/D sky130_fd_sc_hd__a21o_1
X_13668_ _14618_/A vssd1 vssd1 vccd1 vccd1 _13668_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15407_ _15407_/A vssd1 vssd1 vccd1 vccd1 _19208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19175_ _19572_/CLK _19175_/D vssd1 vssd1 vccd1 vccd1 _19175_/Q sky130_fd_sc_hd__dfxtp_1
X_12619_ _12618_/A _12618_/B _12618_/C vssd1 vssd1 vccd1 vccd1 _12620_/B sky130_fd_sc_hd__a21o_4
XANTENNA__12213__A1 _19529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16387_ _13128_/X _19552_/Q _16393_/S vssd1 vssd1 vccd1 vccd1 _16388_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13599_ _13599_/A vssd1 vssd1 vccd1 vccd1 _18505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18126_ _19924_/Q _17558_/X _18125_/X vssd1 vssd1 vccd1 vccd1 _19924_/D sky130_fd_sc_hd__o21a_1
X_15338_ _15338_/A vssd1 vssd1 vccd1 vccd1 _19177_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12764__A2 _13142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10194__B _12661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18057_ _18055_/Y _18056_/X _18089_/S vssd1 vssd1 vccd1 vccd1 _18057_/X sky130_fd_sc_hd__mux2_1
X_15269_ _15269_/A vssd1 vssd1 vccd1 vccd1 _19151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17008_ _19759_/Q _17004_/C _17007_/Y vssd1 vssd1 vccd1 vccd1 _19759_/D sky130_fd_sc_hd__o21a_1
XFILLER_172_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09830_ _19381_/Q _18995_/Q _19445_/Q _18564_/Q _09812_/X _09822_/X vssd1 vssd1 vccd1
+ vccd1 _09831_/B sky130_fd_sc_hd__mux4_2
XFILLER_112_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _18823_/Q _19158_/Q _09761_/S vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__mux2_1
XFILLER_101_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18959_ _19478_/CLK _18959_/D vssd1 vssd1 vccd1 vccd1 _18959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _10056_/A vssd1 vssd1 vccd1 vccd1 _09693_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_172_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16337__A _19950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15241__A _15241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10766__A1 _11399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13696__A _15263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_97_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17168__A _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10861__S1 _10010_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13468__A0 _19919_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09959_ _11204_/A vssd1 vssd1 vccd1 vccd1 _10955_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12970_ _18457_/Q _12966_/X _10363_/A _12969_/X vssd1 vssd1 vccd1 vccd1 _18457_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10377__S0 _09505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__A _13748_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _12492_/A _11919_/Y _11920_/X vssd1 vssd1 vccd1 vccd1 _11921_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14640_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _20040_/Q vssd1 vssd1 vccd1 vccd1 _18321_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10129__S0 _10702_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _10746_/A _10802_/X _09979_/A vssd1 vssd1 vccd1 vccd1 _10803_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14571_/A vssd1 vssd1 vccd1 vccd1 _18862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14466__S _14466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12775__A _12989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ _12444_/A vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16310_ _12215_/X _15770_/X _16300_/A vssd1 vssd1 vccd1 vccd1 _16310_/X sky130_fd_sc_hd__a21bo_1
XFILLER_14_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13522_ _13060_/X _13509_/X _13513_/Y _13521_/X vssd1 vssd1 vccd1 vccd1 _15292_/A
+ sky130_fd_sc_hd__a22o_4
X_10734_ _10734_/A _10734_/B vssd1 vssd1 vccd1 vccd1 _10734_/X sky130_fd_sc_hd__and2_1
XANTENNA__12994__A2 _13546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17290_ _17290_/A vssd1 vssd1 vccd1 vccd1 _19868_/D sky130_fd_sc_hd__clkbuf_1
X_16241_ _17127_/A _16240_/Y _16262_/S vssd1 vssd1 vccd1 vccd1 _16241_/X sky130_fd_sc_hd__mux2_1
X_13453_ _15279_/A vssd1 vssd1 vccd1 vccd1 _13453_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10665_ _10665_/A vssd1 vssd1 vccd1 vccd1 _10665_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__14990__A _15046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12404_ _17389_/A _12428_/A vssd1 vssd1 vccd1 vccd1 _12405_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12746__A2 _12741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16172_ _19500_/Q _14628_/A _16178_/S vssd1 vssd1 vccd1 vccd1 _16173_/A sky130_fd_sc_hd__mux2_1
X_13384_ _19345_/Q _13154_/A _12704_/X _19535_/Q _13383_/X vssd1 vssd1 vccd1 vccd1
+ _13384_/X sky130_fd_sc_hd__a221o_1
X_10596_ _11464_/A _10595_/X _09707_/A vssd1 vssd1 vccd1 vccd1 _10596_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15123_ _14663_/X _19093_/Q _15127_/S vssd1 vssd1 vccd1 vccd1 _15124_/A sky130_fd_sc_hd__mux2_1
X_12335_ _12335_/A _12335_/B vssd1 vssd1 vccd1 vccd1 _12336_/A sky130_fd_sc_hd__xnor2_2
XFILLER_154_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10852__S1 _10054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15054_ _15054_/A vssd1 vssd1 vccd1 vccd1 _19062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19931_ _19956_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 _19931_/Q sky130_fd_sc_hd__dfxtp_1
X_12266_ _17199_/A _12267_/C _19834_/Q vssd1 vssd1 vccd1 vccd1 _12266_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11706__A0 _20042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14005_ _18635_/Q _13608_/X _14013_/S vssd1 vssd1 vccd1 vccd1 _14006_/A sky130_fd_sc_hd__mux2_1
X_11217_ _19455_/Q _19293_/Q _18702_/Q _18472_/Q _10968_/S _11164_/X vssd1 vssd1 vccd1
+ vccd1 _11217_/X sky130_fd_sc_hd__mux4_1
X_19862_ _19881_/CLK _19862_/D vssd1 vssd1 vccd1 vccd1 _19862_/Q sky130_fd_sc_hd__dfxtp_1
X_12197_ _17933_/B _12197_/B vssd1 vssd1 vccd1 vccd1 _12229_/A sky130_fd_sc_hd__xor2_1
XFILLER_110_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput81 _12309_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[19] sky130_fd_sc_hd__buf_2
Xoutput92 _12559_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[29] sky130_fd_sc_hd__buf_2
X_18813_ _19439_/CLK _18813_/D vssd1 vssd1 vccd1 vccd1 _18813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11148_ _11083_/S _11146_/Y _11147_/Y _10974_/A vssd1 vssd1 vccd1 vccd1 _11148_/X
+ sky130_fd_sc_hd__a211o_1
X_19793_ _19803_/CLK _19793_/D vssd1 vssd1 vccd1 vccd1 _19793_/Q sky130_fd_sc_hd__dfxtp_1
X_18744_ _19572_/CLK _18744_/D vssd1 vssd1 vccd1 vccd1 _18744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15956_ _19404_/Q _15251_/X _15962_/S vssd1 vssd1 vccd1 vccd1 _15957_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11079_ _11317_/A _11079_/B vssd1 vssd1 vccd1 vccd1 _11079_/X sky130_fd_sc_hd__or2_1
XANTENNA__12669__B _12669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ _14663_/X _18997_/Q _14911_/S vssd1 vssd1 vccd1 vccd1 _14908_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11573__B _12647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15887_ _15887_/A vssd1 vssd1 vccd1 vccd1 _19373_/D sky130_fd_sc_hd__clkbuf_1
X_18675_ _19493_/CLK _18675_/D vssd1 vssd1 vccd1 vccd1 _18675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10693__B1 _09475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17626_ _17827_/A vssd1 vssd1 vccd1 vccd1 _17626_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14838_ input43/X vssd1 vssd1 vccd1 vccd1 _14838_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14769_ _18939_/Q _14392_/X _14775_/S vssd1 vssd1 vccd1 vccd1 _14770_/A sky130_fd_sc_hd__mux2_1
X_17557_ _18127_/A vssd1 vssd1 vccd1 vccd1 _18019_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16508_ _16528_/A _16508_/B _16508_/C vssd1 vssd1 vccd1 vccd1 _19610_/D sky130_fd_sc_hd__nor3_1
X_17488_ _12331_/A _12145_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17488_/X sky130_fd_sc_hd__mux2_2
X_19227_ _19389_/CLK _19227_/D vssd1 vssd1 vccd1 vccd1 _19227_/Q sky130_fd_sc_hd__dfxtp_1
X_16439_ _13540_/X _19576_/Q _16441_/S vssd1 vssd1 vccd1 vccd1 _16440_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18372__A _18380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19158_ _19416_/CLK _19158_/D vssd1 vssd1 vccd1 vccd1 _19158_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10748__A1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18109_ _18111_/A _18111_/B _18109_/S vssd1 vssd1 vccd1 vccd1 _18109_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19089_ _19476_/CLK _19089_/D vssd1 vssd1 vccd1 vccd1 _19089_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10933__A _19901_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14405__A _14472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15000__S _15000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20002_ _20048_/CLK _20002_/D vssd1 vssd1 vccd1 vccd1 _20002_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12370__B1 _16303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09813_ _09813_/A vssd1 vssd1 vccd1 vccd1 _09814_/A sky130_fd_sc_hd__buf_6
XFILLER_59_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13455__S _13524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09744_ _09751_/A _09751_/B _09751_/C _09319_/X vssd1 vssd1 vccd1 vccd1 _09745_/A
+ sky130_fd_sc_hd__o31ai_4
XFILLER_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18389__B1 _18374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09675_ _11091_/A vssd1 vssd1 vccd1 vccd1 _10986_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10133__C1 _10063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14286__S _14290_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12595__A _12600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10450_ _10490_/A _10449_/X _09695_/A vssd1 vssd1 vccd1 vccd1 _10450_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10739__A1 _09577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10381_ _18654_/Q _19245_/Q _19407_/Q _18622_/Q _10416_/S _09520_/A vssd1 vssd1 vccd1
+ vccd1 _10381_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ _12120_/A vssd1 vssd1 vccd1 vccd1 _12120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12051_ _12051_/A vssd1 vssd1 vccd1 vccd1 _12055_/A sky130_fd_sc_hd__clkinv_2
XFILLER_81_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ _11002_/A vssd1 vssd1 vccd1 vccd1 _11003_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15810_ _15810_/A vssd1 vssd1 vccd1 vccd1 _19349_/D sky130_fd_sc_hd__clkbuf_1
X_16790_ _19701_/Q _19700_/Q _16790_/C vssd1 vssd1 vccd1 vccd1 _16795_/C sky130_fd_sc_hd__and3_1
XFILLER_133_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15741_ _15741_/A vssd1 vssd1 vccd1 vccd1 _19337_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _18446_/Q _12951_/X _10869_/A _12947_/X vssd1 vssd1 vccd1 vccd1 _18446_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11904_ _19962_/Q _11082_/X _11966_/A vssd1 vssd1 vccd1 vccd1 _17421_/A sky130_fd_sc_hd__mux2_4
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ _19985_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_2
X_15672_ _11187_/Y _16303_/A _13592_/B vssd1 vssd1 vccd1 vccd1 _15672_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_73_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12884_/A vssd1 vssd1 vccd1 vccd1 _16678_/A sky130_fd_sc_hd__buf_4
XFILLER_61_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14623_ _14623_/A vssd1 vssd1 vccd1 vccd1 _18878_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _17772_/B _12455_/A _17460_/S vssd1 vssd1 vccd1 vccd1 _17411_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18391_ input37/X vssd1 vssd1 vccd1 vccd1 _18391_/Y sky130_fd_sc_hd__inv_12
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _12693_/A _12893_/A _11952_/B _11952_/C _11952_/D vssd1 vssd1 vccd1 vccd1
+ _11835_/X sky130_fd_sc_hd__o2111a_1
XANTENNA__14196__S _14196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output103_A _09202_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11613__S _11657_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17342_ _11624_/A _17342_/B _17342_/C _17342_/D vssd1 vssd1 vccd1 vccd1 _17342_/X
+ sky130_fd_sc_hd__and4b_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14554_/A vssd1 vssd1 vccd1 vccd1 _18854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _11766_/A _11766_/B vssd1 vssd1 vccd1 vccd1 _11767_/A sky130_fd_sc_hd__xor2_2
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10522__S0 _10470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _13324_/X _13490_/X _13493_/Y _13504_/X vssd1 vssd1 vccd1 vccd1 _15289_/A
+ sky130_fd_sc_hd__a22o_2
X_10717_ _11399_/A _10716_/X _10056_/X vssd1 vssd1 vccd1 vccd1 _10717_/Y sky130_fd_sc_hd__o21ai_1
X_17273_ _17273_/A vssd1 vssd1 vccd1 vccd1 _19860_/D sky130_fd_sc_hd__clkbuf_1
X_14485_ _18198_/A vssd1 vssd1 vccd1 vccd1 _14485_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14924__S _14928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_120_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11697_ _11704_/A _11697_/B vssd1 vssd1 vccd1 vccd1 _12639_/A sky130_fd_sc_hd__nor2_4
XFILLER_9_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19012_ _19366_/CLK _19012_/D vssd1 vssd1 vccd1 vccd1 _19012_/Q sky130_fd_sc_hd__dfxtp_1
X_16224_ _16224_/A vssd1 vssd1 vccd1 vccd1 _19518_/D sky130_fd_sc_hd__clkbuf_1
X_13436_ _13436_/A vssd1 vssd1 vccd1 vccd1 _13436_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10648_ _10648_/A vssd1 vssd1 vccd1 vccd1 _11448_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11078__S1 _11065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16155_ _16155_/A vssd1 vssd1 vccd1 vccd1 _19492_/D sky130_fd_sc_hd__clkbuf_1
X_13367_ _19758_/Q _12892_/X _13366_/X _12896_/X vssd1 vssd1 vccd1 vccd1 _13367_/X
+ sky130_fd_sc_hd__a211o_1
X_10579_ _10588_/A _10579_/B vssd1 vssd1 vccd1 vccd1 _10579_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14225__A _14281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15669__A1 _09345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15106_ _15106_/A vssd1 vssd1 vccd1 vccd1 _19085_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16866__B1 _18365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12318_ _12339_/C _12115_/X _12313_/X _12317_/Y vssd1 vssd1 vccd1 vccd1 _12318_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_154_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16086_ _16132_/S vssd1 vssd1 vccd1 vccd1 _16095_/S sky130_fd_sc_hd__buf_6
XFILLER_170_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13298_ _16278_/A _13282_/A _13271_/B _19941_/Q vssd1 vssd1 vccd1 vccd1 _13299_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_142_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15037_ _15037_/A vssd1 vssd1 vccd1 vccd1 _19054_/D sky130_fd_sc_hd__clkbuf_1
X_19914_ _19914_/CLK _19914_/D vssd1 vssd1 vccd1 vccd1 _19914_/Q sky130_fd_sc_hd__dfxtp_4
X_12249_ _12243_/X _12248_/Y _16474_/A _11771_/X vssd1 vssd1 vccd1 vccd1 _12249_/X
+ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__11155__A1 _11141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19845_ _19876_/CLK _19845_/D vssd1 vssd1 vccd1 vccd1 _19845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17291__A0 _15770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19776_ _19877_/CLK _19776_/D vssd1 vssd1 vccd1 vccd1 _19776_/Q sky130_fd_sc_hd__dfxtp_1
X_16988_ _19754_/Q vssd1 vssd1 vccd1 vccd1 _16994_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18727_ _19511_/CLK _18727_/D vssd1 vssd1 vccd1 vccd1 _18727_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10115__C1 _10794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15939_ _15939_/A vssd1 vssd1 vccd1 vccd1 _19396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09989__A _09989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09460_ _14477_/A vssd1 vssd1 vccd1 vccd1 _12420_/A sky130_fd_sc_hd__clkbuf_2
X_18658_ _19411_/CLK _18658_/D vssd1 vssd1 vccd1 vccd1 _18658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17609_ _17958_/A vssd1 vssd1 vccd1 vccd1 _18110_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09391_ _18338_/A _09391_/B _12797_/B _12798_/B vssd1 vssd1 vccd1 vccd1 _12677_/A
+ sky130_fd_sc_hd__nor4_4
X_18589_ _19564_/CLK _18589_/D vssd1 vssd1 vccd1 vccd1 _18589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10513__S0 _10470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10816__S1 _10074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13974__A _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12894__B2 _19537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17880__S _18009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15832__A1 _09339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09727_ _09727_/A _09727_/B vssd1 vssd1 vccd1 vccd1 _09727_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09899__A _09899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09658_ _09658_/A vssd1 vssd1 vccd1 vccd1 _09659_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09589_ _09479_/X _09525_/X _09566_/X _09581_/X _10205_/A vssd1 vssd1 vccd1 vccd1
+ _09589_/X sky130_fd_sc_hd__a311o_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _12475_/B _11910_/A vssd1 vssd1 vccd1 vccd1 _17391_/C sky130_fd_sc_hd__nand2_1
XFILLER_70_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12949__A2 _12946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11551_ _11554_/A _11552_/C _11552_/A vssd1 vssd1 vccd1 vccd1 _11551_/X sky130_fd_sc_hd__a21o_1
XANTENNA__14744__S _14746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10502_ _18780_/Q _19051_/Q _19275_/Q _19019_/Q _10496_/S _09855_/A vssd1 vssd1 vccd1
+ vccd1 _10502_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14270_ _14281_/A vssd1 vssd1 vccd1 vccd1 _14279_/S sky130_fd_sc_hd__buf_2
X_11482_ _11482_/A _11482_/B vssd1 vssd1 vccd1 vccd1 _11482_/X sky130_fd_sc_hd__and2_1
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12772__B _12772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13221_ _18479_/Q _13219_/X _13278_/S vssd1 vssd1 vccd1 vccd1 _13222_/A sky130_fd_sc_hd__mux2_1
X_10433_ _10314_/X _10426_/X _10428_/X _10432_/X _09604_/A vssd1 vssd1 vccd1 vccd1
+ _10433_/X sky130_fd_sc_hd__a311o_1
XFILLER_164_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input64_A io_ibus_inst[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ _19714_/Q vssd1 vssd1 vccd1 vccd1 _16864_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10364_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10365_/A sky130_fd_sc_hd__or2_1
XFILLER_151_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15575__S _15583_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12103_ _12195_/A vssd1 vssd1 vccd1 vccd1 _17884_/A sky130_fd_sc_hd__buf_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _16617_/B _12752_/X _12753_/X _17053_/B _13082_/X vssd1 vssd1 vccd1 vccd1
+ _15679_/B sky130_fd_sc_hd__a221o_2
X_17960_ _17985_/A _17960_/B vssd1 vssd1 vccd1 vccd1 _17960_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10295_ _18815_/Q _19150_/Q _10417_/S vssd1 vssd1 vccd1 vccd1 _10295_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16911_ _19735_/Q vssd1 vssd1 vccd1 vccd1 _16925_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_12034_ _19826_/Q _19825_/Q _12034_/C vssd1 vssd1 vccd1 vccd1 _12092_/C sky130_fd_sc_hd__and3_1
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17891_ _17886_/X _17890_/Y _12117_/B _17754_/A vssd1 vssd1 vccd1 vccd1 _17891_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_19630_ _19768_/CLK _19630_/D vssd1 vssd1 vccd1 vccd1 _19630_/Q sky130_fd_sc_hd__dfxtp_1
X_16842_ _16845_/A _16853_/D vssd1 vssd1 vccd1 vccd1 _16842_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19561_ _19561_/CLK _19561_/D vssd1 vssd1 vccd1 vccd1 _19561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13985_ _13985_/A vssd1 vssd1 vccd1 vccd1 _13994_/S sky130_fd_sc_hd__buf_4
X_16773_ _16773_/A _16773_/B _16774_/B vssd1 vssd1 vccd1 vccd1 _19695_/D sky130_fd_sc_hd__nor3_1
XFILLER_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13823__S _13829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18512_ _19491_/CLK _18512_/D vssd1 vssd1 vccd1 vccd1 _18512_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15724_ _13587_/X _15722_/X _15723_/Y _12903_/X _18447_/Q vssd1 vssd1 vccd1 vccd1
+ _15724_/X sky130_fd_sc_hd__a32o_4
X_12936_ _18438_/Q _09464_/X _11302_/A _12947_/A _12935_/X vssd1 vssd1 vccd1 vccd1
+ _18438_/D sky130_fd_sc_hd__a221o_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19492_ _19493_/CLK _19492_/D vssd1 vssd1 vccd1 vccd1 _19492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09602__A _09602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18443_ _19930_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_2
X_15655_ _14669_/X _19319_/Q _15655_/S vssd1 vssd1 vccd1 vccd1 _15656_/A sky130_fd_sc_hd__mux2_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _19862_/Q _12842_/X _12863_/X _17187_/A _12866_/X vssd1 vssd1 vccd1 vccd1
+ _12867_/X sky130_fd_sc_hd__a221o_1
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11818_ _12029_/C vssd1 vssd1 vccd1 vccd1 _11818_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14606_ _14605_/X _18873_/Q _14606_/S vssd1 vssd1 vccd1 vccd1 _14607_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18374_ _18414_/A vssd1 vssd1 vccd1 vccd1 _18374_/X sky130_fd_sc_hd__clkbuf_2
X_15586_ _15586_/A vssd1 vssd1 vccd1 vccd1 _19288_/D sky130_fd_sc_hd__clkbuf_1
X_12798_ _12818_/B _12798_/B vssd1 vssd1 vccd1 vccd1 _12798_/Y sky130_fd_sc_hd__nor2_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _14559_/A vssd1 vssd1 vccd1 vccd1 _14546_/S sky130_fd_sc_hd__buf_2
XFILLER_105_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17325_ _17325_/A _17325_/B vssd1 vssd1 vccd1 vccd1 _17325_/X sky130_fd_sc_hd__or2_1
XANTENNA__14654__S _14654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ _11778_/A _11749_/B _11920_/A vssd1 vssd1 vccd1 vccd1 _11749_/X sky130_fd_sc_hd__and3_1
XFILLER_30_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17256_ _13595_/A _19853_/Q _17258_/S vssd1 vssd1 vccd1 vccd1 _17257_/A sky130_fd_sc_hd__mux2_1
X_14468_ _14672_/A vssd1 vssd1 vccd1 vccd1 _14468_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16207_ _11890_/X _16206_/Y _13592_/B vssd1 vssd1 vccd1 vccd1 _16207_/Y sky130_fd_sc_hd__o21ai_1
X_13419_ _19916_/Q _12901_/B _13483_/A vssd1 vssd1 vccd1 vccd1 _13419_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17187_ _17187_/A _17195_/B vssd1 vssd1 vccd1 vccd1 _17187_/X sky130_fd_sc_hd__or2_1
X_14399_ _18803_/Q _14398_/X _14402_/S vssd1 vssd1 vccd1 vccd1 _14400_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16138_ _16138_/A vssd1 vssd1 vccd1 vccd1 _19484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15485__S _15489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16069_ _13056_/X _19454_/Q _16073_/S vssd1 vssd1 vccd1 vccd1 _16070_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12876__A1 _16528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19828_ _19865_/CLK _19828_/D vssd1 vssd1 vccd1 vccd1 _19828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19759_ _19759_/CLK _19759_/D vssd1 vssd1 vccd1 vccd1 _19759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09512_ _09512_/A vssd1 vssd1 vccd1 vccd1 _09513_/A sky130_fd_sc_hd__buf_2
XANTENNA__11300__A1 _09745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09443_ _09608_/A vssd1 vssd1 vccd1 vccd1 _18311_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11761__B _17429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__A _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10658__A _10849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11851__A2 _11144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09374_ _09374_/A _09375_/A _12720_/A vssd1 vssd1 vccd1 vccd1 _12888_/A sky130_fd_sc_hd__nor3_4
XFILLER_21_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14564__S _14568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10575__C1 _10307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17176__A _17176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10080_ _10872_/S vssd1 vssd1 vccd1 vccd1 _11483_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12867__B2 _17187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11428__S _11428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15805__A1 _18462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13770_ _13770_/A vssd1 vssd1 vccd1 vccd1 _18544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10982_ _11025_/A _10975_/X _10981_/X vssd1 vssd1 vccd1 vccd1 _10982_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12721_ _17247_/B _12837_/B vssd1 vssd1 vccd1 vccd1 _12776_/A sky130_fd_sc_hd__nor2_2
XFILLER_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15440_ _15440_/A vssd1 vssd1 vccd1 vccd1 _19223_/D sky130_fd_sc_hd__clkbuf_1
X_12652_ _12664_/A vssd1 vssd1 vccd1 vccd1 _12657_/A sky130_fd_sc_hd__buf_6
XFILLER_90_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13044__B2 _19819_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11603_ _11603_/A _11789_/A _11598_/X vssd1 vssd1 vccd1 vccd1 _11603_/X sky130_fd_sc_hd__or3b_1
XFILLER_90_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15371_ _19193_/Q _15298_/X _15371_/S vssd1 vssd1 vccd1 vccd1 _15372_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12583_ _12579_/X _12582_/Y _12583_/S vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14322_ _18773_/Q _13655_/X _14330_/S vssd1 vssd1 vccd1 vccd1 _14323_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17110_ _17112_/A _17112_/C _17101_/X vssd1 vssd1 vccd1 vccd1 _17110_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18090_ _18090_/A _18090_/B vssd1 vssd1 vccd1 vccd1 _18090_/Y sky130_fd_sc_hd__nor2_1
X_11534_ _11534_/A _11534_/B vssd1 vssd1 vccd1 vccd1 _11534_/X sky130_fd_sc_hd__and2_1
XFILLER_157_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17041_ _17044_/A _17041_/B vssd1 vssd1 vccd1 vccd1 _19774_/D sky130_fd_sc_hd__nor2_1
X_14253_ _13790_/X _18743_/Q _14257_/S vssd1 vssd1 vccd1 vccd1 _14254_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11399__A _11399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11465_ _19481_/Q _19319_/Q _18728_/Q _18498_/Q _10649_/X _10754_/A vssd1 vssd1 vccd1
+ vccd1 _11465_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13204_ _13204_/A vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__clkbuf_2
X_10416_ _18813_/Q _19148_/Q _10416_/S vssd1 vssd1 vccd1 vccd1 _10416_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14184_ _14184_/A vssd1 vssd1 vccd1 vccd1 _18712_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output170_A _16458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10566__C1 _09577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11396_ _19497_/Q _18909_/Q _18946_/Q _18520_/Q _10702_/S _09662_/A vssd1 vssd1 vccd1
+ vccd1 _11396_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13135_ _19781_/Q vssd1 vssd1 vccd1 vccd1 _17062_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10347_ _10486_/A vssd1 vssd1 vccd1 vccd1 _10448_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18992_ _19313_/CLK _18992_/D vssd1 vssd1 vccd1 vccd1 _18992_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14503__A _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _13066_/A vssd1 vssd1 vccd1 vccd1 _13066_/X sky130_fd_sc_hd__clkbuf_2
X_17943_ _12204_/Y _17755_/X _17942_/X _17778_/X vssd1 vssd1 vccd1 vccd1 _17943_/X
+ sky130_fd_sc_hd__a211o_1
X_10278_ _19377_/Q _18991_/Q _19441_/Q _18560_/Q _09926_/S _09887_/A vssd1 vssd1 vccd1
+ vccd1 _10279_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11205__S1 _09954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ _17832_/A _12017_/B vssd1 vssd1 vccd1 vccd1 _12020_/A sky130_fd_sc_hd__xnor2_1
XFILLER_79_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17874_ _17521_/X _17995_/B _17776_/X vssd1 vssd1 vccd1 vccd1 _17874_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_120_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19613_ _19879_/CLK _19613_/D vssd1 vssd1 vccd1 vccd1 _19613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16825_ _19709_/Q _16840_/B _16841_/A vssd1 vssd1 vccd1 vccd1 _16863_/C sky130_fd_sc_hd__and3_1
XFILLER_66_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19544_ _19844_/CLK _19544_/D vssd1 vssd1 vccd1 vccd1 _19544_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_47_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16756_ _16773_/A _16756_/B _16757_/B vssd1 vssd1 vccd1 vccd1 _19689_/D sky130_fd_sc_hd__nor3_1
XFILLER_65_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13968_ _18620_/Q _13685_/X _13972_/S vssd1 vssd1 vccd1 vccd1 _13969_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10716__S0 _09647_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15707_ _15707_/A vssd1 vssd1 vccd1 vccd1 _19331_/D sky130_fd_sc_hd__clkbuf_1
X_19475_ _19569_/CLK _19475_/D vssd1 vssd1 vccd1 vccd1 _19475_/Q sky130_fd_sc_hd__dfxtp_1
X_12919_ _19634_/Q _12911_/X _12918_/X vssd1 vssd1 vccd1 vccd1 _12919_/X sky130_fd_sc_hd__o21a_1
X_13899_ _13899_/A vssd1 vssd1 vccd1 vccd1 _18589_/D sky130_fd_sc_hd__clkbuf_1
X_16687_ _16689_/B _16689_/C _16667_/X vssd1 vssd1 vccd1 vccd1 _16687_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18426_ _18426_/A _18426_/B vssd1 vssd1 vccd1 vccd1 _20049_/D sky130_fd_sc_hd__nor2_1
X_15638_ _14644_/X _19311_/Q _15644_/S vssd1 vssd1 vccd1 vccd1 _15639_/A sky130_fd_sc_hd__mux2_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18357_ input56/X vssd1 vssd1 vccd1 vccd1 _18357_/Y sky130_fd_sc_hd__clkinv_4
X_15569_ _15569_/A vssd1 vssd1 vccd1 vccd1 _19280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09885__S1 _09858_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17308_ _17308_/A vssd1 vssd1 vccd1 vccd1 _19876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18288_ _18288_/A _18311_/B vssd1 vssd1 vccd1 vccd1 _18288_/X sky130_fd_sc_hd__or2_1
XFILLER_147_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17239_ _15833_/X _17229_/X _17238_/X _17232_/X vssd1 vssd1 vccd1 vccd1 _19846_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13301__B _13301_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10417__S _10417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18380__A _18380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17485__A0 _17960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13728__S _13736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__A1 _09957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16104__S _16106_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ _19478_/Q _19316_/Q _18725_/Q _18495_/Q _10824_/S _09957_/A vssd1 vssd1 vccd1
+ vccd1 _09993_/B sky130_fd_sc_hd__mux4_1
XFILLER_135_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09507__A _10244_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15943__S _15951_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09226__B _20049_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17788__A1 _17792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11772__A _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15244__A _15244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10707__S0 _10644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09426_ _09426_/A _09426_/B _12601_/B vssd1 vssd1 vccd1 vccd1 _11690_/D sky130_fd_sc_hd__or3_1
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09357_ _18345_/A _19771_/Q _19770_/Q vssd1 vssd1 vccd1 vccd1 _09357_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09896__B _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14294__S _14294_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16075__A _16132_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09288_ _12935_/A vssd1 vssd1 vccd1 vccd1 _18313_/A sky130_fd_sc_hd__clkinv_2
XANTENNA_clkbuf_leaf_167_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11012__A _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11250_ _11250_/A _11250_/B vssd1 vssd1 vccd1 vccd1 _11250_/X sky130_fd_sc_hd__or2_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17476__A0 _12407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ _18785_/Q _19056_/Q _19280_/Q _19024_/Q _10160_/S _09809_/A vssd1 vssd1 vccd1
+ vccd1 _10201_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15419__A _15430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11181_ _11183_/A _11180_/X _10988_/A vssd1 vssd1 vccd1 vccd1 _11181_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_162_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11760__A1 _11348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10132_ _09680_/A _10131_/X _09706_/A vssd1 vssd1 vccd1 vccd1 _10132_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09417__A input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15853__S _15857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ _10063_/A vssd1 vssd1 vccd1 vccd1 _10063_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14940_ _14940_/A vssd1 vssd1 vccd1 vccd1 _19011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11512__A1 _10039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17779__A1 _11940_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10946__S0 _09530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input27_A io_dbus_rdata[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14871_ _14871_/A vssd1 vssd1 vccd1 vccd1 _18980_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14469__S _14472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16610_ _16609_/A _16609_/B _19644_/Q vssd1 vssd1 vccd1 vccd1 _16611_/C sky130_fd_sc_hd__a21oi_1
X_13822_ _14647_/A vssd1 vssd1 vccd1 vccd1 _13822_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17590_ _17496_/X _17498_/X _17590_/S vssd1 vssd1 vccd1 vccd1 _17590_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13265__B2 _19528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13753_ _13746_/X _18539_/Q _13765_/S vssd1 vssd1 vccd1 vccd1 _13754_/A sky130_fd_sc_hd__mux2_1
X_16541_ _16549_/D vssd1 vssd1 vccd1 vccd1 _16547_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10965_ _11025_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10965_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12704_ _12704_/A vssd1 vssd1 vccd1 vccd1 _12704_/X sky130_fd_sc_hd__clkbuf_2
X_19260_ _19392_/CLK _19260_/D vssd1 vssd1 vccd1 vccd1 _19260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13684_ _15254_/A vssd1 vssd1 vccd1 vccd1 _14631_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16472_ _16472_/A vssd1 vssd1 vccd1 vccd1 _19592_/D sky130_fd_sc_hd__clkbuf_1
X_10896_ _11489_/A _10890_/X _10895_/X _09975_/A vssd1 vssd1 vccd1 vccd1 _10896_/X
+ sky130_fd_sc_hd__o211a_1
X_18211_ _18268_/S vssd1 vssd1 vccd1 vccd1 _18220_/S sky130_fd_sc_hd__clkbuf_2
X_15423_ _15423_/A vssd1 vssd1 vccd1 vccd1 _19215_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_184_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19756_/CLK sky130_fd_sc_hd__clkbuf_16
X_12635_ _12635_/A vssd1 vssd1 vccd1 vccd1 _12635_/X sky130_fd_sc_hd__clkbuf_1
X_19191_ _19511_/CLK _19191_/D vssd1 vssd1 vccd1 vccd1 _19191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15354_ _19185_/Q _15273_/X _15356_/S vssd1 vssd1 vccd1 vccd1 _15355_/A sky130_fd_sc_hd__mux2_1
X_18142_ _13115_/A _19963_/Q _18148_/S vssd1 vssd1 vccd1 vccd1 _18143_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12566_ _12588_/B _12565_/Y _12628_/A vssd1 vssd1 vccd1 vccd1 _12566_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11517_ _11470_/A _12668_/B _11584_/A vssd1 vssd1 vccd1 vccd1 _11535_/A sky130_fd_sc_hd__a21boi_1
XFILLER_8_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14305_ _14305_/A vssd1 vssd1 vccd1 vccd1 _18765_/D sky130_fd_sc_hd__clkbuf_1
X_15285_ _15285_/A vssd1 vssd1 vccd1 vccd1 _19156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18073_ _18054_/X _17745_/Y _18071_/X _18072_/X vssd1 vssd1 vccd1 vccd1 _18073_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12497_ _12473_/X _12666_/B _12474_/X _12496_/X vssd1 vssd1 vccd1 vccd1 _18079_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_144_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output95_A _12620_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17024_ _17027_/C _17025_/C _19764_/Q vssd1 vssd1 vccd1 vccd1 _17026_/B sky130_fd_sc_hd__a21oi_1
X_14236_ _14236_/A vssd1 vssd1 vccd1 vccd1 _18735_/D sky130_fd_sc_hd__clkbuf_1
X_11448_ _11448_/A _11448_/B vssd1 vssd1 vccd1 vccd1 _11448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11426__S1 _11371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14167_ _14167_/A vssd1 vssd1 vccd1 vccd1 _18704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11379_ _10730_/A _11376_/X _11378_/X _09976_/X vssd1 vssd1 vccd1 vccd1 _11379_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _19648_/Q _13116_/X _13117_/X _19780_/Q vssd1 vssd1 vccd1 vccd1 _15693_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09327__A _13578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_122_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19293_/CLK sky130_fd_sc_hd__clkbuf_16
X_14098_ _18676_/Q _13651_/X _14098_/S vssd1 vssd1 vccd1 vccd1 _14099_/A sky130_fd_sc_hd__mux2_1
X_18975_ _19553_/CLK _18975_/D vssd1 vssd1 vccd1 vccd1 _18975_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _19907_/Q _17925_/X _18085_/S vssd1 vssd1 vccd1 vccd1 _17927_/A sky130_fd_sc_hd__mux2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13049_ _18931_/Q vssd1 vssd1 vccd1 vccd1 _13371_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09761__S _09761_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17857_ _17560_/X _17847_/Y _17856_/X _17598_/X vssd1 vssd1 vccd1 vccd1 _17857_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16808_ _16808_/A _16808_/B _20018_/Q _16808_/D vssd1 vssd1 vccd1 vccd1 _16809_/D
+ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_137_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19392_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10700__S _10700_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17788_ _17792_/A _17792_/B _18077_/S vssd1 vssd1 vccd1 vccd1 _17788_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19527_ _19542_/CLK _19527_/D vssd1 vssd1 vccd1 vccd1 _19527_/Q sky130_fd_sc_hd__dfxtp_2
X_16739_ _16783_/A vssd1 vssd1 vccd1 vccd1 _16775_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10165__S1 _10148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13008__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19458_ _19552_/CLK _19458_/D vssd1 vssd1 vccd1 vccd1 _19458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13008__B2 _13007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09211_ _11648_/A _11638_/A _11601_/A vssd1 vssd1 vccd1 vccd1 _11673_/A sky130_fd_sc_hd__nor3_4
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18409_ _18409_/A _18409_/B vssd1 vssd1 vccd1 vccd1 _20042_/D sky130_fd_sc_hd__nor2_1
XFILLER_50_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ _19389_/CLK _19389_/D vssd1 vssd1 vccd1 vccd1 _19389_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15003__S _15011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10778__C1 _10010_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15705__A0 _19900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17458__A0 _17820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__A _10672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09975_ _09975_/A vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10950__C1 _10949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10928__S0 _10040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11706__S _12937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13247__B2 _19527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10750_ _11359_/A vssd1 vssd1 vccd1 vccd1 _12076_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ _19812_/Q _19807_/Q vssd1 vssd1 vccd1 vccd1 _09409_/X sky130_fd_sc_hd__and2_1
X_10681_ _09814_/A _10678_/X _10680_/X vssd1 vssd1 vccd1 vccd1 _10681_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10846__A _10846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12420_ _12420_/A vssd1 vssd1 vccd1 vccd1 _15806_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_166_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12222__A2 _12653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11430__B1 _09989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ _12429_/A vssd1 vssd1 vccd1 vccd1 _17525_/A sky130_fd_sc_hd__buf_2
XFILLER_126_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16533__A _18281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ _11302_/A _12632_/B vssd1 vssd1 vccd1 vccd1 _11302_/Y sky130_fd_sc_hd__nand2_1
X_15070_ _14586_/X _19069_/Q _15072_/S vssd1 vssd1 vccd1 vccd1 _15071_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12282_ _12232_/A _12232_/B _12259_/A _12281_/X vssd1 vssd1 vccd1 vccd1 _12283_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_142_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13183__B1 _13343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14021_ _14021_/A vssd1 vssd1 vccd1 vccd1 _18642_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11677__A _12670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ _09746_/A _11219_/X _11231_/X _09753_/A _11232_/Y vssd1 vssd1 vccd1 vccd1
+ _12634_/B sky130_fd_sc_hd__o32ai_4
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11164_ _11283_/A vssd1 vssd1 vccd1 vccd1 _11164_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__15583__S _15583_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10115_ _11387_/A _10110_/Y _10114_/Y _10794_/A vssd1 vssd1 vccd1 vccd1 _10115_/X
+ sky130_fd_sc_hd__o211a_1
X_18760_ _19063_/CLK _18760_/D vssd1 vssd1 vccd1 vccd1 _18760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15972_ _15972_/A vssd1 vssd1 vccd1 vccd1 _19411_/D sky130_fd_sc_hd__clkbuf_1
X_11095_ _11087_/X _11089_/X _11094_/X _10994_/X vssd1 vssd1 vccd1 vccd1 _11095_/Y
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__13486__A1 _13007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_54_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19411_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_103_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17711_ _17469_/X _17428_/X _17800_/S vssd1 vssd1 vccd1 vccd1 _17711_/X sky130_fd_sc_hd__mux2_1
X_10046_ _10000_/X _10012_/Y _10032_/X _10045_/Y _09738_/A vssd1 vssd1 vccd1 vccd1
+ _10046_/X sky130_fd_sc_hd__o311a_1
X_14923_ _14923_/A vssd1 vssd1 vccd1 vccd1 _19003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18691_ _19058_/CLK _18691_/D vssd1 vssd1 vccd1 vccd1 _18691_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output133_A _12671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10395__S1 _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17642_ _17803_/S _17642_/B vssd1 vssd1 vccd1 vccd1 _17642_/Y sky130_fd_sc_hd__nor2_1
X_14854_ _14586_/X _18973_/Q _14856_/S vssd1 vssd1 vccd1 vccd1 _14855_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13805_ _13805_/A vssd1 vssd1 vccd1 vccd1 _18555_/D sky130_fd_sc_hd__clkbuf_1
X_17573_ _17465_/X _17450_/X _17573_/S vssd1 vssd1 vccd1 vccd1 _17573_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_69_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19027_/CLK sky130_fd_sc_hd__clkbuf_16
X_14785_ _14785_/A vssd1 vssd1 vccd1 vccd1 _18946_/D sky130_fd_sc_hd__clkbuf_1
X_11997_ _11997_/A vssd1 vssd1 vccd1 vccd1 _12002_/A sky130_fd_sc_hd__clkinv_2
XFILLER_91_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19312_ _19476_/CLK _19312_/D vssd1 vssd1 vccd1 vccd1 _19312_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12997__B1 _12996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16524_ _16527_/B _16527_/C _12908_/X vssd1 vssd1 vccd1 vccd1 _16524_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13736_ _18536_/Q _13735_/X _13736_/S vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10948_ _11319_/A _10948_/B vssd1 vssd1 vccd1 vccd1 _10948_/X sky130_fd_sc_hd__or2_1
X_19243_ _19405_/CLK _19243_/D vssd1 vssd1 vccd1 vccd1 _19243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16455_ _17123_/A vssd1 vssd1 vccd1 vccd1 _16455_/X sky130_fd_sc_hd__clkbuf_4
X_13667_ _15241_/A vssd1 vssd1 vccd1 vccd1 _14618_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10879_ _11319_/A vssd1 vssd1 vccd1 vccd1 _11250_/A sky130_fd_sc_hd__clkbuf_2
X_15406_ _14621_/X _19208_/Q _15406_/S vssd1 vssd1 vccd1 vccd1 _15407_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19174_ _19402_/CLK _19174_/D vssd1 vssd1 vccd1 vccd1 _19174_/Q sky130_fd_sc_hd__dfxtp_1
X_12618_ _12618_/A _12618_/B _12618_/C vssd1 vssd1 vccd1 vccd1 _12620_/A sky130_fd_sc_hd__nand3_4
X_13598_ _13597_/X _18505_/Q _13598_/S vssd1 vssd1 vccd1 vccd1 _13599_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17137__C1 _16480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16386_ _16386_/A vssd1 vssd1 vccd1 vccd1 _19551_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13410__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18125_ _12620_/Y _17755_/A _18124_/X _12951_/A vssd1 vssd1 vccd1 vccd1 _18125_/X
+ sky130_fd_sc_hd__a211o_1
X_15337_ _19177_/Q _15247_/X _15345_/S vssd1 vssd1 vccd1 vccd1 _15338_/A sky130_fd_sc_hd__mux2_1
X_12549_ _12473_/X _12668_/B _12474_/X _12548_/X vssd1 vssd1 vccd1 vccd1 _18098_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_172_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18056_ _18058_/A _18058_/B _18088_/S vssd1 vssd1 vccd1 vccd1 _18056_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15268_ _19151_/Q _15267_/X _15277_/S vssd1 vssd1 vccd1 vccd1 _15269_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12690__B _12837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13278__S _13278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17007_ _17007_/A _17013_/C vssd1 vssd1 vccd1 vccd1 _17007_/Y sky130_fd_sc_hd__nor2_1
X_14219_ _14219_/A vssd1 vssd1 vccd1 vccd1 _18728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15199_ hold10/A vssd1 vssd1 vccd1 vccd1 _15299_/S sky130_fd_sc_hd__buf_6
XFILLER_98_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10932__C1 _10063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09760_ _12593_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _11534_/A sky130_fd_sc_hd__or2_1
XANTENNA__17860__B1 _17859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18958_ _19027_/CLK _18958_/D vssd1 vssd1 vccd1 vccd1 _18958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17909_ _17521_/X _17971_/B _17776_/X vssd1 vssd1 vccd1 vccd1 _17909_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09691_ _10988_/A vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__clkbuf_2
X_18889_ _19313_/CLK _18889_/D vssd1 vssd1 vccd1 vccd1 _18889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09520__A _09520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10215__B2 _19915_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14572__S _14572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12881__A _17346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16353__A _19953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11963__B2 _18340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10605__S _10735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11176__C1 _09736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10923__C1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13916__S _13922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09958_ _18821_/Q _19156_/Q _10826_/S vssd1 vssd1 vccd1 vccd1 _09958_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13468__A1 _13467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09767__S0 _09763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _10229_/A _09889_/B vssd1 vssd1 vccd1 vccd1 _09889_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _11920_/A vssd1 vssd1 vccd1 vccd1 _11920_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _09998_/A _11144_/X _11156_/X _10065_/A _11157_/Y vssd1 vssd1 vccd1 vccd1
+ _11899_/B sky130_fd_sc_hd__o32ai_4
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18159__A1 _19971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10129__S1 _09662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16528__A _16528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _19494_/Q _18906_/Q _18943_/Q _18517_/Q _10617_/X _10682_/A vssd1 vssd1 vccd1
+ vccd1 _10802_/X sky130_fd_sc_hd__mux4_2
XANTENNA__12979__B1 _10137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _13847_/X _18862_/Q _14572_/S vssd1 vssd1 vccd1 vccd1 _14571_/A sky130_fd_sc_hd__mux2_1
X_11782_ _12155_/B vssd1 vssd1 vccd1 vccd1 _11782_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09430__A _20042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733_ _18678_/Q _19173_/Q _10735_/S vssd1 vssd1 vccd1 vccd1 _10734_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13521_ _13066_/X _13520_/X _13174_/A vssd1 vssd1 vccd1 vccd1 _13521_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14048__A _14059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16240_ _16248_/C _16240_/B vssd1 vssd1 vccd1 vccd1 _16240_/Y sky130_fd_sc_hd__nand2_1
X_13452_ _13324_/X _13437_/X _13440_/Y _13451_/X vssd1 vssd1 vccd1 vccd1 _15279_/A
+ sky130_fd_sc_hd__a22o_2
X_10664_ _11460_/A _10664_/B vssd1 vssd1 vccd1 vccd1 _10664_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12403_ _12473_/A _12661_/B _12402_/Y vssd1 vssd1 vccd1 vccd1 _18033_/B sky130_fd_sc_hd__o21a_1
X_16171_ _16171_/A vssd1 vssd1 vccd1 vccd1 _19499_/D sky130_fd_sc_hd__clkbuf_1
X_13383_ _19871_/Q _12913_/X _13343_/X _19838_/Q vssd1 vssd1 vccd1 vccd1 _13383_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ _18778_/Q _19049_/Q _19273_/Q _19017_/Q _10591_/S _10396_/A vssd1 vssd1 vccd1
+ vccd1 _10595_/X sky130_fd_sc_hd__mux4_2
XANTENNA__12791__A _16875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15122_ _15122_/A vssd1 vssd1 vccd1 vccd1 _19092_/D sky130_fd_sc_hd__clkbuf_1
X_12334_ _12283_/A _12283_/B _12308_/A _12333_/Y vssd1 vssd1 vccd1 vccd1 _12335_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_114_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15053_ _19062_/Q _14462_/X _15055_/S vssd1 vssd1 vccd1 vccd1 _15054_/A sky130_fd_sc_hd__mux2_1
X_19930_ _19930_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _19930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12265_ _19531_/Q _12206_/X _12262_/X _12264_/X _12212_/X vssd1 vssd1 vccd1 vccd1
+ _12265_/X sky130_fd_sc_hd__o221a_1
XFILLER_142_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11706__A1 _12935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14004_ _14072_/S vssd1 vssd1 vccd1 vccd1 _14013_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_123_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11216_ _11216_/A _11216_/B vssd1 vssd1 vccd1 vccd1 _11216_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18095__B1 _18094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19861_ _19881_/CLK _19861_/D vssd1 vssd1 vccd1 vccd1 _19861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12196_ _12429_/A _12196_/B vssd1 vssd1 vccd1 vccd1 _12197_/B sky130_fd_sc_hd__nand2_1
Xoutput71 _12675_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_68_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13826__S _13829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18812_ _19051_/CLK _18812_/D vssd1 vssd1 vccd1 vccd1 _18812_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17842__A0 _19902_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 _11740_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[1] sky130_fd_sc_hd__buf_2
Xoutput93 _11767_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[2] sky130_fd_sc_hd__buf_2
XANTENNA__09780__C1 _09605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11147_ _11147_/A _18671_/Q vssd1 vssd1 vccd1 vccd1 _11147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19792_ _19792_/CLK _19792_/D vssd1 vssd1 vccd1 vccd1 _19792_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16202__S _16204_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18743_ _19302_/CLK _18743_/D vssd1 vssd1 vccd1 vccd1 _18743_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09605__A _09605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15955_ _15955_/A vssd1 vssd1 vccd1 vccd1 _19403_/D sky130_fd_sc_hd__clkbuf_1
X_11078_ _19457_/Q _19295_/Q _18704_/Q _18474_/Q _10999_/A _11065_/A vssd1 vssd1 vccd1
+ vccd1 _11079_/B sky130_fd_sc_hd__mux4_1
X_14906_ _14906_/A vssd1 vssd1 vccd1 vccd1 _18996_/D sky130_fd_sc_hd__clkbuf_1
X_10029_ _18821_/Q _19156_/Q _11386_/S vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__mux2_1
XFILLER_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12031__A _19523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18674_ _19491_/CLK _18674_/D vssd1 vssd1 vccd1 vccd1 _18674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15886_ _13321_/X _19373_/Q _15890_/S vssd1 vssd1 vccd1 vccd1 _15887_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17625_ _17919_/A vssd1 vssd1 vccd1 vccd1 _17827_/A sky130_fd_sc_hd__clkbuf_2
X_14837_ _18359_/A _18405_/B vssd1 vssd1 vccd1 vccd1 _18967_/D sky130_fd_sc_hd__nor2_4
XANTENNA__12966__A _17861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17556_ _17554_/X _17555_/Y _09341_/X _12946_/X vssd1 vssd1 vccd1 vccd1 _19893_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_14768_ _14768_/A vssd1 vssd1 vccd1 vccd1 _18938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16507_ _19610_/Q _16507_/B _16692_/B vssd1 vssd1 vccd1 vccd1 _16508_/C sky130_fd_sc_hd__and3_1
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09930__S0 _10218_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ _13719_/A vssd1 vssd1 vccd1 vccd1 _13736_/S sky130_fd_sc_hd__buf_4
XANTENNA__15061__B _18297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17487_ _17973_/B _17899_/B _17488_/S vssd1 vssd1 vccd1 vccd1 _17487_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14699_ _14699_/A vssd1 vssd1 vccd1 vccd1 _18903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19226_ _19389_/CLK _19226_/D vssd1 vssd1 vccd1 vccd1 _19226_/Q sky130_fd_sc_hd__dfxtp_1
X_16438_ _16438_/A vssd1 vssd1 vccd1 vccd1 _19575_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12198__A1 _11411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19157_ _19285_/CLK _19157_/D vssd1 vssd1 vccd1 vccd1 _19157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16369_ _19545_/Q _16368_/X _16369_/S vssd1 vssd1 vccd1 vccd1 _16370_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_41_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18108_ _18111_/A _18111_/B vssd1 vssd1 vccd1 vccd1 _18108_/Y sky130_fd_sc_hd__nand2_1
X_19088_ _19476_/CLK _19088_/D vssd1 vssd1 vccd1 vccd1 _19088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18039_ _17626_/X _17811_/X _18038_/X vssd1 vssd1 vccd1 vccd1 _18039_/X sky130_fd_sc_hd__a21o_1
XFILLER_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13736__S _13736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20001_ _20048_/CLK _20001_/D vssd1 vssd1 vccd1 vccd1 _20001_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12370__A1 _19535_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ _10245_/S vssd1 vssd1 vccd1 vccd1 _09812_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14421__A _14453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09515__A _09515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ _18928_/Q vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__inv_2
XFILLER_100_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15951__S _15951_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10160__S _10160_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _18829_/Q vssd1 vssd1 vccd1 vccd1 _11091_/A sky130_fd_sc_hd__inv_2
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15398__S _15406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10380_ _10380_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10380_/X sky130_fd_sc_hd__or2_1
XFILLER_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12050_ _12050_/A _12050_/B vssd1 vssd1 vccd1 vccd1 _12051_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09988__S0 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11001_ _11001_/A _11001_/B vssd1 vssd1 vccd1 vccd1 _11001_/X sky130_fd_sc_hd__and2_1
XFILLER_117_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15740_ _15739_/X _19337_/Q _15747_/S vssd1 vssd1 vccd1 vccd1 _15741_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _18445_/Q _12951_/X _11355_/A _12947_/X vssd1 vssd1 vccd1 vccd1 _18445_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11903_ _17749_/A _11903_/B vssd1 vssd1 vccd1 vccd1 _11905_/A sky130_fd_sc_hd__xnor2_4
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _15671_/A vssd1 vssd1 vccd1 vccd1 _19325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _18345_/B vssd1 vssd1 vccd1 vccd1 _12883_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17419_/A vssd1 vssd1 vccd1 vccd1 _17460_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_60_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14622_ _14621_/X _18878_/Q _14622_/S vssd1 vssd1 vccd1 vccd1 _14623_/A sky130_fd_sc_hd__mux2_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _19770_/Q vssd1 vssd1 vccd1 vccd1 _12893_/A sky130_fd_sc_hd__clkbuf_2
X_18390_ _18396_/A _18390_/B vssd1 vssd1 vccd1 vccd1 _20032_/D sky130_fd_sc_hd__nor2_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17341_ _09307_/B _09215_/A _17396_/B _17340_/X vssd1 vssd1 vccd1 vccd1 _17342_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14553_ _13822_/X _18854_/Q _14557_/S vssd1 vssd1 vccd1 vccd1 _14554_/A sky130_fd_sc_hd__mux2_1
X_11765_ _11764_/Y _12674_/A _11717_/A vssd1 vssd1 vccd1 vccd1 _11766_/B sky130_fd_sc_hd__o21a_2
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10522__S1 _10462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _19496_/Q _18908_/Q _18945_/Q _18519_/Q _09647_/A _11387_/A vssd1 vssd1 vccd1
+ vccd1 _10716_/X sky130_fd_sc_hd__mux4_2
X_13504_ _13066_/X _13503_/X _13174_/A vssd1 vssd1 vccd1 vccd1 _13504_/X sky130_fd_sc_hd__o21a_1
X_17272_ _15724_/X _19860_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17273_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14484_ _17041_/B _18408_/B vssd1 vssd1 vccd1 vccd1 _18827_/D sky130_fd_sc_hd__nor2_2
XFILLER_41_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11696_ _20041_/Q _11690_/X _11693_/X _11695_/X vssd1 vssd1 vccd1 vccd1 _11696_/X
+ sky130_fd_sc_hd__a31o_1
X_19011_ _19204_/CLK _19011_/D vssd1 vssd1 vccd1 vccd1 _19011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16223_ _19518_/Q _16222_/X _16223_/S vssd1 vssd1 vccd1 vccd1 _16224_/A sky130_fd_sc_hd__mux2_1
X_13435_ _13435_/A vssd1 vssd1 vccd1 vccd1 _18493_/D sky130_fd_sc_hd__clkbuf_1
X_10647_ _10764_/A _10646_/X _09694_/A vssd1 vssd1 vccd1 vccd1 _10647_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11388__C1 _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15101__S _15105_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ _19344_/Q _12759_/X _12704_/X _19534_/Q _13365_/X vssd1 vssd1 vccd1 vccd1
+ _13366_/X sky130_fd_sc_hd__a221o_1
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16154_ _19492_/Q _14602_/A _16156_/S vssd1 vssd1 vccd1 vccd1 _16155_/A sky130_fd_sc_hd__mux2_1
X_10578_ _19371_/Q _18985_/Q _19435_/Q _18554_/Q _10494_/S _10332_/A vssd1 vssd1 vccd1
+ vccd1 _10579_/B sky130_fd_sc_hd__mux4_1
XFILLER_6_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15105_ _14637_/X _19085_/Q _15105_/S vssd1 vssd1 vccd1 vccd1 _15106_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10245__S _10245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12317_ _12314_/X _12315_/Y _12373_/C _12218_/X vssd1 vssd1 vccd1 vccd1 _12317_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_142_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13297_ _19940_/Q _19941_/Q _13297_/C vssd1 vssd1 vccd1 vccd1 _13312_/B sky130_fd_sc_hd__and3_1
X_16085_ _16085_/A vssd1 vssd1 vccd1 vccd1 _19461_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12026__A _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10038__S0 _10640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ _19054_/Q _14436_/X _15044_/S vssd1 vssd1 vccd1 vccd1 _15037_/A sky130_fd_sc_hd__mux2_1
X_19913_ _19919_/CLK _19913_/D vssd1 vssd1 vccd1 vccd1 _19913_/Q sky130_fd_sc_hd__dfxtp_4
X_12248_ _12245_/X _12246_/Y _12494_/A vssd1 vssd1 vccd1 vccd1 _12248_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_142_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12352__A1 _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19844_ _19844_/CLK _19844_/D vssd1 vssd1 vccd1 vccd1 _19844_/Q sky130_fd_sc_hd__dfxtp_1
X_12179_ _12179_/A _12338_/C vssd1 vssd1 vccd1 vccd1 _12179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19775_ _19877_/CLK _19775_/D vssd1 vssd1 vccd1 vccd1 _19775_/Q sky130_fd_sc_hd__dfxtp_1
X_16987_ _19753_/Q _16983_/C _16986_/Y vssd1 vssd1 vccd1 vccd1 _19753_/D sky130_fd_sc_hd__o21a_1
XFILLER_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18726_ _19317_/CLK _18726_/D vssd1 vssd1 vccd1 vccd1 _18726_/Q sky130_fd_sc_hd__dfxtp_1
X_15938_ _19396_/Q _15225_/X _15940_/S vssd1 vssd1 vccd1 vccd1 _15939_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18657_ _19411_/CLK _18657_/D vssd1 vssd1 vccd1 vccd1 _18657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15869_ _15869_/A vssd1 vssd1 vccd1 vccd1 _19365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17608_ _17608_/A _17610_/B vssd1 vssd1 vccd1 vccd1 _17616_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09390_ _09398_/A _12702_/A _11833_/A _09398_/B vssd1 vssd1 vccd1 vccd1 _12798_/B
+ sky130_fd_sc_hd__or4b_2
X_18588_ _19308_/CLK _18588_/D vssd1 vssd1 vccd1 vccd1 _18588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09221__B1_N input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10418__A1 _10368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17539_ _17539_/A vssd1 vssd1 vccd1 vccd1 _17607_/A sky130_fd_sc_hd__buf_2
XFILLER_149_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10513__S1 _10462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17751__C1 _17705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19209_ _19306_/CLK _19209_/D vssd1 vssd1 vccd1 vccd1 _19209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15011__S _15011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11759__B _17675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14850__S _14856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09229__B _20050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16631__A _16631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15247__A _15247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input1_A io_dbus_rdata[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09726_ _18826_/Q _19161_/Q _09726_/S vssd1 vssd1 vccd1 vccd1 _09727_/B sky130_fd_sc_hd__mux2_1
XANTENNA__18231__A0 _19971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10201__S0 _10160_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09657_ _11179_/A vssd1 vssd1 vccd1 vccd1 _09658_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09588_ _09588_/A vssd1 vssd1 vccd1 vccd1 _10205_/A sky130_fd_sc_hd__buf_2
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18293__A _18293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ _11550_/A _11550_/B vssd1 vssd1 vccd1 vccd1 _11550_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11082__B2 _19898_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10501_ _18588_/Q _18849_/Q _18748_/Q _19083_/Q _10392_/S _10397_/X vssd1 vssd1 vccd1
+ vccd1 _10501_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11481_ _18697_/Q _19192_/Q _11481_/S vssd1 vssd1 vccd1 vccd1 _11482_/B sky130_fd_sc_hd__mux2_1
XANTENNA__16017__S _16023_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13230__A _15235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13220_ _13558_/S vssd1 vssd1 vccd1 vccd1 _13278_/S sky130_fd_sc_hd__buf_6
X_10432_ _10426_/A _10429_/X _10431_/X _10307_/X vssd1 vssd1 vccd1 vccd1 _10432_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13151_ _13151_/A vssd1 vssd1 vccd1 vccd1 _18476_/D sky130_fd_sc_hd__clkbuf_1
X_10363_ _10363_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _10364_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14760__S _14764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ _12188_/A _12648_/A _12101_/Y vssd1 vssd1 vccd1 vccd1 _12195_/A sky130_fd_sc_hd__a21oi_1
X_13082_ _19710_/Q _12989_/X _12990_/X _19678_/Q _13081_/X vssd1 vssd1 vccd1 vccd1
+ _13082_/X sky130_fd_sc_hd__a221o_1
XFILLER_152_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10294_ _10294_/A _10294_/B vssd1 vssd1 vccd1 vccd1 _10294_/X sky130_fd_sc_hd__and2_1
XANTENNA_input57_A io_ibus_inst[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16910_ _16919_/A _16910_/B _16918_/D vssd1 vssd1 vccd1 vccd1 _19734_/D sky130_fd_sc_hd__nor3_1
X_12033_ _17176_/A _12034_/C _19826_/Q vssd1 vssd1 vccd1 vccd1 _12033_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11685__A _12602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17890_ _17869_/X _17983_/B _17953_/A vssd1 vssd1 vccd1 vccd1 _17890_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12885__A2 _16678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16841_ _16841_/A _16863_/D _16841_/C vssd1 vssd1 vccd1 vccd1 _16853_/D sky130_fd_sc_hd__and3_1
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16481__C1 _16480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19560_ _19560_/CLK _19560_/D vssd1 vssd1 vccd1 vccd1 _19560_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_9_clock_A _19998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16772_ _19695_/Q _19694_/Q _16772_/C vssd1 vssd1 vccd1 vccd1 _16774_/B sky130_fd_sc_hd__and3_1
XFILLER_168_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13984_ _13984_/A vssd1 vssd1 vccd1 vccd1 _18627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18511_ _19488_/CLK _18511_/D vssd1 vssd1 vccd1 vccd1 _18511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15723_ _15737_/A _18447_/Q vssd1 vssd1 vccd1 vccd1 _15723_/Y sky130_fd_sc_hd__nand2_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _12935_/A _18196_/S _12937_/C vssd1 vssd1 vccd1 vccd1 _12935_/X sky130_fd_sc_hd__and3_1
X_19491_ _19491_/CLK _19491_/D vssd1 vssd1 vccd1 vccd1 _19491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _19930_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _15654_/A vssd1 vssd1 vccd1 vccd1 _19318_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _19336_/Q _12864_/X _13099_/A _19526_/Q _12865_/X vssd1 vssd1 vccd1 vccd1
+ _12866_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14605_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14605_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _12066_/B vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__buf_2
X_18373_ _18413_/A vssd1 vssd1 vccd1 vccd1 _18373_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13124__B _19899_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14935__S _14939_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _19288_/Q _15295_/X _15587_/S vssd1 vssd1 vccd1 vccd1 _15586_/A sky130_fd_sc_hd__mux2_1
X_12797_ _16809_/A _12797_/B vssd1 vssd1 vccd1 vccd1 _12818_/B sky130_fd_sc_hd__or2_2
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17324_ _09269_/D _17337_/B _09265_/X _09266_/X _11619_/A vssd1 vssd1 vccd1 vccd1
+ _17324_/X sky130_fd_sc_hd__o221a_1
X_14536_ _14536_/A vssd1 vssd1 vccd1 vccd1 _18846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _14479_/A _14479_/C vssd1 vssd1 vccd1 vccd1 _11920_/A sky130_fd_sc_hd__nor2_1
XFILLER_147_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17255_ _17255_/A vssd1 vssd1 vccd1 vccd1 _19852_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10820__A1 _09612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14467_ _14467_/A vssd1 vssd1 vccd1 vccd1 _18824_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10820__B2 _19903_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _11786_/A _11787_/A vssd1 vssd1 vccd1 vccd1 _11680_/D sky130_fd_sc_hd__and2b_1
XFILLER_146_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16206_ _16206_/A _19322_/Q vssd1 vssd1 vccd1 vccd1 _16206_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_127_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13418_ _13418_/A _13418_/B _13438_/C vssd1 vssd1 vccd1 vccd1 _13418_/X sky130_fd_sc_hd__or3_1
XFILLER_174_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17186_ _12854_/X _17182_/X _17184_/X _17185_/X vssd1 vssd1 vccd1 vccd1 _19828_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14398_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14398_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12573__A1 _11520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _19484_/Q _14574_/A _16145_/S vssd1 vssd1 vccd1 vccd1 _16138_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14670__S _14670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13349_ _16661_/A _12887_/X _12889_/X _17095_/A _13348_/X vssd1 vssd1 vccd1 vccd1
+ _15768_/B sky130_fd_sc_hd__a221o_4
XFILLER_154_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16451__A _18365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16068_ _16068_/A vssd1 vssd1 vccd1 vccd1 _19453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15019_ _15019_/A vssd1 vssd1 vccd1 vccd1 _19046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19827_ _19865_/CLK _19827_/D vssd1 vssd1 vccd1 vccd1 _19827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17282__A _17304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19758_ _19759_/CLK _19758_/D vssd1 vssd1 vccd1 vccd1 _19758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09511_ _09511_/A vssd1 vssd1 vccd1 vccd1 _09512_/A sky130_fd_sc_hd__clkbuf_4
X_18709_ _19430_/CLK _18709_/D vssd1 vssd1 vccd1 vccd1 _18709_/Q sky130_fd_sc_hd__dfxtp_1
X_19689_ _19804_/CLK _19689_/D vssd1 vssd1 vccd1 vccd1 _19689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10103__A3 _10102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11300__A2 _11289_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09442_ _20028_/Q vssd1 vssd1 vccd1 vccd1 _18288_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11851__A3 _11156_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _09398_/A _09398_/B _20010_/Q _20009_/Q vssd1 vssd1 vccd1 vccd1 _12720_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_40_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15530__A _15587_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15750__A1 _18452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13985__A _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16361__A _16361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13196__S _13196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18288__A _18288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13924__S _13926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_163_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _09709_/A vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09703__A _09703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10981_ _10976_/X _10979_/X _10980_/X vssd1 vssd1 vccd1 vccd1 _10981_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12720_ _12720_/A vssd1 vssd1 vccd1 vccd1 _17247_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ _12651_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _12651_/Y sky130_fd_sc_hd__nor2_2
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17131__S _17245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11602_ _11533_/Y _11534_/X _11598_/X _11599_/X _11601_/X vssd1 vssd1 vccd1 vccd1
+ _11604_/B sky130_fd_sc_hd__o221ai_1
XFILLER_168_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10489__S0 _10439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15370_ _15370_/A vssd1 vssd1 vccd1 vccd1 _19192_/D sky130_fd_sc_hd__clkbuf_1
X_12582_ _12582_/A _12622_/B vssd1 vssd1 vccd1 vccd1 _12582_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14321_ _14367_/S vssd1 vssd1 vccd1 vccd1 _14330_/S sky130_fd_sc_hd__buf_2
XFILLER_23_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11533_ _17327_/A _17395_/A vssd1 vssd1 vccd1 vccd1 _11533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17040_ _19774_/Q vssd1 vssd1 vccd1 vccd1 _17044_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14252_ _14252_/A vssd1 vssd1 vccd1 vccd1 _18742_/D sky130_fd_sc_hd__clkbuf_1
X_11464_ _11464_/A _11464_/B vssd1 vssd1 vccd1 vccd1 _11464_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _10428_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10415_/X sky130_fd_sc_hd__or2_1
X_13203_ _13342_/A vssd1 vssd1 vccd1 vccd1 _13203_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_88_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14183_ _13793_/X _18712_/Q _14185_/S vssd1 vssd1 vccd1 vccd1 _14184_/A sky130_fd_sc_hd__mux2_1
X_11395_ _11395_/A _11395_/B vssd1 vssd1 vccd1 vccd1 _11395_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10346_ _10323_/X _10328_/Y _10336_/X _10345_/Y _09741_/A vssd1 vssd1 vccd1 vccd1
+ _10346_/X sky130_fd_sc_hd__o311a_1
X_13134_ _19649_/Q vssd1 vssd1 vccd1 vccd1 _16627_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18991_ _19314_/CLK _18991_/D vssd1 vssd1 vccd1 vccd1 _18991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output163_A _12567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13065_ _11232_/Y _12814_/B _13520_/S vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17942_ _17928_/X _17931_/X _17941_/X _17776_/X vssd1 vssd1 vccd1 vccd1 _17942_/X
+ sky130_fd_sc_hd__o211a_1
X_10277_ _09711_/A _10264_/Y _10272_/X _10276_/Y _09741_/A vssd1 vssd1 vccd1 vccd1
+ _10277_/X sky130_fd_sc_hd__o311a_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12016_ _17820_/A _12104_/A _12194_/A vssd1 vssd1 vccd1 vccd1 _12017_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11603__C_N _11598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17873_ _17871_/Y _17872_/X _17923_/S vssd1 vssd1 vccd1 vccd1 _17995_/B sky130_fd_sc_hd__mux2_2
XFILLER_94_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19612_ _19879_/CLK _19612_/D vssd1 vssd1 vccd1 vccd1 _19612_/Q sky130_fd_sc_hd__dfxtp_1
X_16824_ _16840_/B _16841_/A _16823_/Y vssd1 vssd1 vccd1 vccd1 _19708_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10964__S1 _09659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19543_ _19844_/CLK _19543_/D vssd1 vssd1 vccd1 vccd1 _19543_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16755_ _19689_/Q _19688_/Q _16755_/C vssd1 vssd1 vccd1 vccd1 _16757_/B sky130_fd_sc_hd__and3_1
XFILLER_47_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13967_ _13967_/A vssd1 vssd1 vccd1 vccd1 _18619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10716__S1 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15706_ _15705_/X _19331_/Q _15720_/S vssd1 vssd1 vccd1 vccd1 _15707_/A sky130_fd_sc_hd__mux2_1
X_19474_ _19508_/CLK _19474_/D vssd1 vssd1 vccd1 vccd1 _19474_/Q sky130_fd_sc_hd__dfxtp_1
X_12918_ _19762_/Q _12912_/X _12916_/X _12917_/X vssd1 vssd1 vccd1 vccd1 _12918_/X
+ sky130_fd_sc_hd__a211o_1
X_16686_ _19669_/Q _16682_/B _16685_/Y vssd1 vssd1 vccd1 vccd1 _19669_/D sky130_fd_sc_hd__o21a_1
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13898_ _13809_/X _18589_/Q _13900_/S vssd1 vssd1 vccd1 vccd1 _13899_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18425_ _18343_/A _18413_/X _18414_/X _18424_/Y vssd1 vssd1 vccd1 vccd1 _18426_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15637_ _15637_/A vssd1 vssd1 vccd1 vccd1 _19310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _16868_/C _12775_/X _12777_/X _16747_/B _12848_/X vssd1 vssd1 vccd1 vccd1
+ _12849_/X sky130_fd_sc_hd__a221o_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18356_ _18356_/A vssd1 vssd1 vccd1 vccd1 _20022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15568_ _19280_/Q _15270_/X _15572_/S vssd1 vssd1 vccd1 vccd1 _15569_/A sky130_fd_sc_hd__mux2_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17706__C1 _17705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17307_ _17228_/Y _19876_/Q _17313_/S vssd1 vssd1 vccd1 vccd1 _17308_/A sky130_fd_sc_hd__mux2_1
X_14519_ _14519_/A vssd1 vssd1 vccd1 vccd1 _18838_/D sky130_fd_sc_hd__clkbuf_1
X_18287_ _19995_/Q _18285_/X _18286_/X _17243_/X vssd1 vssd1 vccd1 vccd1 _19995_/D
+ sky130_fd_sc_hd__o211a_1
X_15499_ _15499_/A vssd1 vssd1 vccd1 vccd1 _19249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17238_ _19846_/Q _17240_/B vssd1 vssd1 vccd1 vccd1 _17238_/X sky130_fd_sc_hd__or2_1
XANTENNA__13301__C _13301_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17169_ _17242_/B vssd1 vssd1 vccd1 vccd1 _17180_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_171_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17485__A1 _17914_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09991_ _18661_/Q _19252_/Q _19414_/Q _18629_/Q _09984_/X _09985_/X vssd1 vssd1 vccd1
+ vccd1 _09991_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12214__A _12214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17237__A1 _15828_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17724__B _17729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13744__S _13744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16120__S _16128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09523__A _09569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10669__A _19907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10707__S1 _10645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10493__C1 _09718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09425_ _09264_/B _09425_/B _11675_/A vssd1 vssd1 vccd1 vccd1 _09426_/B sky130_fd_sc_hd__nand3b_2
XFILLER_80_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15260__A _15260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09356_ _20018_/Q vssd1 vssd1 vccd1 vccd1 _18345_/A sky130_fd_sc_hd__inv_2
XFILLER_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09287_ _12935_/A _18293_/A _09285_/Y _09286_/X _19887_/Q vssd1 vssd1 vccd1 vccd1
+ _09287_/X sky130_fd_sc_hd__o221a_1
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10796__B1 _09693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17187__A _17187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10200_ _10196_/X _10198_/X _10199_/X _10156_/A _09820_/X vssd1 vssd1 vccd1 vccd1
+ _10205_/B sky130_fd_sc_hd__o221a_1
XFILLER_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17476__A1 _17820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11180_ _19486_/Q _18898_/Q _18935_/Q _18509_/Q _11161_/X _11179_/X vssd1 vssd1 vccd1
+ vccd1 _11180_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10131_ _18662_/Q _19253_/Q _19415_/Q _18630_/Q _11449_/S _10718_/A vssd1 vssd1 vccd1
+ vccd1 _10131_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09417__B _17346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _11395_/A _10061_/X _10000_/X vssd1 vssd1 vccd1 vccd1 _10062_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10946__S1 _11236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16030__S _16034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870_ _14608_/X _18980_/Q _14878_/S vssd1 vssd1 vccd1 vccd1 _14871_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13821_ _13821_/A vssd1 vssd1 vccd1 vccd1 _18560_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09433__A _20050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16540_ _19620_/Q _19619_/Q _19618_/Q _16540_/D vssd1 vssd1 vccd1 vccd1 _16549_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_90_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13752_ _13851_/S vssd1 vssd1 vccd1 vccd1 _13765_/S sky130_fd_sc_hd__clkbuf_4
X_10964_ _19105_/Q _18871_/Q _19553_/Q _19201_/Q _10903_/A _09659_/A vssd1 vssd1 vccd1
+ vccd1 _10965_/B sky130_fd_sc_hd__mux4_1
XFILLER_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12703_ _12756_/A vssd1 vssd1 vccd1 vccd1 _12704_/A sky130_fd_sc_hd__clkbuf_2
X_16471_ _18352_/A _16471_/B vssd1 vssd1 vccd1 vccd1 _16472_/A sky130_fd_sc_hd__or2_1
X_13683_ _13683_/A vssd1 vssd1 vccd1 vccd1 _18523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10895_ _10955_/A _10895_/B vssd1 vssd1 vccd1 vccd1 _10895_/X sky130_fd_sc_hd__or2_1
X_18210_ _18210_/A vssd1 vssd1 vccd1 vccd1 _19961_/D sky130_fd_sc_hd__clkbuf_1
X_15422_ _14644_/X _19215_/Q _15428_/S vssd1 vssd1 vccd1 vccd1 _15423_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19190_ _19906_/CLK _19190_/D vssd1 vssd1 vccd1 vccd1 _19190_/Q sky130_fd_sc_hd__dfxtp_1
X_12634_ _17391_/B _12634_/B vssd1 vssd1 vccd1 vccd1 _12635_/A sky130_fd_sc_hd__and2_4
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10236__C1 _09719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18141_ _18141_/A vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__clkbuf_1
X_15353_ _15353_/A vssd1 vssd1 vccd1 vccd1 _19184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12565_ _19846_/Q _12564_/B _12421_/X vssd1 vssd1 vccd1 vccd1 _12565_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14304_ _18765_/Q _13622_/X _14308_/S vssd1 vssd1 vccd1 vccd1 _14305_/A sky130_fd_sc_hd__mux2_1
X_11516_ _11520_/A _12669_/B vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__nand2_1
X_18072_ _18072_/A vssd1 vssd1 vccd1 vccd1 _18072_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15284_ _19156_/Q _15283_/X hold9/A vssd1 vssd1 vccd1 vccd1 _15285_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10882__S0 _11305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12496_ _18340_/A _12568_/B vssd1 vssd1 vccd1 vccd1 _12496_/X sky130_fd_sc_hd__or2_2
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13829__S _13829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17023_ _17027_/C _17025_/C _17022_/Y vssd1 vssd1 vccd1 vccd1 _19763_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17097__A _17122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14235_ _13764_/X _18735_/Q _14235_/S vssd1 vssd1 vccd1 vccd1 _14236_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11447_ _19127_/Q _18893_/Q _19575_/Q _19223_/Q _10649_/X _10754_/A vssd1 vssd1 vccd1
+ vccd1 _11448_/B sky130_fd_sc_hd__mux4_1
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output88_A _12463_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ _11378_/A _11378_/B vssd1 vssd1 vccd1 vccd1 _11378_/X sky130_fd_sc_hd__or2_1
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14166_ _13767_/X _18704_/Q _14174_/S vssd1 vssd1 vccd1 vccd1 _14167_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11751__A2 _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10329_ _18687_/Q _19182_/Q _10496_/S vssd1 vssd1 vccd1 vccd1 _10330_/A sky130_fd_sc_hd__mux2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _13117_/A vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__buf_2
XFILLER_124_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _19455_/CLK _18974_/D vssd1 vssd1 vccd1 vccd1 _18974_/Q sky130_fd_sc_hd__dfxtp_1
X_14097_ _14097_/A vssd1 vssd1 vccd1 vccd1 _18675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _19644_/Q _12887_/A _12889_/A _19776_/Q _13047_/X vssd1 vssd1 vccd1 vccd1
+ _13588_/B sky130_fd_sc_hd__a221o_2
X_17925_ _17920_/X _17924_/Y _12175_/Y _17754_/A vssd1 vssd1 vccd1 vccd1 _17925_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12969__A _12976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17856_ _17626_/X _17848_/Y _17855_/X _17667_/A vssd1 vssd1 vccd1 vccd1 _17856_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_120_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10711__B1 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16807_ _17247_/B _16807_/B _16807_/C _16807_/D vssd1 vssd1 vccd1 vccd1 _16807_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17787_ _18009_/A vssd1 vssd1 vccd1 vccd1 _18077_/S sky130_fd_sc_hd__buf_2
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14999_ _14999_/A vssd1 vssd1 vccd1 vccd1 _19037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16738_ _16773_/A _16738_/B _16738_/C vssd1 vssd1 vccd1 vccd1 _19683_/D sky130_fd_sc_hd__nor3_1
X_19526_ _19956_/CLK _19526_/D vssd1 vssd1 vccd1 vccd1 _19526_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19457_ _19551_/CLK _19457_/D vssd1 vssd1 vccd1 vccd1 _19457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16669_ _16670_/B _16670_/C _16668_/Y vssd1 vssd1 vccd1 vccd1 _19664_/D sky130_fd_sc_hd__o21a_1
XFILLER_62_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09210_ _09272_/B _09272_/A vssd1 vssd1 vccd1 vccd1 _11601_/A sky130_fd_sc_hd__or2b_4
X_18408_ _18409_/A _18408_/B vssd1 vssd1 vccd1 vccd1 _20041_/D sky130_fd_sc_hd__nor2_1
X_19388_ _19389_/CLK _19388_/D vssd1 vssd1 vccd1 vccd1 _19388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10227__C1 _09741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18339_ _12475_/A _12883_/X _18338_/Y _18329_/X vssd1 vssd1 vccd1 vccd1 _20015_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_111_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15705__A1 _17127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12519__A1 _19605_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16115__S _16117_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14424__A _14628_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17458__A1 _12407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10671__B _12650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15954__S _15962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _11378_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09974_/X sky130_fd_sc_hd__or2_1
XFILLER_131_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12879__A _14476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10928__S1 _10910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__A0 _18807_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_36_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16086__A _16132_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09408_ _19815_/Q _19811_/Q _19849_/Q _19816_/Q vssd1 vssd1 vccd1 vccd1 _11837_/A
+ sky130_fd_sc_hd__a22o_1
X_10680_ _10734_/A _10679_/X _10630_/A vssd1 vssd1 vccd1 vccd1 _10680_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ _09339_/A _09339_/B vssd1 vssd1 vccd1 vccd1 _12739_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11430__A1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ _12376_/A _12659_/B _12377_/A _12349_/X vssd1 vssd1 vccd1 vccd1 _18012_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_11301_ _11301_/A vssd1 vssd1 vccd1 vccd1 _12632_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11958__A _19823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12281_ _12256_/A _17445_/A _12280_/X vssd1 vssd1 vccd1 vccd1 _12281_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10862__A _11399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11232_ _19896_/Q vssd1 vssd1 vccd1 vccd1 _11232_/Y sky130_fd_sc_hd__inv_2
X_14020_ _18642_/Q _13643_/X _14024_/S vssd1 vssd1 vccd1 vccd1 _14021_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10616__S0 _10614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ _11178_/A _11163_/B vssd1 vssd1 vccd1 vccd1 _11163_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09862__S _10216_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ _10637_/A _10114_/B vssd1 vssd1 vccd1 vccd1 _10114_/Y sky130_fd_sc_hd__nand2_1
X_15971_ _19411_/Q _15273_/X _15973_/S vssd1 vssd1 vccd1 vccd1 _15972_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11094_ _11178_/A _11090_/X _11093_/X _10980_/X vssd1 vssd1 vccd1 vccd1 _11094_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17710_ _19896_/Q _17558_/X _17708_/X _17709_/Y vssd1 vssd1 vccd1 vccd1 _19896_/D
+ sky130_fd_sc_hd__o22a_1
X_10045_ _10757_/A _10038_/X _10044_/X vssd1 vssd1 vccd1 vccd1 _10045_/Y sky130_fd_sc_hd__o21ai_1
X_14922_ _19003_/Q _14376_/X _14928_/S vssd1 vssd1 vccd1 vccd1 _14923_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18690_ _19512_/CLK _18690_/D vssd1 vssd1 vccd1 vccd1 _18690_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11041__S0 _10914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17641_ _17791_/A vssd1 vssd1 vccd1 vccd1 _18121_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_64_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14853_ _14853_/A vssd1 vssd1 vccd1 vccd1 _18972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output126_A _12663_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13804_ _13803_/X _18555_/Q _13813_/S vssd1 vssd1 vccd1 vccd1 _13805_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17572_ _17460_/X _17463_/X _17573_/S vssd1 vssd1 vccd1 vccd1 _17572_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14784_ _18946_/Q _14414_/X _14786_/S vssd1 vssd1 vccd1 vccd1 _14785_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11996_ _12052_/A _11996_/B vssd1 vssd1 vccd1 vccd1 _11997_/A sky130_fd_sc_hd__or2_1
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19311_ _19311_/CLK _19311_/D vssd1 vssd1 vccd1 vccd1 _19311_/Q sky130_fd_sc_hd__dfxtp_1
X_16523_ _19614_/Q _16519_/C _16522_/Y vssd1 vssd1 vccd1 vccd1 _19614_/D sky130_fd_sc_hd__o21a_1
XFILLER_44_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13735_ _14669_/A vssd1 vssd1 vccd1 vccd1 _13735_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10947_ _18578_/Q _18839_/Q _18738_/Q _19073_/Q _09981_/A _09511_/A vssd1 vssd1 vccd1
+ vccd1 _10948_/B sky130_fd_sc_hd__mux4_1
XFILLER_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17924__A2 _17957_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19242_ _19405_/CLK _19242_/D vssd1 vssd1 vccd1 vccd1 _19242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16454_ _16454_/A vssd1 vssd1 vccd1 vccd1 _19581_/D sky130_fd_sc_hd__clkbuf_1
X_13666_ _13666_/A vssd1 vssd1 vccd1 vccd1 _18519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10878_ _18967_/Q vssd1 vssd1 vccd1 vccd1 _11319_/A sky130_fd_sc_hd__buf_2
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15405_ _15405_/A vssd1 vssd1 vccd1 vccd1 _19207_/D sky130_fd_sc_hd__clkbuf_1
X_19173_ _19272_/CLK _19173_/D vssd1 vssd1 vccd1 vccd1 _19173_/Q sky130_fd_sc_hd__dfxtp_1
X_12617_ _12617_/A _12617_/B vssd1 vssd1 vccd1 vccd1 _12618_/C sky130_fd_sc_hd__xor2_2
X_16385_ _13109_/X _19551_/Q _16393_/S vssd1 vssd1 vccd1 vccd1 _16386_/A sky130_fd_sc_hd__mux2_1
X_13597_ _13597_/A _13597_/B vssd1 vssd1 vccd1 vccd1 _13597_/X sky130_fd_sc_hd__or2_1
XFILLER_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18124_ _17869_/X _17530_/Y _18072_/X _18123_/X vssd1 vssd1 vccd1 vccd1 _18124_/X
+ sky130_fd_sc_hd__o211a_1
X_15336_ _15358_/A vssd1 vssd1 vccd1 vccd1 _15345_/S sky130_fd_sc_hd__buf_2
XFILLER_118_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12548_ _17338_/A _12568_/B vssd1 vssd1 vccd1 vccd1 _12548_/X sky130_fd_sc_hd__or2_2
XFILLER_129_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18055_ _18058_/A _18058_/B vssd1 vssd1 vccd1 vccd1 _18055_/Y sky130_fd_sc_hd__nand2_1
X_15267_ _15267_/A vssd1 vssd1 vccd1 vccd1 _15267_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10772__A _19904_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _19983_/Q _10139_/A _17464_/S vssd1 vssd1 vccd1 vccd1 _12480_/A sky130_fd_sc_hd__mux2_4
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17006_ _17016_/D vssd1 vssd1 vccd1 vccd1 _17013_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14218_ _13844_/X _18728_/Q _14218_/S vssd1 vssd1 vccd1 vccd1 _14219_/A sky130_fd_sc_hd__mux2_1
X_15198_ _18293_/A _15198_/B _15301_/A _15373_/C vssd1 vssd1 vccd1 vccd1 hold10/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_141_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14149_ _16371_/D vssd1 vssd1 vccd1 vccd1 _15918_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_141_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17860__A1 _10775_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18957_ _19377_/CLK _18957_/D vssd1 vssd1 vccd1 vccd1 _18957_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17908_ _17906_/Y _17907_/X _17923_/S vssd1 vssd1 vccd1 vccd1 _17971_/B sky130_fd_sc_hd__mux2_2
X_09690_ _18830_/Q vssd1 vssd1 vccd1 vccd1 _10988_/A sky130_fd_sc_hd__inv_2
XFILLER_67_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18888_ _19314_/CLK _18888_/D vssd1 vssd1 vccd1 vccd1 _18888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17839_ _18083_/A _17839_/B vssd1 vssd1 vccd1 vccd1 _17839_/X sky130_fd_sc_hd__or2_1
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12437__B1 _19602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19509_ _19571_/CLK _19509_/D vssd1 vssd1 vccd1 vccd1 _19509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15949__S _15951_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10682__A _10682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14154__A _14222_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16351__A1 _19541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09957_ _09957_/A vssd1 vssd1 vccd1 vccd1 _09957_/X sky130_fd_sc_hd__buf_4
XFILLER_44_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_183_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19762_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_103_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09767__S1 _09526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09888_ _19477_/Q _19315_/Q _18724_/Q _18494_/Q _09881_/X _10219_/A vssd1 vssd1 vccd1
+ vccd1 _09889_/B sky130_fd_sc_hd__mux4_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10687__C1 _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11850_ _11928_/A _11990_/A vssd1 vssd1 vccd1 vccd1 _11857_/A sky130_fd_sc_hd__nand2_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12979__A1 _18464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _10805_/A _10801_/B vssd1 vssd1 vccd1 vccd1 _10801_/X sky130_fd_sc_hd__or2_1
XFILLER_26_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _11827_/A vssd1 vssd1 vccd1 vccd1 _12155_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13520_ _19922_/Q _13519_/X _13520_/S vssd1 vssd1 vccd1 vccd1 _13520_/X sky130_fd_sc_hd__mux2_1
X_10732_ _10732_/A _10732_/B vssd1 vssd1 vccd1 vccd1 _10732_/X sky130_fd_sc_hd__or2_1
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_121_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18973_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13451_ _13054_/A _13450_/X _13036_/X vssd1 vssd1 vccd1 vccd1 _13451_/X sky130_fd_sc_hd__o21a_1
X_10663_ _19466_/Q _19304_/Q _18713_/Q _18483_/Q _10658_/X _10014_/X vssd1 vssd1 vccd1
+ vccd1 _10664_/B sky130_fd_sc_hd__mux4_1
XFILLER_41_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12402_ _17338_/B _12378_/B _12474_/A vssd1 vssd1 vccd1 vccd1 _12402_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16170_ _19499_/Q _14624_/A _16178_/S vssd1 vssd1 vccd1 vccd1 _16171_/A sky130_fd_sc_hd__mux2_1
X_10594_ _18586_/Q _18847_/Q _18746_/Q _19081_/Q _10494_/S _10332_/A vssd1 vssd1 vccd1
+ vccd1 _10594_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10837__S0 _09984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13382_ _16317_/A _13397_/C _13381_/Y vssd1 vssd1 vccd1 vccd1 _13382_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15121_ _14660_/X _19092_/Q _15127_/S vssd1 vssd1 vccd1 vccd1 _15122_/A sky130_fd_sc_hd__mux2_1
X_12333_ _12279_/A _12306_/A _12332_/Y vssd1 vssd1 vccd1 vccd1 _12333_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_136_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19292_/CLK sky130_fd_sc_hd__clkbuf_16
X_15052_ _15052_/A vssd1 vssd1 vccd1 vccd1 _19061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12264_ _12260_/Y _12263_/X _12583_/S vssd1 vssd1 vccd1 vccd1 _12264_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14003_ _14059_/A vssd1 vssd1 vccd1 vccd1 _14072_/S sky130_fd_sc_hd__buf_6
XANTENNA__15594__S _15600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11215_ _18638_/Q _19229_/Q _19391_/Q _18606_/Q _11085_/A _11164_/X vssd1 vssd1 vccd1
+ vccd1 _11216_/B sky130_fd_sc_hd__mux4_1
XANTENNA__18095__A1 _12538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19860_ _19865_/CLK _19860_/D vssd1 vssd1 vccd1 vccd1 _19860_/Q sky130_fd_sc_hd__dfxtp_1
X_12195_ _12195_/A _12195_/B _12136_/A _17918_/B vssd1 vssd1 vccd1 vccd1 _12196_/B
+ sky130_fd_sc_hd__or4bb_1
X_18811_ _19500_/CLK _18811_/D vssd1 vssd1 vccd1 vccd1 _18811_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput72 _12056_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[10] sky130_fd_sc_hd__buf_2
XANTENNA__17842__A1 _17840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 _12336_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[20] sky130_fd_sc_hd__buf_2
XFILLER_1_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _19166_/Q vssd1 vssd1 vccd1 vccd1 _11146_/Y sky130_fd_sc_hd__inv_2
X_19791_ _19792_/CLK _19791_/D vssd1 vssd1 vccd1 vccd1 _19791_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput94 _12579_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[30] sky130_fd_sc_hd__buf_2
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18742_ _19431_/CLK _18742_/D vssd1 vssd1 vccd1 vccd1 _18742_/Q sky130_fd_sc_hd__dfxtp_1
X_15954_ _19403_/Q _15247_/X _15962_/S vssd1 vssd1 vccd1 vccd1 _15955_/A sky130_fd_sc_hd__mux2_1
X_11077_ _18967_/Q vssd1 vssd1 vccd1 vccd1 _11317_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14905_ _14660_/X _18996_/Q _14911_/S vssd1 vssd1 vccd1 vccd1 _14906_/A sky130_fd_sc_hd__mux2_1
X_10028_ _11495_/S vssd1 vssd1 vccd1 vccd1 _11386_/S sky130_fd_sc_hd__buf_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18673_ _19490_/CLK _18673_/D vssd1 vssd1 vccd1 vccd1 _18673_/Q sky130_fd_sc_hd__dfxtp_1
X_15885_ _15885_/A vssd1 vssd1 vccd1 vccd1 _19372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13842__S _13845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14836_ _18316_/A _14485_/X _14825_/X _14835_/Y vssd1 vssd1 vccd1 vccd1 _18405_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_17624_ _18072_/A vssd1 vssd1 vccd1 vccd1 _17624_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09621__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17555_ _12675_/X _17554_/B _09419_/X vssd1 vssd1 vccd1 vccd1 _17555_/Y sky130_fd_sc_hd__o21ai_1
X_14767_ _18938_/Q _14388_/X _14775_/S vssd1 vssd1 vccd1 vccd1 _14768_/A sky130_fd_sc_hd__mux2_1
X_11979_ _19521_/Q _12120_/A _12214_/A vssd1 vssd1 vccd1 vccd1 _11979_/X sky130_fd_sc_hd__o21a_1
X_16506_ _16507_/B _16692_/B _19610_/Q vssd1 vssd1 vccd1 vccd1 _16508_/B sky130_fd_sc_hd__a21oi_1
X_13718_ _14656_/A vssd1 vssd1 vccd1 vccd1 _13718_/X sky130_fd_sc_hd__clkbuf_2
X_17486_ _17484_/X _17485_/X _17486_/S vssd1 vssd1 vccd1 vccd1 _17486_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09930__S1 _09929_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14698_ _18903_/Q _14395_/X _14702_/S vssd1 vssd1 vccd1 vccd1 _14699_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16437_ _13523_/X _19575_/Q _16437_/S vssd1 vssd1 vccd1 vccd1 _16438_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19225_ _19482_/CLK _19225_/D vssd1 vssd1 vccd1 vccd1 _19225_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14673__S _14676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13649_ _13649_/A vssd1 vssd1 vccd1 vccd1 _18515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19156_ _19510_/CLK _19156_/D vssd1 vssd1 vccd1 vccd1 _19156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10828__S0 _11372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16368_ _15668_/X _16367_/Y _13604_/B vssd1 vssd1 vccd1 vccd1 _16368_/X sky130_fd_sc_hd__a21o_1
XFILLER_173_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18107_ _19922_/Q _17558_/X _18106_/X vssd1 vssd1 vccd1 vccd1 _19922_/D sky130_fd_sc_hd__o21a_1
X_15319_ _19169_/Q _15222_/X _15323_/S vssd1 vssd1 vccd1 vccd1 _15320_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19087_ _19311_/CLK _19087_/D vssd1 vssd1 vccd1 vccd1 _19087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16299_ _16299_/A vssd1 vssd1 vccd1 vccd1 _16300_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18038_ _17533_/X _18035_/X _18037_/Y _17646_/A vssd1 vssd1 vccd1 vccd1 _18038_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_114_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10007__A _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20000_ _20000_/CLK _20000_/D vssd1 vssd1 vccd1 vccd1 _20000_/Q sky130_fd_sc_hd__dfxtp_1
X_09811_ _10161_/A _09810_/X _10256_/A vssd1 vssd1 vccd1 vccd1 _09811_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19989_ _20048_/CLK _19989_/D vssd1 vssd1 vccd1 vccd1 _19989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15009__S _15011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ _09712_/X _09722_/Y _09728_/X _09733_/Y _09741_/X vssd1 vssd1 vccd1 vccd1
+ _09742_/X sky130_fd_sc_hd__o311a_1
XANTENNA__13318__A _13353_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__C _11764_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09673_ _09722_/A _09673_/B vssd1 vssd1 vccd1 vccd1 _09673_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14848__S _14856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16629__A _16629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09531__A _09967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09287__C1 _19887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11094__C1 _10980_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12830__B1 _18413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_53_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19412_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11397__B1 _10056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_68_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19443_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09988__S1 _09970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ _18673_/Q _19168_/Q _11000_/S vssd1 vssd1 vccd1 vccd1 _11001_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09706__A _09706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _12951_/A vssd1 vssd1 vccd1 vccd1 _12951_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17642__B _17642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14758__S _14764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _11898_/X _17690_/A _12137_/A vssd1 vssd1 vccd1 vccd1 _11903_/B sky130_fd_sc_hd__a21o_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15670_ _15669_/X _19325_/Q _15684_/S vssd1 vssd1 vccd1 vccd1 _15671_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _18273_/S vssd1 vssd1 vccd1 vccd1 _18345_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14621_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _11833_/A vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14059__A _14059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _09453_/B _09448_/C _17339_/X _17327_/B _18302_/A vssd1 vssd1 vccd1 vccd1
+ _17340_/X sky130_fd_sc_hd__o32a_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14552_/A vssd1 vssd1 vccd1 vccd1 _18853_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11764_ _11764_/A _11764_/B _11764_/C vssd1 vssd1 vccd1 vccd1 _11764_/Y sky130_fd_sc_hd__nor3_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13503_ _19921_/Q _13502_/X _13520_/S vssd1 vssd1 vccd1 vccd1 _13503_/X sky130_fd_sc_hd__mux2_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _11448_/A _10715_/B vssd1 vssd1 vccd1 vccd1 _10715_/Y sky130_fd_sc_hd__nor2_1
X_17271_ _17317_/S vssd1 vssd1 vccd1 vccd1 _17280_/S sky130_fd_sc_hd__buf_2
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _18324_/A _16811_/A _14481_/X _14482_/Y vssd1 vssd1 vccd1 vccd1 _18408_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11695_ _17391_/B _11853_/S _11690_/X _09608_/A vssd1 vssd1 vccd1 vccd1 _11695_/X
+ sky130_fd_sc_hd__o22a_1
X_19010_ _19493_/CLK _19010_/D vssd1 vssd1 vccd1 vccd1 _19010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16222_ _16222_/A _16222_/B vssd1 vssd1 vccd1 vccd1 _16222_/X sky130_fd_sc_hd__or2_1
X_13434_ _18493_/Q _13433_/X _13434_/S vssd1 vssd1 vccd1 vccd1 _13435_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10646_ _19112_/Q _18878_/Q _19560_/Q _19208_/Q _10644_/X _10645_/X vssd1 vssd1 vccd1
+ vccd1 _10646_/X sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_5_clock_A _19998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_158_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16153_ _16153_/A vssd1 vssd1 vccd1 vccd1 _19491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13365_ _19870_/Q _12913_/X _13343_/X _19837_/Q vssd1 vssd1 vccd1 vccd1 _13365_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10577_ _09615_/A _10567_/X _10576_/X _09622_/A _19908_/Q vssd1 vssd1 vccd1 vccd1
+ _11411_/A sky130_fd_sc_hd__a32o_4
X_15104_ _15104_/A vssd1 vssd1 vccd1 vccd1 _19084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12316_ _19836_/Q _19835_/Q _12316_/C vssd1 vssd1 vccd1 vccd1 _12373_/C sky130_fd_sc_hd__and3_2
XFILLER_142_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16084_ _13195_/X _19461_/Q _16084_/S vssd1 vssd1 vccd1 vccd1 _16085_/A sky130_fd_sc_hd__mux2_1
X_13296_ _13296_/A vssd1 vssd1 vccd1 vccd1 _18484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17817__B _17820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12450__A2_N _12663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15035_ _15046_/A vssd1 vssd1 vccd1 vccd1 _15044_/S sky130_fd_sc_hd__buf_2
X_19912_ _19919_/CLK _19912_/D vssd1 vssd1 vccd1 vccd1 _19912_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10038__S1 _10037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ _12247_/A vssd1 vssd1 vccd1 vccd1 _12494_/A sky130_fd_sc_hd__buf_2
XFILLER_107_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19843_ _19876_/CLK _19843_/D vssd1 vssd1 vccd1 vccd1 _19843_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_111_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12178_ _19591_/Q hold18/A _12178_/C vssd1 vssd1 vccd1 vccd1 _12338_/C sky130_fd_sc_hd__and3_1
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11129_ _11191_/S vssd1 vssd1 vccd1 vccd1 _11129_/X sky130_fd_sc_hd__buf_4
X_19774_ _19877_/CLK _19774_/D vssd1 vssd1 vccd1 vccd1 _19774_/Q sky130_fd_sc_hd__dfxtp_1
X_16986_ _17007_/A _16992_/C vssd1 vssd1 vccd1 vccd1 _16986_/Y sky130_fd_sc_hd__nor2_1
X_18725_ _19092_/CLK _18725_/D vssd1 vssd1 vccd1 vccd1 _18725_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10115__A1 _11387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15937_ _15937_/A vssd1 vssd1 vccd1 vccd1 _19395_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16449__A _16487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10210__S1 _10196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18656_ _19412_/CLK _18656_/D vssd1 vssd1 vccd1 vccd1 _18656_/Q sky130_fd_sc_hd__dfxtp_1
X_15868_ _13195_/X _19365_/Q _15868_/S vssd1 vssd1 vccd1 vccd1 _15869_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16251__A0 _15718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14819_ _18962_/Q _14465_/X _14819_/S vssd1 vssd1 vccd1 vccd1 _14820_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17607_ _17607_/A vssd1 vssd1 vccd1 vccd1 _17607_/X sky130_fd_sc_hd__clkbuf_2
X_18587_ _19306_/CLK _18587_/D vssd1 vssd1 vccd1 vccd1 _18587_/Q sky130_fd_sc_hd__dfxtp_1
X_15799_ _15799_/A vssd1 vssd1 vccd1 vccd1 _15799_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17538_ _17538_/A _17545_/B _17538_/C vssd1 vssd1 vccd1 vccd1 _17539_/A sky130_fd_sc_hd__nor3_2
XANTENNA__12812__B1 _12810_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17469_ _17461_/X _17466_/X _17608_/A vssd1 vssd1 vccd1 vccd1 _17469_/X sky130_fd_sc_hd__mux2_1
X_19208_ _19560_/CLK _19208_/D vssd1 vssd1 vccd1 vccd1 _19208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16306__A1 _19532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__A1 _12097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19139_ _19288_/CLK _19139_/D vssd1 vssd1 vccd1 vccd1 _19139_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17503__A0 _12574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11474__S0 _09532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09229__C _20049_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__A _09526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15962__S _15962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09725_ _09725_/A vssd1 vssd1 vccd1 vccd1 _09725_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14578__S _14590_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15263__A _15263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18231__A1 hold18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10201__S1 _09809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09656_ _18828_/Q vssd1 vssd1 vccd1 vccd1 _11179_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16242__A0 _19521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _10519_/A vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18293__B _18326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10500_ _10500_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10500_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13511__A _16361_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11480_ _09964_/X _11473_/X _11475_/X _11479_/X _09601_/A vssd1 vssd1 vccd1 vccd1
+ _11480_/X sky130_fd_sc_hd__a311o_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10431_ _10476_/A _10431_/B vssd1 vssd1 vccd1 vccd1 _10431_/X sky130_fd_sc_hd__or2_1
XANTENNA__11465__S0 _10649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13150_ _18476_/Q _13149_/X _13196_/S vssd1 vssd1 vccd1 vccd1 _13151_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10362_ _10363_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _10364_/A sky130_fd_sc_hd__and2_1
XFILLER_109_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17637__B _17642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13657__S _13673_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ _12606_/A _12189_/A _12190_/A vssd1 vssd1 vccd1 vccd1 _12101_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10293_ _18687_/Q _19182_/Q _10417_/S vssd1 vssd1 vccd1 vccd1 _10294_/B sky130_fd_sc_hd__mux2_1
X_13081_ _19614_/Q _12861_/X _13080_/X vssd1 vssd1 vccd1 vccd1 _13081_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11217__S0 _10968_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12032_ _12032_/A vssd1 vssd1 vccd1 vccd1 _12855_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11685__B _12600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16840_ _19709_/Q _16840_/B _16848_/D vssd1 vssd1 vccd1 vccd1 _16841_/C sky130_fd_sc_hd__and3_1
XFILLER_77_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16771_ _19694_/Q _16772_/C _19695_/Q vssd1 vssd1 vccd1 vccd1 _16773_/B sky130_fd_sc_hd__a21oi_1
XFILLER_93_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13983_ _18627_/Q _13714_/X _13983_/S vssd1 vssd1 vccd1 vccd1 _13984_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18510_ _19489_/CLK _18510_/D vssd1 vssd1 vccd1 vccd1 _18510_/Q sky130_fd_sc_hd__dfxtp_1
X_15722_ _18447_/Q _15722_/B vssd1 vssd1 vccd1 vccd1 _15722_/X sky130_fd_sc_hd__or2_1
XFILLER_74_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12947_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _19490_/CLK _19490_/D vssd1 vssd1 vccd1 vccd1 _19490_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_84_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ _14666_/X _19318_/Q _15655_/S vssd1 vssd1 vccd1 vccd1 _15654_/A sky130_fd_sc_hd__mux2_1
X_18441_ _19930_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _19773_/Q _12914_/B vssd1 vssd1 vccd1 vccd1 _12865_/X sky130_fd_sc_hd__and2_1
XFILLER_34_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14604_/A vssd1 vssd1 vccd1 vccd1 _18872_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _11816_/A vssd1 vssd1 vccd1 vccd1 _11816_/Y sky130_fd_sc_hd__clkinv_4
X_18372_ _18380_/A _18372_/B vssd1 vssd1 vccd1 vccd1 _20027_/D sky130_fd_sc_hd__nor2_1
XFILLER_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15584_ _15584_/A vssd1 vssd1 vccd1 vccd1 _19287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _19806_/Q input70/X vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__or2_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17323_ _17323_/A _17323_/B vssd1 vssd1 vccd1 vccd1 _17337_/B sky130_fd_sc_hd__or2_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _13796_/X _18846_/Q _14535_/S vssd1 vssd1 vccd1 vccd1 _14536_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11747_ input66/X vssd1 vssd1 vccd1 vccd1 _14479_/A sky130_fd_sc_hd__inv_2
XANTENNA__12270__A1 _18319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15112__S _15116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10281__B1 _09696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17254_ _13591_/B _19852_/Q _17258_/S vssd1 vssd1 vccd1 vccd1 _17255_/A sky130_fd_sc_hd__mux2_1
X_14466_ _18824_/Q _14465_/X _14466_/S vssd1 vssd1 vccd1 vccd1 _14467_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10820__A2 _10808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _11678_/A vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__buf_2
X_16205_ _16205_/A vssd1 vssd1 vccd1 vccd1 _19515_/D sky130_fd_sc_hd__clkbuf_1
X_13417_ _19948_/Q _13417_/B vssd1 vssd1 vccd1 vccd1 _13438_/C sky130_fd_sc_hd__and2_1
X_10629_ _10296_/A _10628_/X _09979_/X vssd1 vssd1 vccd1 vccd1 _10629_/X sky130_fd_sc_hd__o21a_1
X_17185_ _17185_/A vssd1 vssd1 vccd1 vccd1 _17185_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14397_ _14397_/A vssd1 vssd1 vccd1 vccd1 _18802_/D sky130_fd_sc_hd__clkbuf_1
X_16136_ _16204_/S vssd1 vssd1 vccd1 vccd1 _16145_/S sky130_fd_sc_hd__buf_2
X_13348_ _16922_/C _13341_/X _13342_/X _19693_/Q _13347_/X vssd1 vssd1 vccd1 vccd1
+ _13348_/X sky130_fd_sc_hd__a221o_2
XFILLER_6_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16067_ _13033_/X _19453_/Q _16073_/S vssd1 vssd1 vccd1 vccd1 _16068_/A sky130_fd_sc_hd__mux2_1
X_13279_ _13279_/A vssd1 vssd1 vccd1 vccd1 _18483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15018_ _19046_/Q _14411_/X _15022_/S vssd1 vssd1 vccd1 vccd1 _15019_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13522__A1 _13060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19826_ _19859_/CLK _19826_/D vssd1 vssd1 vccd1 vccd1 _19826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold10_A hold10/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19757_ _19759_/CLK _19757_/D vssd1 vssd1 vccd1 vccd1 _19757_/Q sky130_fd_sc_hd__dfxtp_1
X_16969_ _16970_/B _16969_/B vssd1 vssd1 vccd1 vccd1 _19748_/D sky130_fd_sc_hd__nor2_1
XFILLER_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09510_ _10880_/A vssd1 vssd1 vccd1 vccd1 _09511_/A sky130_fd_sc_hd__buf_4
X_18708_ _19555_/CLK _18708_/D vssd1 vssd1 vccd1 vccd1 _18708_/Q sky130_fd_sc_hd__dfxtp_1
X_19688_ _19804_/CLK _19688_/D vssd1 vssd1 vccd1 vccd1 _19688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _12378_/A vssd1 vssd1 vccd1 vccd1 _18328_/A sky130_fd_sc_hd__buf_2
XANTENNA__11300__A3 _11298_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18639_ _19486_/CLK _18639_/D vssd1 vssd1 vccd1 vccd1 _18639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11049__C1 _10063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09372_ _12804_/A _12700_/A _12700_/B vssd1 vssd1 vccd1 vccd1 _13077_/B sky130_fd_sc_hd__and3b_1
XFILLER_80_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09888__S0 _09881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14427__A _14631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13331__A _15257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12013__A1 _16226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__S0 _10649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10690__A _10826_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16463__B1 _16455_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09708_ _10322_/A vssd1 vssd1 vccd1 vccd1 _09709_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13506__A _15289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ _10980_/A vssd1 vssd1 vccd1 vccd1 _10980_/X sky130_fd_sc_hd__buf_2
XFILLER_71_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09639_ _10184_/A vssd1 vssd1 vccd1 vccd1 _09722_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16817__A _16832_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12650_ _12650_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _12650_/Y sky130_fd_sc_hd__nor2_4
XFILLER_130_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11601_ _11601_/A _11601_/B _11519_/B _11534_/B vssd1 vssd1 vccd1 vccd1 _11601_/X
+ sky130_fd_sc_hd__or4bb_1
XFILLER_12_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10489__S1 _10397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12581_ _19607_/Q _19608_/Q _12581_/C vssd1 vssd1 vccd1 vccd1 _12622_/B sky130_fd_sc_hd__and3_1
XFILLER_168_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16028__S _16034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14320_ _14320_/A vssd1 vssd1 vccd1 vccd1 _18772_/D sky130_fd_sc_hd__clkbuf_1
X_11532_ _11532_/A _11603_/A vssd1 vssd1 vccd1 vccd1 _17395_/A sky130_fd_sc_hd__nor2_1
XFILLER_168_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ _13787_/X _18742_/Q _14257_/S vssd1 vssd1 vccd1 vccd1 _14252_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11463_ _18664_/Q _19255_/Q _19417_/Q _18632_/Q _10658_/X _10703_/A vssd1 vssd1 vccd1
+ vccd1 _11464_/B sky130_fd_sc_hd__mux4_1
XFILLER_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14771__S _14775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13202_ _13341_/A vssd1 vssd1 vccd1 vccd1 _13202_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10414_ _19116_/Q _18882_/Q _19564_/Q _19212_/Q _10367_/S _09841_/A vssd1 vssd1 vccd1
+ vccd1 _10415_/B sky130_fd_sc_hd__mux4_1
Xclkbuf_opt_4_0_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_14182_ _14182_/A vssd1 vssd1 vccd1 vccd1 _18711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11394_ _19369_/Q _18983_/Q _19433_/Q _18552_/Q _10640_/S _10637_/A vssd1 vssd1 vccd1
+ vccd1 _11395_/B sky130_fd_sc_hd__mux4_1
XFILLER_99_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ _13133_/A _13170_/B vssd1 vssd1 vccd1 vccd1 _13133_/Y sky130_fd_sc_hd__nor2_1
X_10345_ _10407_/A _10338_/X _10344_/X vssd1 vssd1 vccd1 vccd1 _10345_/Y sky130_fd_sc_hd__o21ai_1
X_18990_ _19311_/CLK _18990_/D vssd1 vssd1 vccd1 vccd1 _18990_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10661__S1 _10645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _13163_/A vssd1 vssd1 vccd1 vccd1 _13520_/S sky130_fd_sc_hd__clkbuf_2
X_17941_ _17765_/X _17932_/Y _17939_/X _17940_/X vssd1 vssd1 vccd1 vccd1 _17941_/X
+ sky130_fd_sc_hd__a211o_1
X_10276_ _09884_/A _10273_/X _10275_/X vssd1 vssd1 vccd1 vccd1 _10276_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11515__B1 _10065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output156_A _12401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ _12069_/A _12644_/A _12039_/C _20050_/Q vssd1 vssd1 vccd1 vccd1 _17832_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_79_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17872_ _17687_/X _17676_/A _17887_/S vssd1 vssd1 vccd1 vccd1 _17872_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19611_ _19769_/CLK _19611_/D vssd1 vssd1 vccd1 vccd1 _19611_/Q sky130_fd_sc_hd__dfxtp_1
X_16823_ _16845_/A _16823_/B vssd1 vssd1 vccd1 vccd1 _16823_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19542_ _19542_/CLK _19542_/D vssd1 vssd1 vccd1 vccd1 _19542_/Q sky130_fd_sc_hd__dfxtp_2
X_13966_ _18619_/Q _13681_/X _13972_/S vssd1 vssd1 vccd1 vccd1 _13967_/A sky130_fd_sc_hd__mux2_1
X_16754_ _19688_/Q _16755_/C _19689_/Q vssd1 vssd1 vccd1 vccd1 _16756_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14011__S _14013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12917_ _12995_/A vssd1 vssd1 vccd1 vccd1 _12917_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15705_ _19900_/Q _17127_/A _15719_/S vssd1 vssd1 vccd1 vccd1 _15705_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19473_ _19570_/CLK _19473_/D vssd1 vssd1 vccd1 vccd1 _19473_/Q sky130_fd_sc_hd__dfxtp_1
X_16685_ _16731_/A _16689_/C vssd1 vssd1 vccd1 vccd1 _16685_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13897_ _13897_/A vssd1 vssd1 vccd1 vccd1 _18588_/D sky130_fd_sc_hd__clkbuf_1
X_18424_ input54/X vssd1 vssd1 vccd1 vccd1 _18424_/Y sky130_fd_sc_hd__inv_8
XFILLER_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15636_ _14640_/X _19310_/Q _15644_/S vssd1 vssd1 vccd1 vccd1 _15637_/A sky130_fd_sc_hd__mux2_1
X_12848_ _16547_/B _12839_/X _12847_/X vssd1 vssd1 vccd1 vccd1 _12848_/X sky130_fd_sc_hd__o21a_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15567_ _15567_/A vssd1 vssd1 vccd1 vccd1 _19279_/D sky130_fd_sc_hd__clkbuf_1
X_18355_ _18365_/A _18355_/B vssd1 vssd1 vccd1 vccd1 _18356_/A sky130_fd_sc_hd__or2_1
XANTENNA__12243__A1 _11749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ _19660_/Q _13527_/B _12888_/A _19792_/Q vssd1 vssd1 vccd1 vccd1 _12786_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10775__A _19903_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11370__S _11372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17306_ _17306_/A vssd1 vssd1 vccd1 vccd1 _19875_/D sky130_fd_sc_hd__clkbuf_1
X_14518_ _13771_/X _18838_/Q _14524_/S vssd1 vssd1 vccd1 vccd1 _14519_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15498_ _19249_/Q _15273_/X _15500_/S vssd1 vssd1 vccd1 vccd1 _15499_/A sky130_fd_sc_hd__mux2_1
X_18286_ _18286_/A _18311_/B vssd1 vssd1 vccd1 vccd1 _18286_/X sky130_fd_sc_hd__or2_1
XFILLER_30_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14449_ _14653_/A vssd1 vssd1 vccd1 vccd1 _14449_/X sky130_fd_sc_hd__clkbuf_2
X_17237_ _15828_/X _17229_/X _17236_/X _17232_/X vssd1 vssd1 vccd1 vccd1 _19845_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17558__A _18019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17168_ _17230_/A vssd1 vssd1 vccd1 vccd1 _17242_/B sky130_fd_sc_hd__buf_2
XFILLER_171_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16119_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16128_/S sky130_fd_sc_hd__buf_4
X_09990_ _11475_/A vssd1 vssd1 vccd1 vccd1 _10730_/A sky130_fd_sc_hd__buf_2
X_17099_ _17108_/A _17104_/C vssd1 vssd1 vccd1 vccd1 _17099_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17293__A _17304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15806__A _15806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10404__S1 _10440_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18434__B2 _18433_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09804__A _19921_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19809_ _19881_/CLK _19809_/D vssd1 vssd1 vccd1 vccd1 _19809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14856__S _14856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15541__A _15587_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _11694_/A vssd1 vssd1 vccd1 vccd1 _17327_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09355_ _20017_/Q vssd1 vssd1 vccd1 vccd1 _16808_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__10685__A _10805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12785__A2 _13142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09286_ _20038_/Q _19998_/Q vssd1 vssd1 vccd1 vccd1 _09286_/X sky130_fd_sc_hd__and2_1
XFILLER_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11993__A0 _19965_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17468__A _17601_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16372__A _16428_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_32_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09938__B1 _09696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10130_ _10846_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _10130_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13498__B1 _13099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18299__A _18299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13935__S _13939_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10061_ _19478_/Q _19316_/Q _18725_/Q _18495_/Q _10777_/A _10010_/X vssd1 vssd1 vccd1
+ vccd1 _10061_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18425__B2 _18424_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13820_ _13819_/X _18560_/Q _13829_/S vssd1 vssd1 vccd1 vccd1 _13821_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09433__B _20049_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10159__S0 _09508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ _13832_/A vssd1 vssd1 vccd1 vccd1 _13851_/S sky130_fd_sc_hd__buf_4
XFILLER_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10963_ _11178_/A vssd1 vssd1 vccd1 vccd1 _11025_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12702_ _12702_/A _15662_/A vssd1 vssd1 vccd1 vccd1 _12756_/A sky130_fd_sc_hd__nor2_4
XFILLER_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10484__B1 _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16470_ _12160_/A _12160_/B _17041_/B vssd1 vssd1 vccd1 vccd1 _19591_/D sky130_fd_sc_hd__a21o_1
X_13682_ _18523_/Q _13681_/X _13694_/S vssd1 vssd1 vccd1 vccd1 _13683_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10894_ _18643_/Q _19234_/Q _19396_/Q _18611_/Q _10893_/X _09512_/A vssd1 vssd1 vccd1
+ vccd1 _10895_/B sky130_fd_sc_hd__mux4_1
X_15421_ _15421_/A vssd1 vssd1 vccd1 vccd1 _19214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12633_ _12637_/A _12633_/B vssd1 vssd1 vccd1 vccd1 _12633_/Y sky130_fd_sc_hd__nor2_4
XFILLER_169_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15352_ _19184_/Q _15270_/X _15356_/S vssd1 vssd1 vccd1 vccd1 _15353_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18140_ _16232_/A _19962_/Q _18148_/S vssd1 vssd1 vccd1 vccd1 _18141_/A sky130_fd_sc_hd__mux2_1
X_12564_ _19846_/Q _12564_/B vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__and2_1
XFILLER_157_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14303_ _14303_/A vssd1 vssd1 vccd1 vccd1 _18764_/D sky130_fd_sc_hd__clkbuf_1
X_11515_ _09998_/A _11504_/X _11513_/X _10065_/A _11514_/Y vssd1 vssd1 vccd1 vccd1
+ _12669_/B sky130_fd_sc_hd__o32a_4
XFILLER_8_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18071_ _17781_/X _17743_/X _18070_/X _17796_/X vssd1 vssd1 vccd1 vccd1 _18071_/X
+ sky130_fd_sc_hd__a211o_1
X_15283_ _15283_/A vssd1 vssd1 vccd1 vccd1 _15283_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12495_ _12490_/Y _12494_/Y _19604_/Q _11771_/X vssd1 vssd1 vccd1 vccd1 _12495_/X
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_7_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10882__S1 _11236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17022_ _17027_/C _17025_/C _17021_/X vssd1 vssd1 vccd1 vccd1 _17022_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14234_ _14234_/A vssd1 vssd1 vccd1 vccd1 _18734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11446_ _09614_/A _11436_/X _11445_/X _09621_/A _19922_/Q vssd1 vssd1 vccd1 vccd1
+ _11470_/A sky130_fd_sc_hd__a32o_4
XFILLER_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14165_ _14222_/S vssd1 vssd1 vccd1 vccd1 _14174_/S sky130_fd_sc_hd__buf_2
X_11377_ _18584_/Q _18845_/Q _18744_/Q _19079_/Q _10073_/X _09957_/A vssd1 vssd1 vccd1
+ vccd1 _11378_/B sky130_fd_sc_hd__mux4_1
XFILLER_113_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15478__A1 _15244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13116_ _13116_/A vssd1 vssd1 vccd1 vccd1 _13116_/X sky130_fd_sc_hd__buf_2
X_10328_ _10436_/A _10328_/B vssd1 vssd1 vccd1 vccd1 _10328_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ _18973_/CLK _18973_/D vssd1 vssd1 vccd1 vccd1 _18973_/Q sky130_fd_sc_hd__dfxtp_1
X_14096_ _18675_/Q _13647_/X _14098_/S vssd1 vssd1 vccd1 vccd1 _14097_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13845__S _13845_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14150__A1 _14844_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _16840_/B _13144_/S _12723_/A _16717_/B _13046_/X vssd1 vssd1 vccd1 vccd1
+ _13047_/X sky130_fd_sc_hd__a221o_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17924_ _17869_/X _17957_/B _17953_/A vssd1 vssd1 vccd1 vccd1 _17924_/Y sky130_fd_sc_hd__o21ai_1
X_10259_ _10373_/A _10259_/B vssd1 vssd1 vccd1 vccd1 _10259_/X sky130_fd_sc_hd__or2_1
XFILLER_67_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10398__S0 _10392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17855_ _17850_/X _17852_/Y _17854_/X vssd1 vssd1 vccd1 vccd1 _17855_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16806_ _20003_/Q _20002_/Q _20001_/Q _19998_/Q vssd1 vssd1 vccd1 vccd1 _16807_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_94_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17841__A _18127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17786_ _17792_/A _17792_/B vssd1 vssd1 vccd1 vccd1 _17786_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14998_ _19037_/Q _14382_/X _15000_/S vssd1 vssd1 vccd1 vccd1 _14999_/A sky130_fd_sc_hd__mux2_1
X_19525_ _19542_/CLK _19525_/D vssd1 vssd1 vccd1 vccd1 _19525_/Q sky130_fd_sc_hd__dfxtp_2
X_16737_ _19683_/Q _16737_/B _16737_/C vssd1 vssd1 vccd1 vccd1 _16738_/C sky130_fd_sc_hd__and3_1
XANTENNA__14676__S _14676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12985__A _19890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13949_ _13949_/A vssd1 vssd1 vccd1 vccd1 _18611_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_3_5_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19456_ _19794_/CLK _19456_/D vssd1 vssd1 vccd1 vccd1 _19456_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11672__C1 _09420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16668_ _16670_/B _16670_/C _16667_/X vssd1 vssd1 vccd1 vccd1 _16668_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10570__S0 _10560_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18407_ _18409_/A _18407_/B vssd1 vssd1 vccd1 vccd1 _20040_/D sky130_fd_sc_hd__nor2_1
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15619_ _15619_/A vssd1 vssd1 vccd1 vccd1 _19302_/D sky130_fd_sc_hd__clkbuf_1
X_19387_ _19576_/CLK _19387_/D vssd1 vssd1 vccd1 vccd1 _19387_/Q sky130_fd_sc_hd__dfxtp_1
X_16599_ _19639_/Q _16593_/B _16598_/Y vssd1 vssd1 vccd1 vccd1 _19639_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18338_ _18338_/A _18345_/B vssd1 vssd1 vccd1 vccd1 _18338_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10778__A1 _10644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18269_ _18269_/A vssd1 vssd1 vccd1 vccd1 _19988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09973_ _18597_/Q _18858_/Q _18757_/Q _19092_/Q _10675_/A _09985_/A vssd1 vssd1 vccd1
+ vccd1 _09974_/B sky130_fd_sc_hd__mux4_1
XFILLER_143_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09534__A _10678_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13056__A _15206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ _19813_/Q _19808_/Q _19809_/Q _19814_/Q vssd1 vssd1 vccd1 vccd1 _09407_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09338_ _20006_/Q _20004_/Q _09338_/C vssd1 vssd1 vccd1 vccd1 _16809_/B sky130_fd_sc_hd__or3_2
XFILLER_138_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17198__A _17242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ _18306_/A _09269_/B _09269_/C _09269_/D vssd1 vssd1 vccd1 vccd1 _09301_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA__14615__A _14615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11300_ _09745_/A _11289_/X _11298_/X _09752_/A _11299_/Y vssd1 vssd1 vccd1 vccd1
+ _11301_/A sky130_fd_sc_hd__o32a_1
XANTENNA__15210__S _15213_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12280_ _12228_/A _12257_/A _12256_/A _17445_/A vssd1 vssd1 vccd1 vccd1 _12280_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11231_ _10920_/X _11221_/Y _11226_/X _11230_/Y _09736_/A vssd1 vssd1 vccd1 vccd1
+ _11231_/X sky130_fd_sc_hd__o311a_2
XFILLER_134_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10616__S1 _11371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11194__B2 _11319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11162_ _19100_/Q _18866_/Q _19548_/Q _19196_/Q _11161_/X _10974_/A vssd1 vssd1 vccd1
+ vccd1 _11163_/B sky130_fd_sc_hd__mux4_1
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13665__S _13673_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _18822_/Q _19157_/Q _10751_/S vssd1 vssd1 vccd1 vccd1 _10114_/B sky130_fd_sc_hd__mux2_1
XANTENNA__15446__A _15502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16041__S _16045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15970_ _15970_/A vssd1 vssd1 vccd1 vccd1 _19410_/D sky130_fd_sc_hd__clkbuf_1
X_11093_ _11170_/A _11093_/B vssd1 vssd1 vccd1 vccd1 _11093_/X sky130_fd_sc_hd__or2_1
XFILLER_103_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input32_A io_dbus_rdata[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09444__A _18311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _10652_/A _10042_/X _10043_/X vssd1 vssd1 vccd1 vccd1 _10044_/X sky130_fd_sc_hd__o21a_1
X_14921_ _14921_/A vssd1 vssd1 vccd1 vccd1 _19002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11041__S1 _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17640_ _17607_/A _17637_/Y _17639_/X _17543_/X vssd1 vssd1 vccd1 vccd1 _17640_/X
+ sky130_fd_sc_hd__a211o_1
X_14852_ _14583_/X _18972_/Q _14856_/S vssd1 vssd1 vccd1 vccd1 _14853_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13803_ _14628_/A vssd1 vssd1 vccd1 vccd1 _13803_/X sky130_fd_sc_hd__clkbuf_1
X_14783_ _14783_/A vssd1 vssd1 vccd1 vccd1 _18945_/D sky130_fd_sc_hd__clkbuf_1
X_17571_ _17568_/X _17569_/X _17660_/S vssd1 vssd1 vccd1 vccd1 _17571_/X sky130_fd_sc_hd__mux2_1
X_11995_ _11995_/A _17457_/A vssd1 vssd1 vccd1 vccd1 _11996_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output119_A _12656_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19310_ _19311_/CLK _19310_/D vssd1 vssd1 vccd1 vccd1 _19310_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10457__B1 _09756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ _15292_/A vssd1 vssd1 vccd1 vccd1 _14669_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16522_ _16550_/A _16527_/C vssd1 vssd1 vccd1 vccd1 _16522_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10946_ _18770_/Q _19041_/Q _19265_/Q _19009_/Q _09530_/A _11236_/A vssd1 vssd1 vccd1
+ vccd1 _10946_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19241_ _19405_/CLK _19241_/D vssd1 vssd1 vccd1 vccd1 _19241_/Q sky130_fd_sc_hd__dfxtp_1
X_13665_ _18519_/Q _13664_/X _13673_/S vssd1 vssd1 vccd1 vccd1 _13666_/A sky130_fd_sc_hd__mux2_1
X_16453_ _18404_/A _16453_/B vssd1 vssd1 vccd1 vccd1 _16454_/A sky130_fd_sc_hd__or2_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10877_ _18771_/Q _19042_/Q _19266_/Q _19010_/Q _09983_/A _10084_/A vssd1 vssd1 vccd1
+ vccd1 _10877_/X sky130_fd_sc_hd__mux4_1
X_15404_ _14618_/X _19207_/Q _15406_/S vssd1 vssd1 vccd1 vccd1 _15405_/A sky130_fd_sc_hd__mux2_1
X_12616_ _18111_/A _12572_/B _17542_/A vssd1 vssd1 vccd1 vccd1 _12617_/B sky130_fd_sc_hd__o21ai_1
X_19172_ _19268_/CLK _19172_/D vssd1 vssd1 vccd1 vccd1 _19172_/Q sky130_fd_sc_hd__dfxtp_1
X_16384_ _16441_/S vssd1 vssd1 vccd1 vccd1 _16393_/S sky130_fd_sc_hd__buf_2
X_13596_ _15806_/A _13596_/B vssd1 vssd1 vccd1 vccd1 _13597_/B sky130_fd_sc_hd__nor2_2
XANTENNA__17137__A1 _19813_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15335_ _15335_/A vssd1 vssd1 vccd1 vccd1 _19176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18123_ _17516_/X _17626_/X _18122_/X vssd1 vssd1 vccd1 vccd1 _18123_/X sky130_fd_sc_hd__a21o_1
X_12547_ _19606_/Q _12537_/X _12543_/Y _12546_/Y vssd1 vssd1 vccd1 vccd1 _12547_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15266_ _15266_/A vssd1 vssd1 vccd1 vccd1 _19150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18054_ _18054_/A vssd1 vssd1 vccd1 vccd1 _18054_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12478_ _18068_/A _12478_/B vssd1 vssd1 vccd1 vccd1 _12481_/A sky130_fd_sc_hd__xnor2_4
X_14217_ _14217_/A vssd1 vssd1 vccd1 vccd1 _18727_/D sky130_fd_sc_hd__clkbuf_1
X_17005_ _19759_/Q _19758_/Q _17005_/C _17005_/D vssd1 vssd1 vccd1 vccd1 _17016_/D
+ sky130_fd_sc_hd__and4_1
X_11429_ _18696_/Q _19191_/Q _11429_/S vssd1 vssd1 vccd1 vccd1 _11429_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_12_0_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15197_ _15197_/A vssd1 vssd1 vccd1 vccd1 _15197_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14148_ _14148_/A _15198_/B vssd1 vssd1 vccd1 vccd1 _16371_/D sky130_fd_sc_hd__nand2_1
XFILLER_140_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11590__D1 _11589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18956_ _19507_/CLK _18956_/D vssd1 vssd1 vccd1 vccd1 _18956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14079_ _18667_/Q _13608_/X _14087_/S vssd1 vssd1 vccd1 vccd1 _14080_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17907_ _17737_/X _17740_/A _17922_/S vssd1 vssd1 vccd1 vccd1 _17907_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18887_ _19313_/CLK _18887_/D vssd1 vssd1 vccd1 vccd1 _18887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17838_ _17836_/Y _17837_/X _17931_/S vssd1 vssd1 vccd1 vccd1 _17839_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10791__S0 _10048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15803__B _18462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17769_ _17772_/A _17772_/B _18109_/S vssd1 vssd1 vccd1 vccd1 _17769_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19508_ _19508_/CLK _19508_/D vssd1 vssd1 vccd1 vccd1 _19508_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10543__S0 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19439_ _19439_/CLK _19439_/D vssd1 vssd1 vccd1 vccd1 _19439_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10439__S _10439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17128__B2 _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11412__A2 _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16126__S _16128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09529__A _09981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11176__A1 _09703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09956_ _10074_/A vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__buf_4
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09887_ _09887_/A vssd1 vssd1 vccd1 vccd1 _10219_/A sky130_fd_sc_hd__buf_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16809__B _16809_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16097__A _16119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _19366_/Q _18980_/Q _19430_/Q _18549_/Q _10073_/X _10609_/A vssd1 vssd1 vccd1
+ vccd1 _10801_/B sky130_fd_sc_hd__mux4_2
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11773_/X _11957_/A _19819_/Q vssd1 vssd1 vccd1 vccd1 _11780_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10731_ _18582_/Q _18843_/Q _18742_/Q _19077_/Q _10675_/X _10609_/X vssd1 vssd1 vccd1
+ vccd1 _10732_/B sky130_fd_sc_hd__mux4_2
XFILLER_159_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13450_ _19918_/Q _13449_/X _13468_/S vssd1 vssd1 vccd1 vccd1 _13450_/X sky130_fd_sc_hd__mux2_1
X_10662_ _10768_/A _10661_/X _09694_/A vssd1 vssd1 vccd1 vccd1 _10662_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _19600_/Q _12363_/X _12397_/X _12400_/Y vssd1 vssd1 vccd1 vccd1 _12401_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_51_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11969__A _11969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ _16317_/A _13397_/C _13054_/A vssd1 vssd1 vccd1 vccd1 _13381_/Y sky130_fd_sc_hd__o21ai_1
X_10593_ _09855_/A _10590_/Y _10592_/Y _10339_/A vssd1 vssd1 vccd1 vccd1 _10593_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10837__S1 _09985_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15120_ _15120_/A vssd1 vssd1 vccd1 vccd1 _19091_/D sky130_fd_sc_hd__clkbuf_1
X_12332_ _12332_/A _17985_/B vssd1 vssd1 vccd1 vccd1 _12332_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09439__A _17339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15875__S _15879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15051_ _19061_/Q _14459_/X _15055_/S vssd1 vssd1 vccd1 vccd1 _15052_/A sky130_fd_sc_hd__mux2_1
X_12263_ _12263_/A _12288_/C vssd1 vssd1 vccd1 vccd1 _12263_/X sky130_fd_sc_hd__xor2_1
XFILLER_135_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14002_ _16134_/A _15918_/A vssd1 vssd1 vccd1 vccd1 _14059_/A sky130_fd_sc_hd__nor2_4
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ _11141_/A _11213_/X _10988_/X vssd1 vssd1 vccd1 vccd1 _11214_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_107_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12194_ _12194_/A vssd1 vssd1 vccd1 vccd1 _12429_/A sky130_fd_sc_hd__buf_2
X_18810_ _19500_/CLK _18810_/D vssd1 vssd1 vccd1 vccd1 _18810_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput73 _12084_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[11] sky130_fd_sc_hd__buf_2
X_11145_ _19102_/Q _18868_/Q _19550_/Q _19198_/Q _11030_/A _09658_/A vssd1 vssd1 vccd1
+ vccd1 _11145_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10812__S _10812_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 _12362_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[21] sky130_fd_sc_hd__buf_2
X_19790_ _19792_/CLK _19790_/D vssd1 vssd1 vccd1 vccd1 _19790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput95 _12620_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[31] sky130_fd_sc_hd__buf_2
XFILLER_96_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18741_ _19268_/CLK _18741_/D vssd1 vssd1 vccd1 vccd1 _18741_/Q sky130_fd_sc_hd__dfxtp_1
X_15953_ _15975_/A vssd1 vssd1 vccd1 vccd1 _15962_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11076_ _18640_/Q _19231_/Q _19393_/Q _18608_/Q _11000_/S _11065_/X vssd1 vssd1 vccd1
+ vccd1 _11076_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10678__A0 _18807_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14904_ _14904_/A vssd1 vssd1 vccd1 vccd1 _18995_/D sky130_fd_sc_hd__clkbuf_1
X_10027_ _10665_/A vssd1 vssd1 vccd1 vccd1 _10030_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_1_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18672_ _19489_/CLK _18672_/D vssd1 vssd1 vccd1 vccd1 _18672_/Q sky130_fd_sc_hd__dfxtp_1
X_15884_ _13309_/X _19372_/Q _15890_/S vssd1 vssd1 vccd1 vccd1 _15885_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17623_ _09345_/X _17558_/X _17621_/X _17622_/Y vssd1 vssd1 vccd1 vccd1 _19894_/D
+ sky130_fd_sc_hd__o22a_1
X_14835_ input42/X vssd1 vssd1 vccd1 vccd1 _14835_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_45_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17554_ _17554_/A _17554_/B _17554_/C vssd1 vssd1 vccd1 vccd1 _17554_/X sky130_fd_sc_hd__and3_1
X_14766_ _14823_/S vssd1 vssd1 vccd1 vccd1 _14775_/S sky130_fd_sc_hd__buf_2
X_11978_ _12116_/A _11972_/Y _11976_/X _11977_/X vssd1 vssd1 vccd1 vccd1 _11978_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10525__S0 _10509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16505_ _16511_/D vssd1 vssd1 vccd1 vccd1 _16692_/B sky130_fd_sc_hd__clkbuf_2
X_13717_ _15279_/A vssd1 vssd1 vccd1 vccd1 _14656_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10929_ _10929_/A _10929_/B vssd1 vssd1 vccd1 vccd1 _10929_/Y sky130_fd_sc_hd__nor2_1
X_17485_ _17960_/B _17914_/B _17488_/S vssd1 vssd1 vccd1 vccd1 _17485_/X sky130_fd_sc_hd__mux2_1
X_14697_ _14697_/A vssd1 vssd1 vccd1 vccd1 _18902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19224_ _19299_/CLK _19224_/D vssd1 vssd1 vccd1 vccd1 _19224_/Q sky130_fd_sc_hd__dfxtp_1
X_16436_ _16436_/A vssd1 vssd1 vccd1 vccd1 _19574_/D sky130_fd_sc_hd__clkbuf_1
X_13648_ _18515_/Q _13647_/X _13652_/S vssd1 vssd1 vccd1 vccd1 _13649_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19155_ _19287_/CLK _19155_/D vssd1 vssd1 vccd1 vccd1 _19155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10828__S1 _09515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13579_ _15818_/A _18438_/Q vssd1 vssd1 vccd1 vccd1 _13579_/Y sky130_fd_sc_hd__nand2_1
X_16367_ _19956_/Q _16367_/B vssd1 vssd1 vccd1 vccd1 _16367_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_12_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18106_ _12559_/Y _17755_/A _18105_/X _12951_/A vssd1 vssd1 vccd1 vccd1 _18106_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09349__A _09349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15318_ _15318_/A vssd1 vssd1 vccd1 vccd1 _19168_/D sky130_fd_sc_hd__clkbuf_1
X_19086_ _19311_/CLK _19086_/D vssd1 vssd1 vccd1 vccd1 _19086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16298_ _16298_/A vssd1 vssd1 vccd1 vccd1 _19531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_79_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18037_ _18121_/B _18032_/Y _18036_/Y vssd1 vssd1 vccd1 vccd1 _18037_/Y sky130_fd_sc_hd__a21oi_1
X_15249_ _19145_/Q _15247_/X _15261_/S vssd1 vssd1 vccd1 vccd1 _15250_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09810_ _18692_/Q _19187_/Q _10195_/S vssd1 vssd1 vccd1 vccd1 _09810_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19988_ _19988_/CLK _19988_/D vssd1 vssd1 vccd1 vccd1 _19988_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12107__A0 _19969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09741_ _09741_/A vssd1 vssd1 vccd1 vccd1 _09741_/X sky130_fd_sc_hd__buf_2
XFILLER_101_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18939_ _19042_/CLK _18939_/D vssd1 vssd1 vccd1 vccd1 _18939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09672_ _19387_/Q _19001_/Q _19451_/Q _18570_/Q _09655_/X _09727_/A vssd1 vssd1 vccd1
+ vccd1 _09673_/B sky130_fd_sc_hd__mux4_1
XFILLER_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09812__A _10245_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10958__A _11202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15025__S _15033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10516__S0 _10509_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12830__A1 _13591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09958__S _10826_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14165__A _14222_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11397__A1 _10052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13138__A2 _12992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17285__A0 _12741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09939_ _18659_/Q _19250_/Q _19412_/Q _18627_/Q _09653_/A _09929_/X vssd1 vssd1 vccd1
+ vccd1 _09940_/B sky130_fd_sc_hd__mux4_1
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12950_ _18444_/Q _12946_/X _10961_/X _12947_/X vssd1 vssd1 vccd1 vccd1 _18444_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _11901_/A _11901_/B _17397_/B _11901_/D vssd1 vssd1 vccd1 vccd1 _12137_/A
+ sky130_fd_sc_hd__or4_4
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _17346_/B vssd1 vssd1 vccd1 vccd1 _18273_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11872__A2 _11864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10868__A _10869_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _14620_/A vssd1 vssd1 vccd1 vccd1 _18877_/D sky130_fd_sc_hd__clkbuf_1
X_11832_ _19819_/Q vssd1 vssd1 vccd1 vccd1 _11843_/A sky130_fd_sc_hd__inv_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _13819_/X _18853_/Q _14557_/S vssd1 vssd1 vccd1 vccd1 _14552_/A sky130_fd_sc_hd__mux2_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11763_/A _11763_/B vssd1 vssd1 vccd1 vccd1 _11766_/A sky130_fd_sc_hd__nor2_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11180__S0 _11161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _19368_/Q _18982_/Q _19432_/Q _18551_/Q _10653_/X _10665_/X vssd1 vssd1 vccd1
+ vccd1 _10715_/B sky130_fd_sc_hd__mux4_1
X_13502_ _16689_/B _12832_/X _12833_/X _17120_/B _13501_/X vssd1 vssd1 vccd1 vccd1
+ _13502_/X sky130_fd_sc_hd__a221o_4
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14482_ input46/X vssd1 vssd1 vccd1 vccd1 _14482_/Y sky130_fd_sc_hd__inv_2
X_17270_ _17270_/A vssd1 vssd1 vccd1 vccd1 _19859_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11694_/A _11895_/C vssd1 vssd1 vccd1 vccd1 _11853_/S sky130_fd_sc_hd__nand2_1
XFILLER_158_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13433_ _15276_/A vssd1 vssd1 vccd1 vccd1 _13433_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16221_ _16232_/C _16220_/Y _12492_/A vssd1 vssd1 vccd1 vccd1 _16222_/B sky130_fd_sc_hd__a21oi_1
X_10645_ _10665_/A vssd1 vssd1 vccd1 vccd1 _10645_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15771__A0 _19912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11388__A1 _10665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16152_ _19491_/Q _14599_/A _16156_/S vssd1 vssd1 vccd1 vccd1 _16153_/A sky130_fd_sc_hd__mux2_1
X_13364_ _19726_/Q vssd1 vssd1 vccd1 vccd1 _16922_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_155_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10576_ _10314_/A _10569_/X _10571_/X _10575_/X _09604_/A vssd1 vssd1 vccd1 vccd1
+ _10576_/X sky130_fd_sc_hd__a311o_2
X_15103_ _14634_/X _19084_/Q _15105_/S vssd1 vssd1 vccd1 vccd1 _15104_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_80_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12315_ _17205_/A _12316_/C _19836_/Q vssd1 vssd1 vccd1 vccd1 _12315_/Y sky130_fd_sc_hd__a21oi_1
X_16083_ _16083_/A vssd1 vssd1 vccd1 vccd1 _19460_/D sky130_fd_sc_hd__clkbuf_1
X_13295_ _18484_/Q _13293_/X _13358_/S vssd1 vssd1 vccd1 vccd1 _13296_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15034_ _15034_/A vssd1 vssd1 vccd1 vccd1 _19053_/D sky130_fd_sc_hd__clkbuf_1
X_19911_ _19919_/CLK _19911_/D vssd1 vssd1 vccd1 vccd1 _19911_/Q sky130_fd_sc_hd__dfxtp_4
X_12246_ _17199_/A _12267_/C _11890_/X vssd1 vssd1 vccd1 vccd1 _12246_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17276__A0 _12874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19842_ _19876_/CLK _19842_/D vssd1 vssd1 vccd1 vccd1 _19842_/Q sky130_fd_sc_hd__dfxtp_1
X_12177_ _12152_/A _12178_/C hold18/A vssd1 vssd1 vccd1 vccd1 _12179_/A sky130_fd_sc_hd__a21oi_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _11317_/A vssd1 vssd1 vccd1 vccd1 _11304_/A sky130_fd_sc_hd__clkbuf_2
X_19773_ _19857_/CLK _19773_/D vssd1 vssd1 vccd1 vccd1 _19773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16985_ _16994_/D vssd1 vssd1 vccd1 vccd1 _16992_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12042__B _17832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18724_ _19481_/CLK _18724_/D vssd1 vssd1 vccd1 vccd1 _18724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11059_ _11059_/A vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__buf_4
X_15936_ _19395_/Q _15222_/X _15940_/S vssd1 vssd1 vccd1 vccd1 _15937_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09632__A _11460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18655_ _19409_/CLK _18655_/D vssd1 vssd1 vccd1 vccd1 _18655_/Q sky130_fd_sc_hd__dfxtp_1
X_15867_ _15867_/A vssd1 vssd1 vccd1 vccd1 _19364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17606_ _17600_/X _17921_/A _17530_/A vssd1 vssd1 vccd1 vccd1 _17606_/Y sky130_fd_sc_hd__a21oi_1
X_14818_ _14818_/A vssd1 vssd1 vccd1 vccd1 _18961_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13065__A1 _12814_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18586_ _19305_/CLK _18586_/D vssd1 vssd1 vccd1 vccd1 _18586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15798_ _15798_/A vssd1 vssd1 vccd1 vccd1 _19347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17537_ _17725_/A vssd1 vssd1 vccd1 vccd1 _17748_/S sky130_fd_sc_hd__clkbuf_2
X_14749_ _14749_/A vssd1 vssd1 vccd1 vccd1 _18926_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16465__A _18352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__S0 _11147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17468_ _17601_/S vssd1 vssd1 vccd1 vccd1 _17608_/A sky130_fd_sc_hd__clkbuf_2
X_19207_ _19559_/CLK _19207_/D vssd1 vssd1 vccd1 vccd1 _19207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16419_ _16419_/A vssd1 vssd1 vccd1 vccd1 _19566_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_182_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19759_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_165_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11379__A1 _10730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17399_ _17504_/S vssd1 vssd1 vccd1 vccd1 _17419_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19138_ _19288_/CLK _19138_/D vssd1 vssd1 vccd1 vccd1 _19138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12040__A2 _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17503__A1 _11764_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18830__D _18830_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19069_ _19391_/CLK _19069_/D vssd1 vssd1 vccd1 vccd1 _19069_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16404__S _16404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10018__A _10018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_120_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19455_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09724_ _18698_/Q _19193_/Q _09724_/S vssd1 vssd1 vccd1 vccd1 _09725_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16490__A1 _19605_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10737__S0 _10614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _09787_/S vssd1 vssd1 vccd1 vccd1 _09655_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_135_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _18836_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09586_ _10623_/A vssd1 vssd1 vccd1 vccd1 _10519_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11162__S0 _11161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_102_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10430_ _19470_/Q _19308_/Q _18717_/Q _18487_/Q _10466_/S _10312_/A vssd1 vssd1 vccd1
+ vccd1 _10431_/B sky130_fd_sc_hd__mux4_1
XFILLER_155_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18298__A2 _18291_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11465__S1 _10754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ _09750_/A _10346_/X _10359_/X _09757_/A _10360_/Y vssd1 vssd1 vccd1 vccd1
+ _12657_/B sky130_fd_sc_hd__o32a_4
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12100_ _12098_/A _12319_/B _12376_/A vssd1 vssd1 vccd1 vccd1 _12190_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__09717__A _09717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13080_ _16958_/B _12991_/X _13079_/X _12995_/X vssd1 vssd1 vccd1 vccd1 _13080_/X
+ sky130_fd_sc_hd__a211o_1
X_10292_ _19118_/Q _18884_/Q _19566_/Q _19214_/Q _10465_/S _10291_/X vssd1 vssd1 vccd1
+ vccd1 _10292_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11217__S1 _11164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _19523_/Q _12120_/A vssd1 vssd1 vccd1 vccd1 _12031_/X sky130_fd_sc_hd__or2_1
XANTENNA__13239__A _15238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09830__S1 _09822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_1_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14769__S _14775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__S _13673_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16770_ _19694_/Q _16772_/C _16769_/Y vssd1 vssd1 vccd1 vccd1 _19694_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13982_ _13982_/A vssd1 vssd1 vccd1 vccd1 _18626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ _15721_/A vssd1 vssd1 vccd1 vccd1 _19333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09452__A _17338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_27_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12933_ _12933_/A _12937_/C vssd1 vssd1 vccd1 vccd1 _12976_/A sky130_fd_sc_hd__nor2_4
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17430__A0 _17642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18440_ _20000_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _15652_/A vssd1 vssd1 vccd1 vccd1 _19317_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12864_/A vssd1 vssd1 vccd1 vccd1 _12864_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17981__A1 _12287_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14602_/X _18872_/Q _14606_/S vssd1 vssd1 vccd1 vccd1 _14604_/A sky130_fd_sc_hd__mux2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _18286_/A _12795_/X _14831_/X _18370_/Y vssd1 vssd1 vccd1 vccd1 _18372_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_11815_ _11815_/A _11815_/B vssd1 vssd1 vccd1 vccd1 _11816_/A sky130_fd_sc_hd__xnor2_4
X_15583_ _19287_/Q _15292_/X _15583_/S vssd1 vssd1 vccd1 vccd1 _15584_/A sky130_fd_sc_hd__mux2_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output101_A _12003_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12795_ _18413_/A vssd1 vssd1 vccd1 vccd1 _12795_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17322_ _17322_/A vssd1 vssd1 vccd1 vccd1 _18301_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ _14534_/A vssd1 vssd1 vccd1 vccd1 _18845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11746_ _16208_/S vssd1 vssd1 vccd1 vccd1 _11778_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17253_ _17253_/A vssd1 vssd1 vccd1 vccd1 _19851_/D sky130_fd_sc_hd__clkbuf_1
X_14465_ _14669_/A vssd1 vssd1 vccd1 vccd1 _14465_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14009__S _14013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11677_ _12670_/A _11692_/C _11693_/C _11676_/X vssd1 vssd1 vccd1 vccd1 _17397_/B
+ sky130_fd_sc_hd__or4b_2
XANTENNA__10820__A3 _10819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16204_ _19515_/Q _14675_/A _16204_/S vssd1 vssd1 vccd1 vccd1 _16205_/A sky130_fd_sc_hd__mux2_1
X_10628_ _19498_/Q _18910_/Q _18947_/Q _18521_/Q _10678_/S _09813_/A vssd1 vssd1 vccd1
+ vccd1 _10628_/X sky130_fd_sc_hd__mux4_2
X_13416_ _16332_/A _13417_/B vssd1 vssd1 vccd1 vccd1 _13418_/B sky130_fd_sc_hd__nor2_1
XFILLER_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17184_ _19828_/Q _17195_/B vssd1 vssd1 vccd1 vccd1 _17184_/X sky130_fd_sc_hd__or2_1
X_14396_ _18802_/Q _14395_/X _14402_/S vssd1 vssd1 vccd1 vccd1 _14397_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13848__S _13851_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16135_ _16191_/A vssd1 vssd1 vccd1 vccd1 _16204_/S sky130_fd_sc_hd__buf_6
X_13347_ _19629_/Q _12891_/X _13346_/X vssd1 vssd1 vccd1 vccd1 _13347_/X sky130_fd_sc_hd__o21a_1
X_10559_ _18810_/Q _19145_/Q _10559_/S vssd1 vssd1 vccd1 vccd1 _10559_/X sky130_fd_sc_hd__mux2_1
X_13278_ _18483_/Q _13277_/X _13278_/S vssd1 vssd1 vccd1 vccd1 _13279_/A sky130_fd_sc_hd__mux2_1
X_16066_ _16066_/A vssd1 vssd1 vccd1 vccd1 _19452_/D sky130_fd_sc_hd__clkbuf_1
X_15017_ _15017_/A vssd1 vssd1 vccd1 vccd1 _19045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13149__A _15222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ _12229_/A _17447_/A vssd1 vssd1 vccd1 vccd1 _12229_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19825_ _19865_/CLK _19825_/D vssd1 vssd1 vccd1 vccd1 _19825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19756_ _19756_/CLK _19756_/D vssd1 vssd1 vccd1 vccd1 _19756_/Q sky130_fd_sc_hd__dfxtp_1
X_16968_ _19748_/Q _16975_/D _16833_/X vssd1 vssd1 vccd1 vccd1 _16969_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12089__A2 _12084_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10719__S0 _10649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19409_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18707_ _19552_/CLK _18707_/D vssd1 vssd1 vccd1 vccd1 _18707_/Q sky130_fd_sc_hd__dfxtp_1
X_15919_ _15975_/A vssd1 vssd1 vccd1 vccd1 _15988_/S sky130_fd_sc_hd__buf_6
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19687_ _19720_/CLK _19687_/D vssd1 vssd1 vccd1 vccd1 _19687_/Q sky130_fd_sc_hd__dfxtp_1
X_16899_ _16924_/C _16906_/D vssd1 vssd1 vccd1 vccd1 _16901_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09440_ _20044_/Q vssd1 vssd1 vccd1 vccd1 _17338_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18638_ _19487_/CLK _18638_/D vssd1 vssd1 vccd1 vccd1 _18638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09371_ _09389_/A _12688_/A _12688_/B _20015_/Q vssd1 vssd1 vccd1 vccd1 _12700_/B
+ sky130_fd_sc_hd__nor4b_1
XFILLER_52_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18569_ _19482_/CLK _18569_/D vssd1 vssd1 vccd1 vccd1 _18569_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15811__B _18463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19286_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09888__S1 _10219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10272__A1 _09929_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16923__A _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11447__S1 _10754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09965__B2 _10840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09537__A _10417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09707_ _09707_/A vssd1 vssd1 vccd1 vccd1 _10322_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09638_ _09936_/A vssd1 vssd1 vccd1 vccd1 _10184_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09569_ _09569_/A vssd1 vssd1 vccd1 vccd1 _09762_/A sky130_fd_sc_hd__buf_2
XFILLER_128_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15213__S _15213_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ _11600_/A _11603_/A vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__or2_1
XFILLER_71_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12580_ _12561_/A _12581_/C _19608_/Q vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__a21oi_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18425__A1_N _18343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15726__A0 _19903_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ _11600_/A vssd1 vssd1 vccd1 vccd1 _17327_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16833__A _16939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__A _11046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14250_ _14250_/A vssd1 vssd1 vccd1 vccd1 _18741_/D sky130_fd_sc_hd__clkbuf_1
X_11462_ _11464_/A _11461_/X _09694_/A vssd1 vssd1 vccd1 vccd1 _11462_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17479__A0 _12328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13201_ _19716_/Q vssd1 vssd1 vccd1 vccd1 _16864_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10413_ _11415_/A _12656_/B vssd1 vssd1 vccd1 vccd1 _11558_/A sky130_fd_sc_hd__or2_1
XFILLER_99_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14181_ _13790_/X _18711_/Q _14185_/S vssd1 vssd1 vccd1 vccd1 _14182_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11393_ _10000_/X _11383_/Y _11388_/X _11392_/Y _09738_/A vssd1 vssd1 vccd1 vccd1
+ _11393_/X sky130_fd_sc_hd__o311a_2
XANTENNA__10881__A _11260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18140__A1 _19962_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13132_ _19931_/Q _19932_/Q _13132_/C vssd1 vssd1 vccd1 vccd1 _13170_/B sky130_fd_sc_hd__and3_1
XANTENNA__12960__B1 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10344_ _10486_/A _10343_/X _09709_/A vssd1 vssd1 vccd1 vccd1 _10344_/X sky130_fd_sc_hd__o21a_1
XANTENNA_input62_A io_ibus_inst[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09447__A _18288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _16206_/A _16219_/A _13066_/A vssd1 vssd1 vccd1 vccd1 _13063_/Y sky130_fd_sc_hd__o21ai_1
X_17940_ _17940_/A vssd1 vssd1 vccd1 vccd1 _17940_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10275_ _10403_/A _10274_/X _09891_/A vssd1 vssd1 vccd1 vccd1 _10275_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11515__A1 _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ _12027_/A _11920_/X _12009_/X _12013_/X vssd1 vssd1 vccd1 vccd1 _16461_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17871_ _17871_/A vssd1 vssd1 vccd1 vccd1 _17871_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__10723__C1 _09717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output149_A _12249_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19610_ _19877_/CLK _19610_/D vssd1 vssd1 vccd1 vccd1 _19610_/Q sky130_fd_sc_hd__dfxtp_1
X_16822_ _16840_/B _16841_/A vssd1 vssd1 vccd1 vccd1 _16823_/B sky130_fd_sc_hd__and2_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19541_ _19956_/CLK _19541_/D vssd1 vssd1 vccd1 vccd1 _19541_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16753_ _19688_/Q _16755_/C _16752_/Y vssd1 vssd1 vccd1 vccd1 _19688_/D sky130_fd_sc_hd__o21a_1
XFILLER_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13965_ _13965_/A vssd1 vssd1 vccd1 vccd1 _18618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11374__S0 _11429_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15704_ _15700_/X _15701_/X _15703_/Y _13577_/A _18444_/Q vssd1 vssd1 vccd1 vccd1
+ _17127_/A sky130_fd_sc_hd__a32o_2
XFILLER_80_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19472_ _19570_/CLK _19472_/D vssd1 vssd1 vccd1 vccd1 _19472_/Q sky130_fd_sc_hd__dfxtp_1
X_12916_ _19874_/Q _12913_/X _12863_/X _19841_/Q _12915_/X vssd1 vssd1 vccd1 vccd1
+ _12916_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16684_ _16684_/A vssd1 vssd1 vccd1 vccd1 _16689_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13896_ _13806_/X _18588_/Q _13900_/S vssd1 vssd1 vccd1 vccd1 _13897_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18423_ _18426_/A _18423_/B vssd1 vssd1 vccd1 vccd1 _20048_/D sky130_fd_sc_hd__nor2_1
XFILLER_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15635_ _15646_/A vssd1 vssd1 vccd1 vccd1 _15644_/S sky130_fd_sc_hd__buf_2
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _19749_/Q _12840_/X _12845_/X _12846_/X vssd1 vssd1 vccd1 vccd1 _12847_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15123__S _15127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11126__S0 _11004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__B1 _12888_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _09328_/C _14476_/A _18414_/A input45/X vssd1 vssd1 vccd1 vccd1 _18355_/B
+ sky130_fd_sc_hd__o22a_1
X_15566_ _19279_/Q _15267_/X _15572_/S vssd1 vssd1 vccd1 vccd1 _15567_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _19724_/Q _12775_/X _12777_/X _19692_/Q vssd1 vssd1 vccd1 vccd1 _12786_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17225_/Y _19875_/Q _17313_/S vssd1 vssd1 vccd1 vccd1 _17306_/A sky130_fd_sc_hd__mux2_1
X_14517_ _14517_/A vssd1 vssd1 vccd1 vccd1 _18837_/D sky130_fd_sc_hd__clkbuf_1
X_18285_ _18323_/A vssd1 vssd1 vccd1 vccd1 _18285_/X sky130_fd_sc_hd__clkbuf_2
X_11729_ _11729_/A _17325_/B vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__or2_1
X_15497_ _15497_/A vssd1 vssd1 vccd1 vccd1 _19248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17236_ _19845_/Q _17240_/B vssd1 vssd1 vccd1 vccd1 _17236_/X sky130_fd_sc_hd__or2_1
X_14448_ _14448_/A vssd1 vssd1 vccd1 vccd1 _18818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ _17197_/A vssd1 vssd1 vccd1 vccd1 _17167_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14379_ _14583_/A vssd1 vssd1 vccd1 vccd1 _14379_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16118_ _16118_/A vssd1 vssd1 vccd1 vccd1 _19476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17098_ _17098_/A vssd1 vssd1 vccd1 vccd1 _17104_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16049_ _16049_/A vssd1 vssd1 vccd1 vccd1 _19445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13607__A _15197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19808_ _19881_/CLK _19808_/D vssd1 vssd1 vccd1 vccd1 _19808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19739_ _19745_/CLK _19739_/D vssd1 vssd1 vccd1 vccd1 _19739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11365__S0 _10690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16918__A _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09423_ _09426_/A _11532_/A _12601_/B vssd1 vssd1 vccd1 vccd1 _11694_/A sky130_fd_sc_hd__or3_1
XFILLER_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15033__S _15033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09354_ _11839_/C _09354_/B vssd1 vssd1 vccd1 vccd1 _11952_/D sky130_fd_sc_hd__and2b_1
XFILLER_40_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13431__B2 _13554_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _20038_/Q _19998_/Q vssd1 vssd1 vccd1 vccd1 _09285_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14872__S _14878_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11993__A1 _11355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13488__S _13524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09938__A1 _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12942__A0 _18321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13498__B2 _19542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18299__B _18326_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ _11399_/A _10060_/B vssd1 vssd1 vccd1 vccd1 _10060_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09797__S0 _09724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15716__B _15716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10640__S _10640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14112__S _14120_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12421__A _15806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10159__S1 _10148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13750_ _18299_/A _14917_/B _15373_/A _15373_/B vssd1 vssd1 vccd1 vccd1 _13832_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10962_ _11096_/A vssd1 vssd1 vccd1 vccd1 _11178_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10484__A1 _09615_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ _12701_/A _17247_/A vssd1 vssd1 vccd1 vccd1 _15662_/A sky130_fd_sc_hd__or2_2
XFILLER_44_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10484__B2 _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16039__S _16045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13681_ _14628_/A vssd1 vssd1 vccd1 vccd1 _13681_/X sky130_fd_sc_hd__clkbuf_2
X_10893_ _11114_/S vssd1 vssd1 vccd1 vccd1 _10893_/X sky130_fd_sc_hd__clkbuf_4
X_15420_ _14640_/X _19214_/Q _15428_/S vssd1 vssd1 vccd1 vccd1 _15421_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12632_ _12637_/A _12632_/B vssd1 vssd1 vccd1 vccd1 _12632_/Y sky130_fd_sc_hd__nor2_4
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15351_ _15351_/A vssd1 vssd1 vccd1 vccd1 _19183_/D sky130_fd_sc_hd__clkbuf_1
X_12563_ _19543_/Q _12122_/X _14477_/B _12562_/X _12123_/X vssd1 vssd1 vccd1 vccd1
+ _12563_/X sky130_fd_sc_hd__o221a_1
XANTENNA__14782__S _14786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11514_ _19923_/Q vssd1 vssd1 vccd1 vccd1 _11514_/Y sky130_fd_sc_hd__inv_2
X_14302_ _18764_/Q _13618_/X _14308_/S vssd1 vssd1 vccd1 vccd1 _14303_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18070_ _17785_/X _18067_/X _18069_/Y _17705_/A vssd1 vssd1 vccd1 vccd1 _18070_/X
+ sky130_fd_sc_hd__o211a_1
X_15282_ _15282_/A vssd1 vssd1 vccd1 vccd1 _19155_/D sky130_fd_sc_hd__clkbuf_1
X_12494_ _12494_/A _12494_/B vssd1 vssd1 vccd1 vccd1 _12494_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17021_ _17101_/A vssd1 vssd1 vccd1 vccd1 _17021_/X sky130_fd_sc_hd__buf_2
X_11445_ _09476_/A _11438_/X _11440_/X _11444_/X _09603_/A vssd1 vssd1 vccd1 vccd1
+ _11445_/X sky130_fd_sc_hd__a311o_1
X_14233_ _13761_/X _18734_/Q _14235_/S vssd1 vssd1 vccd1 vccd1 _14234_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11736__A1 _12097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10095__S0 _10081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ _14164_/A vssd1 vssd1 vccd1 vccd1 _18703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11376_ _18776_/Q _19047_/Q _19271_/Q _19015_/Q _10675_/X _09957_/X vssd1 vssd1 vccd1
+ vccd1 _11376_/X sky130_fd_sc_hd__mux4_2
XFILLER_124_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10327_ _19118_/Q _18884_/Q _19566_/Q _19214_/Q _10325_/X _10326_/X vssd1 vssd1 vccd1
+ vccd1 _10328_/B sky130_fd_sc_hd__mux4_1
X_13115_ _13115_/A _13132_/C vssd1 vssd1 vccd1 vccd1 _13115_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18972_ _19196_/CLK _18972_/D vssd1 vssd1 vccd1 vccd1 _18972_/Q sky130_fd_sc_hd__dfxtp_1
X_14095_ _14095_/A vssd1 vssd1 vccd1 vccd1 _18674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _16518_/B _12911_/X _13045_/X vssd1 vssd1 vccd1 vccd1 _13046_/X sky130_fd_sc_hd__o21a_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _17921_/Y _17922_/X _17923_/S vssd1 vssd1 vccd1 vccd1 _17957_/B sky130_fd_sc_hd__mux2_2
X_10258_ _19473_/Q _19311_/Q _18720_/Q _18490_/Q _09901_/A _09842_/A vssd1 vssd1 vccd1
+ vccd1 _10259_/B sky130_fd_sc_hd__mux4_1
XANTENNA__14150__A2 _16809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10398__S1 _10397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17854_ _17976_/A _17851_/X _17853_/X _17533_/A vssd1 vssd1 vccd1 vccd1 _17854_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14022__S _14024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10189_ _19475_/Q _19313_/Q _18722_/Q _18492_/Q _09881_/X _10219_/A vssd1 vssd1 vccd1
+ vccd1 _10189_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16805_ _19995_/Q _19994_/Q _19992_/Q _19993_/Q vssd1 vssd1 vccd1 vccd1 _16807_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17785_ _17785_/A vssd1 vssd1 vccd1 vccd1 _17785_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14957__S _14961_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14997_ _14997_/A vssd1 vssd1 vccd1 vccd1 _19036_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13861__S _13867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19524_ _19542_/CLK _19524_/D vssd1 vssd1 vccd1 vccd1 _19524_/Q sky130_fd_sc_hd__dfxtp_2
X_16736_ _16737_/B _16737_/C _19683_/Q vssd1 vssd1 vccd1 vccd1 _16738_/B sky130_fd_sc_hd__a21oi_1
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13948_ _18611_/Q _13647_/X _13950_/S vssd1 vssd1 vccd1 vccd1 _13949_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19455_ _19455_/CLK _19455_/D vssd1 vssd1 vccd1 vccd1 _19455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16667_ _16860_/A vssd1 vssd1 vccd1 vccd1 _16667_/X sky130_fd_sc_hd__buf_2
XANTENNA__11672__B1 _11910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13879_ _13879_/A vssd1 vssd1 vccd1 vccd1 _18580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18406_ _18409_/A _18406_/B vssd1 vssd1 vccd1 vccd1 _20039_/D sky130_fd_sc_hd__nor2_1
X_15618_ _14615_/X _19302_/Q _15622_/S vssd1 vssd1 vccd1 vccd1 _15619_/A sky130_fd_sc_hd__mux2_1
X_19386_ _19576_/CLK _19386_/D vssd1 vssd1 vccd1 vccd1 _19386_/Q sky130_fd_sc_hd__dfxtp_1
X_16598_ _16631_/A _16600_/B vssd1 vssd1 vccd1 vccd1 _16598_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18337_ _12688_/A _18323_/X _18336_/X _18329_/X vssd1 vssd1 vccd1 vccd1 _20014_/D
+ sky130_fd_sc_hd__o211a_1
X_15549_ _15549_/A vssd1 vssd1 vccd1 vccd1 _19271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18268_ _19988_/Q _19609_/Q _18268_/S vssd1 vssd1 vccd1 vccd1 _18269_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_149_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17219_ _17217_/Y _17212_/X _17218_/X _17215_/X vssd1 vssd1 vccd1 vccd1 _19839_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18199_ _18255_/A vssd1 vssd1 vccd1 vccd1 _18268_/S sky130_fd_sc_hd__buf_2
XANTENNA__18104__A1 _17705_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10086__S0 _10081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09972_ _11489_/A vssd1 vssd1 vccd1 vccd1 _11378_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12940__S _17808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13101__B1 _13099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15552__A _15574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09550__A _10368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09406_ _19883_/Q _11952_/C vssd1 vssd1 vccd1 vccd1 _09406_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09337_ _20008_/Q _20007_/Q _20005_/Q vssd1 vssd1 vccd1 vccd1 _09338_/C sky130_fd_sc_hd__or3_1
XFILLER_40_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13800__A _13832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _09272_/B vssd1 vssd1 vccd1 vccd1 _18306_/A sky130_fd_sc_hd__inv_2
XFILLER_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09199_ _09272_/A _09272_/B vssd1 vssd1 vccd1 vccd1 _11627_/C sky130_fd_sc_hd__and2_1
XFILLER_147_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12915__B1 _12756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ _11221_/A _11227_/X _11229_/X vssd1 vssd1 vccd1 vccd1 _11230_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13946__S _13950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ _11327_/S vssd1 vssd1 vccd1 vccd1 _11161_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14631__A _14631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10112_ _10112_/A vssd1 vssd1 vccd1 vccd1 _10637_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11092_ _18768_/Q _19039_/Q _19263_/Q _19007_/Q _11035_/A _11179_/A vssd1 vssd1 vccd1
+ vccd1 _11093_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10043_ _10043_/A vssd1 vssd1 vccd1 vccd1 _10043_/X sky130_fd_sc_hd__clkbuf_4
X_14920_ _19002_/Q _14369_/X _14928_/S vssd1 vssd1 vccd1 vccd1 _14921_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input25_A io_dbus_rdata[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851_ _14851_/A vssd1 vssd1 vccd1 vccd1 _18971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13802_ _13802_/A vssd1 vssd1 vccd1 vccd1 _18554_/D sky130_fd_sc_hd__clkbuf_1
X_17570_ _17674_/S vssd1 vssd1 vccd1 vccd1 _17660_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14782_ _18945_/Q _14411_/X _14786_/S vssd1 vssd1 vccd1 vccd1 _14783_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11994_ _11995_/A _17457_/A vssd1 vssd1 vccd1 vccd1 _12052_/A sky130_fd_sc_hd__and2_1
XFILLER_17_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10457__A1 _09749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16521_ _16529_/D vssd1 vssd1 vccd1 vccd1 _16527_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13733_ _13733_/A vssd1 vssd1 vccd1 vccd1 _18535_/D sky130_fd_sc_hd__clkbuf_1
X_10945_ _10938_/X _10942_/X _10944_/X _11250_/A _09472_/A vssd1 vssd1 vccd1 vccd1
+ _10951_/B sky130_fd_sc_hd__o221a_1
XFILLER_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14078__A _14146_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19240_ _19402_/CLK _19240_/D vssd1 vssd1 vccd1 vccd1 _19240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16452_ _16449_/X _11796_/X _11798_/X _18412_/A vssd1 vssd1 vccd1 vccd1 _19580_/D
+ sky130_fd_sc_hd__a211o_1
X_13664_ _14615_/A vssd1 vssd1 vccd1 vccd1 _13664_/X sky130_fd_sc_hd__clkbuf_2
X_10876_ _10871_/X _10873_/X _10874_/X _11014_/A _10875_/X vssd1 vssd1 vccd1 vccd1
+ _10885_/B sky130_fd_sc_hd__o221a_1
X_15403_ _15403_/A vssd1 vssd1 vccd1 vccd1 _19206_/D sky130_fd_sc_hd__clkbuf_1
X_19171_ _19288_/CLK _19171_/D vssd1 vssd1 vccd1 vccd1 _19171_/Q sky130_fd_sc_hd__dfxtp_1
X_12615_ _18121_/A _12615_/B vssd1 vssd1 vccd1 vccd1 _12617_/A sky130_fd_sc_hd__nand2_2
X_16383_ _16383_/A vssd1 vssd1 vccd1 vccd1 _19550_/D sky130_fd_sc_hd__clkbuf_1
X_13595_ _13595_/A vssd1 vssd1 vccd1 vccd1 _13596_/B sky130_fd_sc_hd__inv_2
XFILLER_12_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11501__S0 _10040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13710__A _14650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18122_ _12615_/B _17634_/X _18120_/X _18121_/Y _17646_/A vssd1 vssd1 vccd1 vccd1
+ _18122_/X sky130_fd_sc_hd__a41o_1
X_15334_ _19176_/Q _15244_/X _15334_/S vssd1 vssd1 vccd1 vccd1 _15335_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16345__A0 _19540_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12546_ _12314_/X _12544_/Y _12564_/B _12537_/A vssd1 vssd1 vccd1 vccd1 _12546_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_150_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18053_ _18053_/A vssd1 vssd1 vccd1 vccd1 _19917_/D sky130_fd_sc_hd__clkbuf_1
X_15265_ _19150_/Q _15263_/X _15277_/S vssd1 vssd1 vccd1 vccd1 _15266_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12477_ _12427_/A _12429_/B _18058_/A _17525_/A vssd1 vssd1 vccd1 vccd1 _12478_/B
+ sky130_fd_sc_hd__o31a_2
X_17004_ _17046_/A _17004_/B _17004_/C vssd1 vssd1 vccd1 vccd1 _19758_/D sky130_fd_sc_hd__nor3_1
XANTENNA_output93_A _11767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _13841_/X _18727_/Q _14218_/S vssd1 vssd1 vccd1 vccd1 _14217_/A sky130_fd_sc_hd__mux2_1
X_11428_ _18824_/Q _19159_/Q _11428_/S vssd1 vssd1 vccd1 vccd1 _11428_/X sky130_fd_sc_hd__mux2_1
X_15196_ _15196_/A vssd1 vssd1 vccd1 vccd1 _19129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14147_ _14147_/A vssd1 vssd1 vccd1 vccd1 _18698_/D sky130_fd_sc_hd__clkbuf_1
X_11359_ _11359_/A _12647_/A vssd1 vssd1 vccd1 vccd1 _11359_/X sky130_fd_sc_hd__and2_1
XFILLER_152_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11590__C1 _11571_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18955_ _19508_/CLK _18955_/D vssd1 vssd1 vccd1 vccd1 _18955_/Q sky130_fd_sc_hd__dfxtp_1
X_14078_ _14146_/S vssd1 vssd1 vccd1 vccd1 _14087_/S sky130_fd_sc_hd__buf_2
XFILLER_141_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12134__A1 _12600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _16609_/B _12752_/X _12753_/X _17044_/B _13028_/X vssd1 vssd1 vccd1 vccd1
+ _13029_/X sky130_fd_sc_hd__a221o_1
X_17906_ _17906_/A vssd1 vssd1 vccd1 vccd1 _17906_/Y sky130_fd_sc_hd__clkinv_2
X_18886_ _19313_/CLK _18886_/D vssd1 vssd1 vccd1 vccd1 _18886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17837_ _17576_/X _17585_/X _17930_/S vssd1 vssd1 vccd1 vccd1 _17837_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14687__S _14691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16468__A _16939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10791__S1 _10037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17768_ _17772_/A _17772_/B vssd1 vssd1 vccd1 vccd1 _17768_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_75_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19507_ _19507_/CLK _19507_/D vssd1 vssd1 vccd1 vccd1 _19507_/Q sky130_fd_sc_hd__dfxtp_1
X_16719_ _19678_/Q _19677_/Q _19676_/Q _16719_/D vssd1 vssd1 vccd1 vccd1 _16729_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13604__B _13604_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17699_ _18009_/A vssd1 vssd1 vccd1 vccd1 _18109_/S sky130_fd_sc_hd__buf_2
X_19438_ _19470_/CLK _19438_/D vssd1 vssd1 vccd1 vccd1 _19438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11405__A _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19369_ _19369_/CLK _19369_/D vssd1 vssd1 vccd1 vccd1 _19369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16407__S _16415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17128__A2 _12026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18325__A1 _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16931__A _16946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__D_N _11585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10059__S0 _11451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17746__B _17749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09955_ _09955_/A vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09886_ _10233_/A _09885_/X _09696_/X vssd1 vssd1 vccd1 vccd1 _09886_/Y sky130_fd_sc_hd__o21ai_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10687__A1 _09979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16809__C _16809_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10730_ _10730_/A _10730_/B vssd1 vssd1 vccd1 vccd1 _10730_/X sky130_fd_sc_hd__or2_1
XFILLER_41_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19998__CLK _19998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13389__A0 _19914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ _19498_/Q _18910_/Q _18947_/Q _18521_/Q _10653_/X _10645_/X vssd1 vssd1 vccd1
+ vccd1 _10661_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _12314_/X _12398_/Y _12399_/X _12218_/X vssd1 vssd1 vccd1 vccd1 _12400_/Y
+ sky130_fd_sc_hd__o31ai_4
X_13380_ _19946_/Q vssd1 vssd1 vccd1 vccd1 _16317_/A sky130_fd_sc_hd__clkbuf_2
X_10592_ _10592_/A _10592_/B vssd1 vssd1 vccd1 vccd1 _10592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _12331_/A vssd1 vssd1 vccd1 vccd1 _17985_/B sky130_fd_sc_hd__buf_2
XANTENNA__09439__B _18324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17937__A _17937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11050__A _19899_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15050_ _15050_/A vssd1 vssd1 vccd1 vccd1 _19060_/D sky130_fd_sc_hd__clkbuf_1
X_12262_ _14477_/B vssd1 vssd1 vccd1 vccd1 _12262_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15550__A1 _15244_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14001_ _14151_/B _15301_/A vssd1 vssd1 vccd1 vccd1 _15918_/A sky130_fd_sc_hd__or2_2
XFILLER_107_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11213_ _19487_/Q _18899_/Q _18936_/Q _18510_/Q _10968_/S _10024_/A vssd1 vssd1 vccd1
+ vccd1 _11213_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16052__S _16056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12193_ _12272_/D vssd1 vssd1 vccd1 vccd1 _17933_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10375__B1 _09826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11144_ _11137_/Y _11139_/Y _11141_/Y _11143_/Y _10994_/X vssd1 vssd1 vccd1 vccd1
+ _11144_/X sky130_fd_sc_hd__o221a_4
Xoutput74 _12117_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[12] sky130_fd_sc_hd__buf_2
Xoutput85 _12391_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[22] sky130_fd_sc_hd__buf_2
XFILLER_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput96 _11816_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_150_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18740_ _19203_/CLK _18740_/D vssd1 vssd1 vccd1 vccd1 _18740_/Q sky130_fd_sc_hd__dfxtp_1
X_15952_ _15952_/A vssd1 vssd1 vccd1 vccd1 _19402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11075_ _11127_/A _11075_/B vssd1 vssd1 vccd1 vccd1 _11075_/X sky130_fd_sc_hd__or2_1
XANTENNA__10127__B1 _09693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14903_ _14656_/X _18995_/Q _14911_/S vssd1 vssd1 vccd1 vccd1 _14904_/A sky130_fd_sc_hd__mux2_1
X_10026_ _10041_/A vssd1 vssd1 vccd1 vccd1 _10665_/A sky130_fd_sc_hd__clkbuf_2
X_18671_ _19488_/CLK _18671_/D vssd1 vssd1 vccd1 vccd1 _18671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17391__B _17391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ _15883_/A vssd1 vssd1 vccd1 vccd1 _19371_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output131_A _12633_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ _11740_/A _17554_/B _09419_/X vssd1 vssd1 vccd1 vccd1 _17622_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13705__A _15270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14834_ _18359_/A _18403_/B vssd1 vssd1 vccd1 vccd1 _18966_/D sky130_fd_sc_hd__nor2_4
XFILLER_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14300__S _14308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17553_ _17516_/X _17521_/X _17552_/X _17966_/A vssd1 vssd1 vccd1 vccd1 _17554_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14765_ _14765_/A vssd1 vssd1 vccd1 vccd1 _18937_/D sky130_fd_sc_hd__clkbuf_1
X_11977_ _11977_/A vssd1 vssd1 vccd1 vccd1 _11977_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ _19671_/Q _19670_/Q _19672_/Q _16684_/A vssd1 vssd1 vccd1 vccd1 _16511_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__11225__A _11225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13716_ _13716_/A vssd1 vssd1 vccd1 vccd1 _18531_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15920__A _15988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17484_ _12257_/A _17937_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17484_/X sky130_fd_sc_hd__mux2_2
XFILLER_72_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10928_ _19460_/Q _19298_/Q _18707_/Q _18477_/Q _10040_/A _10910_/A vssd1 vssd1 vccd1
+ vccd1 _10929_/B sky130_fd_sc_hd__mux4_1
XFILLER_44_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14696_ _18902_/Q _14392_/X _14702_/S vssd1 vssd1 vccd1 vccd1 _14697_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19223_ _19481_/CLK _19223_/D vssd1 vssd1 vccd1 vccd1 _19223_/Q sky130_fd_sc_hd__dfxtp_1
X_16435_ _13506_/X _19574_/Q _16437_/S vssd1 vssd1 vccd1 vccd1 _16436_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13647_ _14602_/A vssd1 vssd1 vccd1 vccd1 _13647_/X sky130_fd_sc_hd__clkbuf_1
X_10859_ _19493_/Q _18905_/Q _18942_/Q _18516_/Q _10753_/S _10014_/A vssd1 vssd1 vccd1
+ vccd1 _10859_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15131__S _15131_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19154_ _19412_/CLK _19154_/D vssd1 vssd1 vccd1 vccd1 _19154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16318__A0 _15784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16366_/A vssd1 vssd1 vccd1 vccd1 _19544_/D sky130_fd_sc_hd__clkbuf_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13578_ _13578_/A vssd1 vssd1 vccd1 vccd1 _15818_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18105_ _18054_/X _17633_/Y _18104_/Y _18072_/X vssd1 vssd1 vccd1 vccd1 _18105_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15317_ _19168_/Q _15219_/X _15323_/S vssd1 vssd1 vccd1 vccd1 _15318_/A sky130_fd_sc_hd__mux2_1
X_19085_ _19564_/CLK _19085_/D vssd1 vssd1 vccd1 vccd1 _19085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12529_ _12529_/A vssd1 vssd1 vccd1 vccd1 _18090_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12056__A _12056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16297_ _19531_/Q _16296_/X _16325_/S vssd1 vssd1 vccd1 vccd1 _16298_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18036_ _18036_/A _18036_/B vssd1 vssd1 vccd1 vccd1 _18036_/Y sky130_fd_sc_hd__nor2_1
X_15248_ hold10/A vssd1 vssd1 vccd1 vccd1 _15261_/S sky130_fd_sc_hd__buf_2
XFILLER_160_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11158__A2 _11144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _19121_/Q vssd1 vssd1 vccd1 vccd1 _15180_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_113_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19987_ _19987_/CLK _19987_/D vssd1 vssd1 vccd1 vccd1 _19987_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12107__A1 _10727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _09740_/A vssd1 vssd1 vccd1 vccd1 _09741_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18938_ _19487_/CLK _18938_/D vssd1 vssd1 vccd1 vccd1 _18938_/Q sky130_fd_sc_hd__dfxtp_1
.ends

