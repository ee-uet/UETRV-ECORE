magic
tech sky130A
magscale 1 2
timestamp 1647604978
<< viali >>
rect 2697 17289 2731 17323
rect 7941 17289 7975 17323
rect 10333 17289 10367 17323
rect 14381 17289 14415 17323
rect 18245 17289 18279 17323
rect 3801 17221 3835 17255
rect 8401 17221 8435 17255
rect 2237 17153 2271 17187
rect 2513 17153 2547 17187
rect 6377 17153 6411 17187
rect 6745 17153 6779 17187
rect 6837 17153 6871 17187
rect 7389 17153 7423 17187
rect 8125 17153 8159 17187
rect 9137 17153 9171 17187
rect 10517 17153 10551 17187
rect 12265 17153 12299 17187
rect 12725 17153 12759 17187
rect 13185 17153 13219 17187
rect 14565 17153 14599 17187
rect 15025 17153 15059 17187
rect 15393 17153 15427 17187
rect 15669 17153 15703 17187
rect 16865 17153 16899 17187
rect 17509 17153 17543 17187
rect 18061 17153 18095 17187
rect 1961 17085 1995 17119
rect 9413 17085 9447 17119
rect 10793 17085 10827 17119
rect 12449 17085 12483 17119
rect 16313 17085 16347 17119
rect 6561 17017 6595 17051
rect 15853 17017 15887 17051
rect 17693 17017 17727 17051
rect 2973 16949 3007 16983
rect 7205 16949 7239 16983
rect 12081 16949 12115 16983
rect 14841 16949 14875 16983
rect 16681 16949 16715 16983
rect 2973 16745 3007 16779
rect 6009 16745 6043 16779
rect 8585 16745 8619 16779
rect 1869 16677 1903 16711
rect 3157 16677 3191 16711
rect 8125 16677 8159 16711
rect 11621 16677 11655 16711
rect 2421 16609 2455 16643
rect 7665 16609 7699 16643
rect 9137 16609 9171 16643
rect 11345 16609 11379 16643
rect 12357 16609 12391 16643
rect 14289 16609 14323 16643
rect 16589 16609 16623 16643
rect 4914 16541 4948 16575
rect 5181 16541 5215 16575
rect 5641 16541 5675 16575
rect 7389 16541 7423 16575
rect 7757 16541 7791 16575
rect 7941 16541 7975 16575
rect 11253 16541 11287 16575
rect 11897 16541 11931 16575
rect 14556 16541 14590 16575
rect 16845 16541 16879 16575
rect 1685 16473 1719 16507
rect 2237 16473 2271 16507
rect 3433 16473 3467 16507
rect 7144 16473 7178 16507
rect 9404 16473 9438 16507
rect 12602 16473 12636 16507
rect 15945 16473 15979 16507
rect 16129 16473 16163 16507
rect 3801 16405 3835 16439
rect 5457 16405 5491 16439
rect 10517 16405 10551 16439
rect 12081 16405 12115 16439
rect 13737 16405 13771 16439
rect 15669 16405 15703 16439
rect 16313 16405 16347 16439
rect 17969 16405 18003 16439
rect 1961 16201 1995 16235
rect 2237 16201 2271 16235
rect 3525 16201 3559 16235
rect 3709 16201 3743 16235
rect 6377 16201 6411 16235
rect 9413 16201 9447 16235
rect 10241 16201 10275 16235
rect 10609 16201 10643 16235
rect 14841 16201 14875 16235
rect 15685 16201 15719 16235
rect 15853 16201 15887 16235
rect 17049 16201 17083 16235
rect 3617 16133 3651 16167
rect 3893 16133 3927 16167
rect 6561 16133 6595 16167
rect 10793 16133 10827 16167
rect 13001 16133 13035 16167
rect 13613 16133 13647 16167
rect 13829 16133 13863 16167
rect 14657 16133 14691 16167
rect 15485 16133 15519 16167
rect 16681 16133 16715 16167
rect 16897 16133 16931 16167
rect 17417 16133 17451 16167
rect 1409 16065 1443 16099
rect 2789 16065 2823 16099
rect 2973 16065 3007 16099
rect 3065 16065 3099 16099
rect 4445 16065 4479 16099
rect 5549 16065 5583 16099
rect 5641 16065 5675 16099
rect 6929 16065 6963 16099
rect 7205 16065 7239 16099
rect 7389 16065 7423 16099
rect 7757 16065 7791 16099
rect 8024 16065 8058 16099
rect 9597 16065 9631 16099
rect 10057 16065 10091 16099
rect 10333 16065 10367 16099
rect 11529 16065 11563 16099
rect 14289 16065 14323 16099
rect 16313 16065 16347 16099
rect 17325 16065 17359 16099
rect 17509 16065 17543 16099
rect 4169 15997 4203 16031
rect 5365 15997 5399 16031
rect 5457 15997 5491 16031
rect 9873 15997 9907 16031
rect 11805 15997 11839 16031
rect 17785 15997 17819 16031
rect 2789 15929 2823 15963
rect 3341 15929 3375 15963
rect 5825 15929 5859 15963
rect 9137 15929 9171 15963
rect 11161 15929 11195 15963
rect 12633 15929 12667 15963
rect 13461 15929 13495 15963
rect 16129 15929 16163 15963
rect 6561 15861 6595 15895
rect 7389 15861 7423 15895
rect 10793 15861 10827 15895
rect 13001 15861 13035 15895
rect 13185 15861 13219 15895
rect 13645 15861 13679 15895
rect 14657 15861 14691 15895
rect 15669 15861 15703 15895
rect 16865 15861 16899 15895
rect 3249 15657 3283 15691
rect 3341 15657 3375 15691
rect 6653 15657 6687 15691
rect 10885 15657 10919 15691
rect 12357 15657 12391 15691
rect 15209 15657 15243 15691
rect 18337 15657 18371 15691
rect 2881 15589 2915 15623
rect 7389 15589 7423 15623
rect 11253 15589 11287 15623
rect 14335 15589 14369 15623
rect 3157 15521 3191 15555
rect 3801 15521 3835 15555
rect 4077 15521 4111 15555
rect 5273 15521 5307 15555
rect 11713 15521 11747 15555
rect 16957 15521 16991 15555
rect 1501 15453 1535 15487
rect 3433 15453 3467 15487
rect 5540 15453 5574 15487
rect 7113 15453 7147 15487
rect 7389 15453 7423 15487
rect 7665 15453 7699 15487
rect 8033 15453 8067 15487
rect 9505 15453 9539 15487
rect 9781 15453 9815 15487
rect 10057 15453 10091 15487
rect 10241 15453 10275 15487
rect 10333 15453 10367 15487
rect 11621 15453 11655 15487
rect 12081 15453 12115 15487
rect 12817 15453 12851 15487
rect 13645 15453 13679 15487
rect 14105 15453 14139 15487
rect 15393 15453 15427 15487
rect 15669 15453 15703 15487
rect 16129 15453 16163 15487
rect 1768 15385 1802 15419
rect 7941 15385 7975 15419
rect 11897 15385 11931 15419
rect 13001 15385 13035 15419
rect 13185 15385 13219 15419
rect 16313 15385 16347 15419
rect 17224 15385 17258 15419
rect 7205 15317 7239 15351
rect 7849 15317 7883 15351
rect 8217 15317 8251 15351
rect 10701 15317 10735 15351
rect 10885 15317 10919 15351
rect 11989 15317 12023 15351
rect 12633 15317 12667 15351
rect 12909 15317 12943 15351
rect 13461 15317 13495 15351
rect 15577 15317 15611 15351
rect 16497 15317 16531 15351
rect 4077 15113 4111 15147
rect 4261 15113 4295 15147
rect 7941 15113 7975 15147
rect 11713 15113 11747 15147
rect 12725 15113 12759 15147
rect 14565 15113 14599 15147
rect 15669 15113 15703 15147
rect 17049 15113 17083 15147
rect 17325 15113 17359 15147
rect 5733 15045 5767 15079
rect 10793 15045 10827 15079
rect 12357 15045 12391 15079
rect 12541 15045 12575 15079
rect 13452 15045 13486 15079
rect 15025 15045 15059 15079
rect 15393 15045 15427 15079
rect 15945 15045 15979 15079
rect 16681 15045 16715 15079
rect 16881 15045 16915 15079
rect 1409 14977 1443 15011
rect 2136 14977 2170 15011
rect 4537 14977 4571 15011
rect 4721 14977 4755 15011
rect 4997 14977 5031 15011
rect 5365 14977 5399 15011
rect 6745 14977 6779 15011
rect 6929 14977 6963 15011
rect 7389 14977 7423 15011
rect 7849 14977 7883 15011
rect 7941 14977 7975 15011
rect 8493 14977 8527 15011
rect 8677 14977 8711 15011
rect 8769 14977 8803 15011
rect 8861 14977 8895 15011
rect 9413 14977 9447 15011
rect 10517 14977 10551 15011
rect 10885 14977 10919 15011
rect 12081 14977 12115 15011
rect 15301 14977 15335 15011
rect 15669 14977 15703 15011
rect 17509 14977 17543 15011
rect 18337 14977 18371 15011
rect 1869 14909 1903 14943
rect 3709 14909 3743 14943
rect 5457 14909 5491 14943
rect 5549 14909 5583 14943
rect 7665 14909 7699 14943
rect 9689 14909 9723 14943
rect 10701 14909 10735 14943
rect 13185 14909 13219 14943
rect 15761 14909 15795 14943
rect 3249 14841 3283 14875
rect 9137 14841 9171 14875
rect 15025 14841 15059 14875
rect 15209 14841 15243 14875
rect 4077 14773 4111 14807
rect 4905 14773 4939 14807
rect 6837 14773 6871 14807
rect 7297 14773 7331 14807
rect 10517 14773 10551 14807
rect 11529 14773 11563 14807
rect 11713 14773 11747 14807
rect 16865 14773 16899 14807
rect 3985 14569 4019 14603
rect 5365 14569 5399 14603
rect 6285 14569 6319 14603
rect 6469 14569 6503 14603
rect 10057 14569 10091 14603
rect 10977 14569 11011 14603
rect 11805 14569 11839 14603
rect 16221 14569 16255 14603
rect 17877 14569 17911 14603
rect 7021 14501 7055 14535
rect 8953 14501 8987 14535
rect 14105 14501 14139 14535
rect 3801 14433 3835 14467
rect 7482 14433 7516 14467
rect 7573 14433 7607 14467
rect 9137 14433 9171 14467
rect 14749 14433 14783 14467
rect 16589 14433 16623 14467
rect 1409 14365 1443 14399
rect 4261 14365 4295 14399
rect 5641 14365 5675 14399
rect 5917 14365 5951 14399
rect 6745 14365 6779 14399
rect 7021 14365 7055 14399
rect 7665 14365 7699 14399
rect 7758 14365 7792 14399
rect 9229 14365 9263 14399
rect 11621 14365 11655 14399
rect 12725 14365 12759 14399
rect 12909 14365 12943 14399
rect 13001 14365 13035 14399
rect 13093 14365 13127 14399
rect 14565 14365 14599 14399
rect 15117 14365 15151 14399
rect 15301 14365 15335 14399
rect 15761 14365 15795 14399
rect 16129 14365 16163 14399
rect 16313 14365 16347 14399
rect 18337 14365 18371 14399
rect 4169 14297 4203 14331
rect 4997 14297 5031 14331
rect 5411 14297 5445 14331
rect 6929 14297 6963 14331
rect 8309 14297 8343 14331
rect 8493 14297 8527 14331
rect 9873 14297 9907 14331
rect 10089 14297 10123 14331
rect 11161 14297 11195 14331
rect 11345 14297 11379 14331
rect 6285 14229 6319 14263
rect 7297 14229 7331 14263
rect 8125 14229 8159 14263
rect 9597 14229 9631 14263
rect 10241 14229 10275 14263
rect 13369 14229 13403 14263
rect 14473 14229 14507 14263
rect 15301 14229 15335 14263
rect 15577 14229 15611 14263
rect 5825 14025 5859 14059
rect 9531 14025 9565 14059
rect 9965 14025 9999 14059
rect 14749 14025 14783 14059
rect 18061 14025 18095 14059
rect 6621 13957 6655 13991
rect 6837 13957 6871 13991
rect 9321 13957 9355 13991
rect 10885 13957 10919 13991
rect 12992 13957 13026 13991
rect 3341 13889 3375 13923
rect 3608 13889 3642 13923
rect 5273 13889 5307 13923
rect 5641 13889 5675 13923
rect 7573 13889 7607 13923
rect 7757 13889 7791 13923
rect 7849 13889 7883 13923
rect 8677 13889 8711 13923
rect 8769 13889 8803 13923
rect 8953 13889 8987 13923
rect 9045 13889 9079 13923
rect 9965 13889 9999 13923
rect 10149 13889 10183 13923
rect 12081 13889 12115 13923
rect 12173 13889 12207 13923
rect 12265 13889 12299 13923
rect 12449 13889 12483 13923
rect 12725 13889 12759 13923
rect 15862 13889 15896 13923
rect 16129 13889 16163 13923
rect 16681 13889 16715 13923
rect 16937 13889 16971 13923
rect 7113 13821 7147 13855
rect 10701 13753 10735 13787
rect 4721 13685 4755 13719
rect 5549 13685 5583 13719
rect 6469 13685 6503 13719
rect 6653 13685 6687 13719
rect 8493 13685 8527 13719
rect 9505 13685 9539 13719
rect 9689 13685 9723 13719
rect 11805 13685 11839 13719
rect 14105 13685 14139 13719
rect 3801 13481 3835 13515
rect 5273 13481 5307 13515
rect 5733 13481 5767 13515
rect 6101 13481 6135 13515
rect 7021 13481 7055 13515
rect 8217 13481 8251 13515
rect 9137 13481 9171 13515
rect 18337 13481 18371 13515
rect 4905 13413 4939 13447
rect 8401 13413 8435 13447
rect 11253 13413 11287 13447
rect 13185 13413 13219 13447
rect 15301 13345 15335 13379
rect 15485 13345 15519 13379
rect 16497 13345 16531 13379
rect 16957 13345 16991 13379
rect 2053 13277 2087 13311
rect 3985 13277 4019 13311
rect 4261 13277 4295 13311
rect 4721 13277 4755 13311
rect 5365 13277 5399 13311
rect 5457 13277 5491 13311
rect 5733 13277 5767 13311
rect 5825 13277 5859 13311
rect 7849 13277 7883 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 9873 13277 9907 13311
rect 11529 13277 11563 13311
rect 16405 13277 16439 13311
rect 2320 13209 2354 13243
rect 5181 13209 5215 13243
rect 7205 13209 7239 13243
rect 8217 13209 8251 13243
rect 10140 13209 10174 13243
rect 11796 13209 11830 13243
rect 13369 13209 13403 13243
rect 14381 13209 14415 13243
rect 15209 13209 15243 13243
rect 17202 13209 17236 13243
rect 3433 13141 3467 13175
rect 4445 13141 4479 13175
rect 6837 13141 6871 13175
rect 7005 13141 7039 13175
rect 12909 13141 12943 13175
rect 14473 13141 14507 13175
rect 14841 13141 14875 13175
rect 15945 13141 15979 13175
rect 16313 13141 16347 13175
rect 2605 12937 2639 12971
rect 4353 12937 4387 12971
rect 5825 12937 5859 12971
rect 10425 12937 10459 12971
rect 11897 12937 11931 12971
rect 13185 12937 13219 12971
rect 15209 12937 15243 12971
rect 16313 12937 16347 12971
rect 17141 12937 17175 12971
rect 18245 12937 18279 12971
rect 4445 12869 4479 12903
rect 9873 12869 9907 12903
rect 13093 12869 13127 12903
rect 2237 12801 2271 12835
rect 2789 12801 2823 12835
rect 3249 12801 3283 12835
rect 4813 12801 4847 12835
rect 4997 12801 5031 12835
rect 6561 12801 6595 12835
rect 7950 12801 7984 12835
rect 8217 12801 8251 12835
rect 9321 12801 9355 12835
rect 9689 12801 9723 12835
rect 10701 12801 10735 12835
rect 10793 12801 10827 12835
rect 10885 12801 10919 12835
rect 11069 12801 11103 12835
rect 11989 12801 12023 12835
rect 14565 12801 14599 12835
rect 14749 12801 14783 12835
rect 14841 12801 14875 12835
rect 14933 12801 14967 12835
rect 15669 12801 15703 12835
rect 15832 12804 15866 12838
rect 15964 12804 15998 12838
rect 16057 12801 16091 12835
rect 17049 12801 17083 12835
rect 18061 12801 18095 12835
rect 5181 12733 5215 12767
rect 5641 12733 5675 12767
rect 6009 12733 6043 12767
rect 9045 12733 9079 12767
rect 12173 12733 12207 12767
rect 13369 12733 13403 12767
rect 17233 12733 17267 12767
rect 6377 12665 6411 12699
rect 6837 12665 6871 12699
rect 11529 12665 11563 12699
rect 12725 12665 12759 12699
rect 2053 12597 2087 12631
rect 3065 12597 3099 12631
rect 5457 12597 5491 12631
rect 16681 12597 16715 12631
rect 4813 12393 4847 12427
rect 5733 12393 5767 12427
rect 6285 12393 6319 12427
rect 7205 12393 7239 12427
rect 7665 12393 7699 12427
rect 10609 12393 10643 12427
rect 11897 12393 11931 12427
rect 14749 12393 14783 12427
rect 15393 12393 15427 12427
rect 18337 12393 18371 12427
rect 11253 12325 11287 12359
rect 5733 12257 5767 12291
rect 7021 12257 7055 12291
rect 8953 12257 8987 12291
rect 9229 12257 9263 12291
rect 12449 12257 12483 12291
rect 1685 12189 1719 12223
rect 1952 12189 1986 12223
rect 4261 12189 4295 12223
rect 4353 12189 4387 12223
rect 4997 12189 5031 12223
rect 5181 12189 5215 12223
rect 5457 12189 5491 12223
rect 6469 12189 6503 12223
rect 6837 12189 6871 12223
rect 7205 12189 7239 12223
rect 10885 12189 10919 12223
rect 11529 12189 11563 12223
rect 12173 12189 12207 12223
rect 13461 12189 13495 12223
rect 13737 12189 13771 12223
rect 15025 12189 15059 12223
rect 16037 12189 16071 12223
rect 16221 12189 16255 12223
rect 16313 12189 16347 12223
rect 16405 12189 16439 12223
rect 16957 12189 16991 12223
rect 4537 12121 4571 12155
rect 7573 12121 7607 12155
rect 10241 12121 10275 12155
rect 10425 12121 10459 12155
rect 11069 12121 11103 12155
rect 11713 12121 11747 12155
rect 14381 12121 14415 12155
rect 14565 12121 14599 12155
rect 15209 12121 15243 12155
rect 16681 12121 16715 12155
rect 17202 12121 17236 12155
rect 3065 12053 3099 12087
rect 6009 12053 6043 12087
rect 6929 12053 6963 12087
rect 13277 12053 13311 12087
rect 13645 12053 13679 12087
rect 5733 11849 5767 11883
rect 8769 11849 8803 11883
rect 2136 11781 2170 11815
rect 4068 11781 4102 11815
rect 7021 11781 7055 11815
rect 7656 11781 7690 11815
rect 13452 11781 13486 11815
rect 16313 11781 16347 11815
rect 17018 11781 17052 11815
rect 1869 11713 1903 11747
rect 5825 11713 5859 11747
rect 6745 11713 6779 11747
rect 7389 11713 7423 11747
rect 9045 11713 9079 11747
rect 9312 11713 9346 11747
rect 10701 11713 10735 11747
rect 10885 11713 10919 11747
rect 11785 11713 11819 11747
rect 15025 11713 15059 11747
rect 15209 11713 15243 11747
rect 15669 11713 15703 11747
rect 15853 11713 15887 11747
rect 15945 11713 15979 11747
rect 16037 11713 16071 11747
rect 3801 11645 3835 11679
rect 6837 11645 6871 11679
rect 7021 11645 7055 11679
rect 11529 11645 11563 11679
rect 13185 11645 13219 11679
rect 15393 11645 15427 11679
rect 16773 11645 16807 11679
rect 1409 11577 1443 11611
rect 3249 11509 3283 11543
rect 5181 11509 5215 11543
rect 10425 11509 10459 11543
rect 11069 11509 11103 11543
rect 12909 11509 12943 11543
rect 14565 11509 14599 11543
rect 18153 11509 18187 11543
rect 3985 11305 4019 11339
rect 4629 11305 4663 11339
rect 6009 11305 6043 11339
rect 8585 11305 8619 11339
rect 10977 11305 11011 11339
rect 12173 11305 12207 11339
rect 16129 11305 16163 11339
rect 3433 11237 3467 11271
rect 5181 11237 5215 11271
rect 5273 11237 5307 11271
rect 7757 11237 7791 11271
rect 9597 11237 9631 11271
rect 15853 11237 15887 11271
rect 2605 11169 2639 11203
rect 10241 11169 10275 11203
rect 12725 11169 12759 11203
rect 16681 11169 16715 11203
rect 1409 11101 1443 11135
rect 2421 11101 2455 11135
rect 3249 11101 3283 11135
rect 4537 11101 4571 11135
rect 5273 11101 5307 11135
rect 5549 11101 5583 11135
rect 5733 11101 5767 11135
rect 7389 11101 7423 11135
rect 7849 11101 7883 11135
rect 8401 11101 8435 11135
rect 8953 11101 8987 11135
rect 9137 11101 9171 11135
rect 9321 11101 9355 11135
rect 9965 11101 9999 11135
rect 10793 11101 10827 11135
rect 12541 11101 12575 11135
rect 16589 11101 16623 11135
rect 17877 11101 17911 11135
rect 18337 11101 18371 11135
rect 3801 11033 3835 11067
rect 4017 11033 4051 11067
rect 4997 11033 5031 11067
rect 5641 11033 5675 11067
rect 7144 11033 7178 11067
rect 10057 11033 10091 11067
rect 11345 11033 11379 11067
rect 12633 11033 12667 11067
rect 13277 11033 13311 11067
rect 13461 11033 13495 11067
rect 14749 11033 14783 11067
rect 14933 11033 14967 11067
rect 15485 11033 15519 11067
rect 15669 11033 15703 11067
rect 16497 11033 16531 11067
rect 17509 11033 17543 11067
rect 2237 10965 2271 10999
rect 4169 10965 4203 10999
rect 11437 10965 11471 10999
rect 18153 10965 18187 10999
rect 5733 10761 5767 10795
rect 9781 10761 9815 10795
rect 16129 10761 16163 10795
rect 6929 10693 6963 10727
rect 7573 10693 7607 10727
rect 10977 10693 11011 10727
rect 11989 10693 12023 10727
rect 16037 10693 16071 10727
rect 1777 10625 1811 10659
rect 2044 10625 2078 10659
rect 3893 10625 3927 10659
rect 4160 10625 4194 10659
rect 5641 10625 5675 10659
rect 7297 10625 7331 10659
rect 7389 10625 7423 10659
rect 7849 10625 7883 10659
rect 8033 10625 8067 10659
rect 9689 10625 9723 10659
rect 10609 10625 10643 10659
rect 11897 10625 11931 10659
rect 12173 10625 12207 10659
rect 12817 10625 12851 10659
rect 13001 10625 13035 10659
rect 13093 10625 13127 10659
rect 13185 10625 13219 10659
rect 14289 10625 14323 10659
rect 14556 10625 14590 10659
rect 16681 10625 16715 10659
rect 16948 10625 16982 10659
rect 9873 10557 9907 10591
rect 13461 10557 13495 10591
rect 6745 10489 6779 10523
rect 7573 10489 7607 10523
rect 11161 10489 11195 10523
rect 15669 10489 15703 10523
rect 3157 10421 3191 10455
rect 5273 10421 5307 10455
rect 7849 10421 7883 10455
rect 9321 10421 9355 10455
rect 10425 10421 10459 10455
rect 12173 10421 12207 10455
rect 14013 10421 14047 10455
rect 18061 10421 18095 10455
rect 2145 10217 2179 10251
rect 2697 10217 2731 10251
rect 5365 10217 5399 10251
rect 18337 10217 18371 10251
rect 7941 10149 7975 10183
rect 3341 10081 3375 10115
rect 3985 10081 4019 10115
rect 10517 10081 10551 10115
rect 12265 10081 12299 10115
rect 16129 10081 16163 10115
rect 16957 10081 16991 10115
rect 1409 10013 1443 10047
rect 2329 10013 2363 10047
rect 3065 10013 3099 10047
rect 4169 10013 4203 10047
rect 4537 10013 4571 10047
rect 5457 10013 5491 10047
rect 6009 10013 6043 10047
rect 6285 10013 6319 10047
rect 8125 10013 8159 10047
rect 10261 10013 10295 10047
rect 11345 10013 11379 10047
rect 11529 10013 11563 10047
rect 11805 10013 11839 10047
rect 15485 10013 15519 10047
rect 16313 10013 16347 10047
rect 3157 9945 3191 9979
rect 6552 9945 6586 9979
rect 8585 9945 8619 9979
rect 10977 9945 11011 9979
rect 12510 9945 12544 9979
rect 15218 9945 15252 9979
rect 17224 9945 17258 9979
rect 4721 9877 4755 9911
rect 5825 9877 5859 9911
rect 7665 9877 7699 9911
rect 9137 9877 9171 9911
rect 10885 9877 10919 9911
rect 11989 9877 12023 9911
rect 13645 9877 13679 9911
rect 14105 9877 14139 9911
rect 16221 9877 16255 9911
rect 16681 9877 16715 9911
rect 6837 9673 6871 9707
rect 14657 9673 14691 9707
rect 17325 9673 17359 9707
rect 4353 9605 4387 9639
rect 12642 9605 12676 9639
rect 18245 9605 18279 9639
rect 2145 9537 2179 9571
rect 2329 9537 2363 9571
rect 2513 9537 2547 9571
rect 2973 9537 3007 9571
rect 4169 9537 4203 9571
rect 5742 9537 5776 9571
rect 6009 9537 6043 9571
rect 7021 9537 7055 9571
rect 7113 9537 7147 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 7665 9537 7699 9571
rect 7932 9537 7966 9571
rect 9321 9537 9355 9571
rect 13185 9537 13219 9571
rect 13645 9537 13679 9571
rect 13829 9537 13863 9571
rect 14013 9537 14047 9571
rect 14289 9537 14323 9571
rect 14841 9537 14875 9571
rect 15577 9537 15611 9571
rect 15761 9537 15795 9571
rect 16129 9537 16163 9571
rect 16681 9537 16715 9571
rect 16865 9537 16899 9571
rect 17509 9537 17543 9571
rect 18061 9537 18095 9571
rect 3985 9469 4019 9503
rect 12909 9469 12943 9503
rect 15117 9469 15151 9503
rect 15393 9469 15427 9503
rect 17049 9469 17083 9503
rect 17785 9469 17819 9503
rect 13369 9401 13403 9435
rect 16313 9401 16347 9435
rect 2789 9333 2823 9367
rect 4629 9333 4663 9367
rect 9045 9333 9079 9367
rect 10609 9333 10643 9367
rect 11529 9333 11563 9367
rect 15025 9333 15059 9367
rect 17693 9333 17727 9367
rect 4077 9129 4111 9163
rect 7941 9129 7975 9163
rect 9137 9129 9171 9163
rect 9965 9129 9999 9163
rect 10977 9129 11011 9163
rect 11529 9129 11563 9163
rect 12265 9129 12299 9163
rect 14105 9129 14139 9163
rect 15853 9129 15887 9163
rect 17785 9129 17819 9163
rect 6561 9061 6595 9095
rect 4721 8993 4755 9027
rect 5089 8993 5123 9027
rect 11069 8993 11103 9027
rect 11667 8993 11701 9027
rect 14749 8993 14783 9027
rect 16221 8993 16255 9027
rect 1593 8925 1627 8959
rect 1860 8925 1894 8959
rect 3249 8925 3283 8959
rect 6101 8925 6135 8959
rect 6745 8925 6779 8959
rect 7573 8925 7607 8959
rect 8125 8925 8159 8959
rect 8309 8925 8343 8959
rect 8401 8925 8435 8959
rect 9597 8925 9631 8959
rect 9781 8925 9815 8959
rect 10793 8925 10827 8959
rect 11345 8925 11379 8959
rect 11805 8925 11839 8959
rect 12081 8925 12115 8959
rect 12265 8925 12299 8959
rect 12817 8925 12851 8959
rect 13001 8925 13035 8959
rect 13185 8925 13219 8959
rect 15577 8925 15611 8959
rect 16405 8925 16439 8959
rect 16589 8925 16623 8959
rect 16865 8925 16899 8959
rect 17509 8925 17543 8959
rect 17969 8925 18003 8959
rect 18061 8925 18095 8959
rect 4537 8857 4571 8891
rect 5273 8857 5307 8891
rect 9321 8857 9355 8891
rect 11437 8857 11471 8891
rect 13093 8857 13127 8891
rect 13737 8857 13771 8891
rect 2973 8789 3007 8823
rect 3433 8789 3467 8823
rect 4445 8789 4479 8823
rect 6285 8789 6319 8823
rect 7573 8789 7607 8823
rect 8953 8789 8987 8823
rect 9121 8789 9155 8823
rect 10609 8789 10643 8823
rect 13369 8789 13403 8823
rect 14473 8789 14507 8823
rect 14565 8789 14599 8823
rect 15393 8789 15427 8823
rect 17049 8789 17083 8823
rect 1501 8585 1535 8619
rect 2513 8585 2547 8619
rect 2881 8585 2915 8619
rect 5181 8585 5215 8619
rect 5457 8585 5491 8619
rect 7757 8585 7791 8619
rect 8861 8585 8895 8619
rect 11621 8585 11655 8619
rect 4046 8517 4080 8551
rect 8401 8517 8435 8551
rect 10802 8517 10836 8551
rect 17040 8517 17074 8551
rect 1685 8449 1719 8483
rect 2053 8449 2087 8483
rect 2145 8449 2179 8483
rect 5641 8449 5675 8483
rect 5733 8449 5767 8483
rect 6377 8449 6411 8483
rect 6633 8449 6667 8483
rect 8217 8449 8251 8483
rect 9045 8449 9079 8483
rect 9137 8449 9171 8483
rect 11805 8449 11839 8483
rect 12081 8449 12115 8483
rect 12260 8449 12294 8483
rect 12360 8452 12394 8486
rect 12495 8449 12529 8483
rect 13001 8449 13035 8483
rect 13185 8449 13219 8483
rect 13277 8449 13311 8483
rect 13369 8449 13403 8483
rect 13921 8449 13955 8483
rect 14105 8449 14139 8483
rect 14289 8449 14323 8483
rect 14473 8449 14507 8483
rect 14933 8449 14967 8483
rect 15189 8449 15223 8483
rect 16773 8449 16807 8483
rect 2973 8381 3007 8415
rect 3157 8381 3191 8415
rect 3801 8381 3835 8415
rect 9229 8381 9263 8415
rect 9321 8381 9355 8415
rect 11069 8381 11103 8415
rect 14197 8381 14231 8415
rect 14657 8381 14691 8415
rect 8585 8313 8619 8347
rect 12725 8313 12759 8347
rect 13645 8313 13679 8347
rect 9689 8245 9723 8279
rect 16313 8245 16347 8279
rect 18153 8245 18187 8279
rect 4629 8041 4663 8075
rect 6469 8041 6503 8075
rect 11805 8041 11839 8075
rect 13185 8041 13219 8075
rect 14105 8041 14139 8075
rect 15209 8041 15243 8075
rect 16313 8041 16347 8075
rect 7389 7973 7423 8007
rect 3065 7905 3099 7939
rect 4077 7905 4111 7939
rect 7849 7905 7883 7939
rect 8033 7905 8067 7939
rect 9229 7905 9263 7939
rect 13737 7905 13771 7939
rect 16865 7905 16899 7939
rect 17509 7905 17543 7939
rect 2145 7837 2179 7871
rect 2789 7837 2823 7871
rect 4169 7837 4203 7871
rect 4261 7837 4295 7871
rect 6101 7837 6135 7871
rect 6653 7837 6687 7871
rect 6745 7837 6779 7871
rect 8953 7837 8987 7871
rect 10425 7837 10459 7871
rect 10701 7837 10735 7871
rect 10793 7837 10827 7871
rect 11253 7837 11287 7871
rect 11989 7837 12023 7871
rect 12081 7837 12115 7871
rect 12173 7837 12207 7871
rect 12357 7837 12391 7871
rect 12633 7837 12667 7871
rect 12725 7837 12759 7871
rect 12909 7837 12943 7871
rect 13001 7837 13035 7871
rect 13553 7837 13587 7871
rect 14284 7837 14318 7871
rect 14473 7837 14507 7871
rect 14656 7837 14690 7871
rect 14749 7837 14783 7871
rect 15117 7837 15151 7871
rect 16037 7837 16071 7871
rect 16681 7837 16715 7871
rect 17785 7837 17819 7871
rect 5917 7769 5951 7803
rect 7757 7769 7791 7803
rect 10609 7769 10643 7803
rect 14381 7769 14415 7803
rect 1961 7701 1995 7735
rect 2421 7701 2455 7735
rect 2881 7701 2915 7735
rect 10977 7701 11011 7735
rect 11437 7701 11471 7735
rect 16773 7701 16807 7735
rect 7481 7497 7515 7531
rect 9689 7497 9723 7531
rect 1952 7429 1986 7463
rect 6837 7429 6871 7463
rect 7849 7429 7883 7463
rect 8065 7429 8099 7463
rect 13645 7429 13679 7463
rect 14841 7429 14875 7463
rect 15393 7429 15427 7463
rect 17202 7429 17236 7463
rect 1685 7361 1719 7395
rect 4445 7361 4479 7395
rect 4905 7361 4939 7395
rect 5365 7361 5399 7395
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 7573 7361 7607 7395
rect 8493 7361 8527 7395
rect 9781 7361 9815 7395
rect 10701 7361 10735 7395
rect 10793 7361 10827 7395
rect 10977 7361 11011 7395
rect 11069 7361 11103 7395
rect 11529 7361 11563 7395
rect 12725 7361 12759 7395
rect 13553 7361 13587 7395
rect 13737 7361 13771 7395
rect 13921 7361 13955 7395
rect 14197 7361 14231 7395
rect 14360 7361 14394 7395
rect 14473 7361 14507 7395
rect 14611 7361 14645 7395
rect 15117 7361 15151 7395
rect 15301 7361 15335 7395
rect 15485 7361 15519 7395
rect 16129 7361 16163 7395
rect 16957 7361 16991 7395
rect 4169 7293 4203 7327
rect 4721 7293 4755 7327
rect 8769 7293 8803 7327
rect 11805 7293 11839 7327
rect 16313 7293 16347 7327
rect 5089 7225 5123 7259
rect 6653 7225 6687 7259
rect 8217 7225 8251 7259
rect 12909 7225 12943 7259
rect 3065 7157 3099 7191
rect 5549 7157 5583 7191
rect 8033 7157 8067 7191
rect 10517 7157 10551 7191
rect 13369 7157 13403 7191
rect 15669 7157 15703 7191
rect 15945 7157 15979 7191
rect 18337 7157 18371 7191
rect 1961 6953 1995 6987
rect 4905 6953 4939 6987
rect 8125 6953 8159 6987
rect 8953 6953 8987 6987
rect 14933 6953 14967 6987
rect 16313 6953 16347 6987
rect 12265 6885 12299 6919
rect 1409 6817 1443 6851
rect 2329 6817 2363 6851
rect 3065 6817 3099 6851
rect 4353 6817 4387 6851
rect 6561 6817 6595 6851
rect 9229 6817 9263 6851
rect 12357 6817 12391 6851
rect 12541 6817 12575 6851
rect 12817 6817 12851 6851
rect 16773 6817 16807 6851
rect 16865 6817 16899 6851
rect 17877 6817 17911 6851
rect 2145 6749 2179 6783
rect 2789 6749 2823 6783
rect 3249 6749 3283 6783
rect 6294 6749 6328 6783
rect 7757 6749 7791 6783
rect 9597 6749 9631 6783
rect 9873 6749 9907 6783
rect 10057 6749 10091 6783
rect 10241 6749 10275 6783
rect 10425 6749 10459 6783
rect 11437 6749 11471 6783
rect 11805 6749 11839 6783
rect 12265 6749 12299 6783
rect 13093 6749 13127 6783
rect 14125 6749 14159 6783
rect 14473 6749 14507 6783
rect 15117 6749 15151 6783
rect 15209 6749 15243 6783
rect 15393 6749 15427 6783
rect 15485 6749 15519 6783
rect 15853 6749 15887 6783
rect 17693 6749 17727 6783
rect 3433 6681 3467 6715
rect 9112 6681 9146 6715
rect 10793 6681 10827 6715
rect 11621 6681 11655 6715
rect 11713 6681 11747 6715
rect 14289 6681 14323 6715
rect 14381 6681 14415 6715
rect 17785 6681 17819 6715
rect 2605 6613 2639 6647
rect 4445 6613 4479 6647
rect 4537 6613 4571 6647
rect 5181 6613 5215 6647
rect 8125 6613 8159 6647
rect 8309 6613 8343 6647
rect 9321 6613 9355 6647
rect 10149 6613 10183 6647
rect 10885 6613 10919 6647
rect 11989 6613 12023 6647
rect 14657 6613 14691 6647
rect 16037 6613 16071 6647
rect 16681 6613 16715 6647
rect 17325 6613 17359 6647
rect 2881 6409 2915 6443
rect 4169 6409 4203 6443
rect 4537 6409 4571 6443
rect 6837 6409 6871 6443
rect 7573 6409 7607 6443
rect 9413 6409 9447 6443
rect 10333 6409 10367 6443
rect 11161 6409 11195 6443
rect 15669 6409 15703 6443
rect 18245 6409 18279 6443
rect 2973 6341 3007 6375
rect 4629 6341 4663 6375
rect 5365 6341 5399 6375
rect 6745 6341 6779 6375
rect 7205 6341 7239 6375
rect 7421 6341 7455 6375
rect 8401 6341 8435 6375
rect 8953 6341 8987 6375
rect 9229 6341 9263 6375
rect 13185 6341 13219 6375
rect 13921 6341 13955 6375
rect 14013 6341 14047 6375
rect 17110 6341 17144 6375
rect 1685 6273 1719 6307
rect 3709 6273 3743 6307
rect 5917 6273 5951 6307
rect 7941 6273 7975 6307
rect 8125 6273 8159 6307
rect 8677 6273 8711 6307
rect 10980 6273 11014 6307
rect 11713 6273 11747 6307
rect 11805 6273 11839 6307
rect 11989 6273 12023 6307
rect 12081 6273 12115 6307
rect 12449 6273 12483 6307
rect 12909 6273 12943 6307
rect 13093 6273 13127 6307
rect 13277 6273 13311 6307
rect 13737 6273 13771 6307
rect 14105 6273 14139 6307
rect 14565 6273 14599 6307
rect 14657 6273 14691 6307
rect 14841 6273 14875 6307
rect 14933 6273 14967 6307
rect 15485 6273 15519 6307
rect 15945 6273 15979 6307
rect 16129 6273 16163 6307
rect 16865 6273 16899 6307
rect 1409 6205 1443 6239
rect 3157 6205 3191 6239
rect 3525 6205 3559 6239
rect 4721 6205 4755 6239
rect 9321 6205 9355 6239
rect 9689 6205 9723 6239
rect 9965 6205 9999 6239
rect 10793 6205 10827 6239
rect 16313 6205 16347 6239
rect 5181 6137 5215 6171
rect 12633 6137 12667 6171
rect 14289 6137 14323 6171
rect 2513 6069 2547 6103
rect 3893 6069 3927 6103
rect 5733 6069 5767 6103
rect 7389 6069 7423 6103
rect 10333 6069 10367 6103
rect 10517 6069 10551 6103
rect 11529 6069 11563 6103
rect 13461 6069 13495 6103
rect 15117 6069 15151 6103
rect 2881 5865 2915 5899
rect 3893 5865 3927 5899
rect 6653 5865 6687 5899
rect 10333 5865 10367 5899
rect 11989 5865 12023 5899
rect 12909 5865 12943 5899
rect 11161 5797 11195 5831
rect 4445 5729 4479 5763
rect 5273 5729 5307 5763
rect 6929 5729 6963 5763
rect 10793 5729 10827 5763
rect 11713 5729 11747 5763
rect 12265 5729 12299 5763
rect 16957 5729 16991 5763
rect 17785 5729 17819 5763
rect 1501 5661 1535 5695
rect 1768 5661 1802 5695
rect 4261 5661 4295 5695
rect 5540 5661 5574 5695
rect 9321 5661 9355 5695
rect 9505 5661 9539 5695
rect 10149 5661 10183 5695
rect 10701 5661 10735 5695
rect 10885 5661 10919 5695
rect 10985 5661 11019 5695
rect 11529 5661 11563 5695
rect 11621 5661 11655 5695
rect 11805 5661 11839 5695
rect 12449 5661 12483 5695
rect 13277 5661 13311 5695
rect 13553 5661 13587 5695
rect 14289 5661 14323 5695
rect 14749 5661 14783 5695
rect 16773 5661 16807 5695
rect 16865 5661 16899 5695
rect 17509 5661 17543 5695
rect 7196 5593 7230 5627
rect 9781 5593 9815 5627
rect 9965 5593 9999 5627
rect 14105 5593 14139 5627
rect 15016 5593 15050 5627
rect 4353 5525 4387 5559
rect 8309 5525 8343 5559
rect 9505 5525 9539 5559
rect 10057 5525 10091 5559
rect 12633 5525 12667 5559
rect 13369 5525 13403 5559
rect 13737 5525 13771 5559
rect 16129 5525 16163 5559
rect 16405 5525 16439 5559
rect 1409 5321 1443 5355
rect 2145 5321 2179 5355
rect 2881 5321 2915 5355
rect 5365 5321 5399 5355
rect 6377 5321 6411 5355
rect 6745 5321 6779 5355
rect 13553 5321 13587 5355
rect 15117 5321 15151 5355
rect 18061 5321 18095 5355
rect 1777 5185 1811 5219
rect 1961 5185 1995 5219
rect 2789 5185 2823 5219
rect 3873 5185 3907 5219
rect 5825 5185 5859 5219
rect 7573 5185 7607 5219
rect 8668 5185 8702 5219
rect 10701 5185 10735 5219
rect 10793 5185 10827 5219
rect 10885 5185 10919 5219
rect 11069 5185 11103 5219
rect 11713 5185 11747 5219
rect 12173 5185 12207 5219
rect 12429 5185 12463 5219
rect 13921 5185 13955 5219
rect 14381 5185 14415 5219
rect 14565 5185 14599 5219
rect 14657 5185 14691 5219
rect 14933 5185 14967 5219
rect 15393 5185 15427 5219
rect 15577 5185 15611 5219
rect 15669 5185 15703 5219
rect 15761 5185 15795 5219
rect 16681 5185 16715 5219
rect 16948 5185 16982 5219
rect 3065 5117 3099 5151
rect 3617 5117 3651 5151
rect 5641 5117 5675 5151
rect 6837 5117 6871 5151
rect 6929 5117 6963 5151
rect 8401 5117 8435 5151
rect 11897 5117 11931 5151
rect 14749 5117 14783 5151
rect 4997 5049 5031 5083
rect 2421 4981 2455 5015
rect 6009 4981 6043 5015
rect 7389 4981 7423 5015
rect 9781 4981 9815 5015
rect 10425 4981 10459 5015
rect 11529 4981 11563 5015
rect 14013 4981 14047 5015
rect 16037 4981 16071 5015
rect 3065 4777 3099 4811
rect 3893 4777 3927 4811
rect 6469 4777 6503 4811
rect 12541 4777 12575 4811
rect 15945 4777 15979 4811
rect 9505 4709 9539 4743
rect 1685 4641 1719 4675
rect 4629 4641 4663 4675
rect 4905 4641 4939 4675
rect 9137 4641 9171 4675
rect 9597 4641 9631 4675
rect 11897 4641 11931 4675
rect 13093 4641 13127 4675
rect 4077 4573 4111 4607
rect 5089 4573 5123 4607
rect 5273 4573 5307 4607
rect 5733 4573 5767 4607
rect 6285 4573 6319 4607
rect 7113 4573 7147 4607
rect 7380 4573 7414 4607
rect 10425 4573 10459 4607
rect 10609 4573 10643 4607
rect 10701 4573 10735 4607
rect 10793 4573 10827 4607
rect 12173 4573 12207 4607
rect 13277 4573 13311 4607
rect 15577 4573 15611 4607
rect 16221 4573 16255 4607
rect 16405 4573 16439 4607
rect 16957 4573 16991 4607
rect 1930 4505 1964 4539
rect 3341 4505 3375 4539
rect 13369 4505 13403 4539
rect 15310 4505 15344 4539
rect 17224 4505 17258 4539
rect 5549 4437 5583 4471
rect 8493 4437 8527 4471
rect 11069 4437 11103 4471
rect 12081 4437 12115 4471
rect 13737 4437 13771 4471
rect 14197 4437 14231 4471
rect 16589 4437 16623 4471
rect 18337 4437 18371 4471
rect 1685 4233 1719 4267
rect 3341 4233 3375 4267
rect 7113 4233 7147 4267
rect 9873 4233 9907 4267
rect 12265 4233 12299 4267
rect 16865 4233 16899 4267
rect 17325 4233 17359 4267
rect 16313 4165 16347 4199
rect 1501 4097 1535 4131
rect 1961 4097 1995 4131
rect 2145 4097 2179 4131
rect 4169 4097 4203 4131
rect 4896 4097 4930 4131
rect 7757 4097 7791 4131
rect 8024 4097 8058 4131
rect 9413 4097 9447 4131
rect 10149 4097 10183 4131
rect 10333 4097 10367 4131
rect 10517 4097 10551 4131
rect 10977 4097 11011 4131
rect 11161 4097 11195 4131
rect 11713 4097 11747 4131
rect 11897 4097 11931 4131
rect 12449 4097 12483 4131
rect 13185 4097 13219 4131
rect 13829 4097 13863 4131
rect 14289 4097 14323 4131
rect 14749 4097 14783 4131
rect 16129 4097 16163 4131
rect 16681 4097 16715 4131
rect 17509 4097 17543 4131
rect 17693 4097 17727 4131
rect 18061 4097 18095 4131
rect 2329 4029 2363 4063
rect 2697 4029 2731 4063
rect 3433 4029 3467 4063
rect 3525 4029 3559 4063
rect 3985 4029 4019 4063
rect 4629 4029 4663 4063
rect 7205 4029 7239 4063
rect 7297 4029 7331 4063
rect 10609 4029 10643 4063
rect 11989 4029 12023 4063
rect 13645 4029 13679 4063
rect 14013 4029 14047 4063
rect 15853 4029 15887 4063
rect 17785 4029 17819 4063
rect 6009 3961 6043 3995
rect 12909 3961 12943 3995
rect 15945 3961 15979 3995
rect 18245 3961 18279 3995
rect 2973 3893 3007 3927
rect 4353 3893 4387 3927
rect 6745 3893 6779 3927
rect 9137 3893 9171 3927
rect 9505 3893 9539 3927
rect 11529 3893 11563 3927
rect 13369 3893 13403 3927
rect 14473 3893 14507 3927
rect 14933 3893 14967 3927
rect 15577 3893 15611 3927
rect 3893 3689 3927 3723
rect 4905 3689 4939 3723
rect 7113 3689 7147 3723
rect 8953 3689 8987 3723
rect 11989 3689 12023 3723
rect 13369 3689 13403 3723
rect 16865 3689 16899 3723
rect 17785 3689 17819 3723
rect 3433 3621 3467 3655
rect 13093 3621 13127 3655
rect 16497 3621 16531 3655
rect 2053 3553 2087 3587
rect 4353 3553 4387 3587
rect 4537 3553 4571 3587
rect 5457 3553 5491 3587
rect 6745 3553 6779 3587
rect 7389 3553 7423 3587
rect 11713 3553 11747 3587
rect 14657 3553 14691 3587
rect 18153 3553 18187 3587
rect 1593 3485 1627 3519
rect 4261 3485 4295 3519
rect 5365 3485 5399 3519
rect 6929 3485 6963 3519
rect 9229 3485 9263 3519
rect 9321 3485 9355 3519
rect 9413 3485 9447 3519
rect 9597 3485 9631 3519
rect 11446 3485 11480 3519
rect 12173 3485 12207 3519
rect 12265 3485 12299 3519
rect 12909 3485 12943 3519
rect 13553 3485 13587 3519
rect 15301 3485 15335 3519
rect 15945 3485 15979 3519
rect 16221 3485 16255 3519
rect 16405 3485 16439 3519
rect 17049 3485 17083 3519
rect 17141 3485 17175 3519
rect 17969 3485 18003 3519
rect 2320 3417 2354 3451
rect 13737 3417 13771 3451
rect 14473 3417 14507 3451
rect 14565 3417 14599 3451
rect 1777 3349 1811 3383
rect 5273 3349 5307 3383
rect 6101 3349 6135 3383
rect 10057 3349 10091 3383
rect 10333 3349 10367 3383
rect 14105 3349 14139 3383
rect 15117 3349 15151 3383
rect 3157 3145 3191 3179
rect 6009 3145 6043 3179
rect 9965 3145 9999 3179
rect 13737 3145 13771 3179
rect 14473 3145 14507 3179
rect 16129 3145 16163 3179
rect 18061 3145 18095 3179
rect 7512 3077 7546 3111
rect 10333 3077 10367 3111
rect 10977 3077 11011 3111
rect 15016 3077 15050 3111
rect 16926 3077 16960 3111
rect 2513 3009 2547 3043
rect 2697 3009 2731 3043
rect 2881 3009 2915 3043
rect 3341 3009 3375 3043
rect 3985 3009 4019 3043
rect 4252 3009 4286 3043
rect 5733 3009 5767 3043
rect 5825 3009 5859 3043
rect 7757 3009 7791 3043
rect 8217 3009 8251 3043
rect 8852 3009 8886 3043
rect 10241 3009 10275 3043
rect 10425 3009 10459 3043
rect 11161 3009 11195 3043
rect 12734 3009 12768 3043
rect 13001 3009 13035 3043
rect 13829 3009 13863 3043
rect 14749 3009 14783 3043
rect 16681 3009 16715 3043
rect 1961 2941 1995 2975
rect 2237 2941 2271 2975
rect 8585 2941 8619 2975
rect 13921 2941 13955 2975
rect 3617 2873 3651 2907
rect 5365 2873 5399 2907
rect 8033 2873 8067 2907
rect 10793 2873 10827 2907
rect 6377 2805 6411 2839
rect 11621 2805 11655 2839
rect 13369 2805 13403 2839
rect 11621 2601 11655 2635
rect 12817 2601 12851 2635
rect 13737 2601 13771 2635
rect 15669 2601 15703 2635
rect 4169 2533 4203 2567
rect 6561 2533 6595 2567
rect 9137 2533 9171 2567
rect 10149 2533 10183 2567
rect 10609 2533 10643 2567
rect 16037 2533 16071 2567
rect 2237 2465 2271 2499
rect 5733 2465 5767 2499
rect 7113 2465 7147 2499
rect 9597 2465 9631 2499
rect 12081 2465 12115 2499
rect 12265 2465 12299 2499
rect 14289 2465 14323 2499
rect 1961 2397 1995 2431
rect 2513 2397 2547 2431
rect 3433 2397 3467 2431
rect 3985 2397 4019 2431
rect 4905 2397 4939 2431
rect 6009 2397 6043 2431
rect 6929 2397 6963 2431
rect 7021 2397 7055 2431
rect 8125 2397 8159 2431
rect 9321 2397 9355 2431
rect 9505 2397 9539 2431
rect 9965 2397 9999 2431
rect 10425 2397 10459 2431
rect 11161 2397 11195 2431
rect 12633 2397 12667 2431
rect 13369 2397 13403 2431
rect 13553 2397 13587 2431
rect 14556 2397 14590 2431
rect 16221 2397 16255 2431
rect 17141 2397 17175 2431
rect 17785 2397 17819 2431
rect 18061 2397 18095 2431
rect 8585 2329 8619 2363
rect 7941 2261 7975 2295
rect 10977 2261 11011 2295
rect 11989 2261 12023 2295
rect 16957 2261 16991 2295
rect 18245 2261 18279 2295
<< metal1 >>
rect 1104 17434 18860 17456
rect 1104 17382 6880 17434
rect 6932 17382 6944 17434
rect 6996 17382 7008 17434
rect 7060 17382 7072 17434
rect 7124 17382 7136 17434
rect 7188 17382 12811 17434
rect 12863 17382 12875 17434
rect 12927 17382 12939 17434
rect 12991 17382 13003 17434
rect 13055 17382 13067 17434
rect 13119 17382 18860 17434
rect 1104 17360 18860 17382
rect 2685 17323 2743 17329
rect 2685 17289 2697 17323
rect 2731 17320 2743 17323
rect 4338 17320 4344 17332
rect 2731 17292 4344 17320
rect 2731 17289 2743 17292
rect 2685 17283 2743 17289
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 7742 17280 7748 17332
rect 7800 17320 7806 17332
rect 7929 17323 7987 17329
rect 7929 17320 7941 17323
rect 7800 17292 7941 17320
rect 7800 17280 7806 17292
rect 7929 17289 7941 17292
rect 7975 17289 7987 17323
rect 7929 17283 7987 17289
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 10321 17323 10379 17329
rect 10321 17320 10333 17323
rect 9732 17292 10333 17320
rect 9732 17280 9738 17292
rect 10321 17289 10333 17292
rect 10367 17289 10379 17323
rect 10321 17283 10379 17289
rect 14182 17280 14188 17332
rect 14240 17320 14246 17332
rect 14369 17323 14427 17329
rect 14369 17320 14381 17323
rect 14240 17292 14381 17320
rect 14240 17280 14246 17292
rect 14369 17289 14381 17292
rect 14415 17289 14427 17323
rect 14369 17283 14427 17289
rect 18046 17280 18052 17332
rect 18104 17320 18110 17332
rect 18233 17323 18291 17329
rect 18233 17320 18245 17323
rect 18104 17292 18245 17320
rect 18104 17280 18110 17292
rect 18233 17289 18245 17292
rect 18279 17289 18291 17323
rect 18233 17283 18291 17289
rect 3789 17255 3847 17261
rect 3789 17252 3801 17255
rect 2240 17224 3801 17252
rect 1302 17144 1308 17196
rect 1360 17184 1366 17196
rect 2240 17193 2268 17224
rect 3789 17221 3801 17224
rect 3835 17221 3847 17255
rect 8389 17255 8447 17261
rect 8389 17252 8401 17255
rect 3789 17215 3847 17221
rect 6288 17224 6960 17252
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 1360 17156 2237 17184
rect 1360 17144 1366 17156
rect 2225 17153 2237 17156
rect 2271 17153 2283 17187
rect 2225 17147 2283 17153
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17184 2559 17187
rect 2866 17184 2872 17196
rect 2547 17156 2872 17184
rect 2547 17153 2559 17156
rect 2501 17147 2559 17153
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17085 2007 17119
rect 1949 17079 2007 17085
rect 1964 17048 1992 17079
rect 6288 17048 6316 17224
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17184 6423 17187
rect 6546 17184 6552 17196
rect 6411 17156 6552 17184
rect 6411 17153 6423 17156
rect 6365 17147 6423 17153
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 6730 17184 6736 17196
rect 6691 17156 6736 17184
rect 6730 17144 6736 17156
rect 6788 17144 6794 17196
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 6638 17076 6644 17128
rect 6696 17116 6702 17128
rect 6840 17116 6868 17147
rect 6696 17088 6868 17116
rect 6932 17116 6960 17224
rect 7392 17224 8401 17252
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7392 17193 7420 17224
rect 8389 17221 8401 17224
rect 8435 17221 8447 17255
rect 8389 17215 8447 17221
rect 12434 17212 12440 17264
rect 12492 17252 12498 17264
rect 12492 17224 12756 17252
rect 12492 17212 12498 17224
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7340 17156 7389 17184
rect 7340 17144 7346 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 8113 17187 8171 17193
rect 8113 17153 8125 17187
rect 8159 17153 8171 17187
rect 8113 17147 8171 17153
rect 6932 17088 8064 17116
rect 6696 17076 6702 17088
rect 1964 17020 6316 17048
rect 6549 17051 6607 17057
rect 6549 17017 6561 17051
rect 6595 17048 6607 17051
rect 7926 17048 7932 17060
rect 6595 17020 7932 17048
rect 6595 17017 6607 17020
rect 6549 17011 6607 17017
rect 7926 17008 7932 17020
rect 7984 17008 7990 17060
rect 2958 16980 2964 16992
rect 2919 16952 2964 16980
rect 2958 16940 2964 16952
rect 3016 16940 3022 16992
rect 7190 16980 7196 16992
rect 7151 16952 7196 16980
rect 7190 16940 7196 16952
rect 7248 16940 7254 16992
rect 8036 16980 8064 17088
rect 8128 17048 8156 17147
rect 9030 17144 9036 17196
rect 9088 17184 9094 17196
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 9088 17156 9137 17184
rect 9088 17144 9094 17156
rect 9125 17153 9137 17156
rect 9171 17153 9183 17187
rect 9125 17147 9183 17153
rect 10410 17144 10416 17196
rect 10468 17184 10474 17196
rect 10505 17187 10563 17193
rect 10505 17184 10517 17187
rect 10468 17156 10517 17184
rect 10468 17144 10474 17156
rect 10505 17153 10517 17156
rect 10551 17153 10563 17187
rect 10505 17147 10563 17153
rect 11606 17144 11612 17196
rect 11664 17184 11670 17196
rect 12728 17193 12756 17224
rect 12253 17187 12311 17193
rect 12253 17184 12265 17187
rect 11664 17156 12265 17184
rect 11664 17144 11670 17156
rect 12253 17153 12265 17156
rect 12299 17153 12311 17187
rect 12253 17147 12311 17153
rect 12713 17187 12771 17193
rect 12713 17153 12725 17187
rect 12759 17153 12771 17187
rect 13170 17184 13176 17196
rect 13131 17156 13176 17184
rect 12713 17147 12771 17153
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17153 14611 17187
rect 15010 17184 15016 17196
rect 14971 17156 15016 17184
rect 14553 17147 14611 17153
rect 9401 17119 9459 17125
rect 9401 17085 9413 17119
rect 9447 17116 9459 17119
rect 9490 17116 9496 17128
rect 9447 17088 9496 17116
rect 9447 17085 9459 17088
rect 9401 17079 9459 17085
rect 9490 17076 9496 17088
rect 9548 17076 9554 17128
rect 10318 17076 10324 17128
rect 10376 17116 10382 17128
rect 10781 17119 10839 17125
rect 10781 17116 10793 17119
rect 10376 17088 10793 17116
rect 10376 17076 10382 17088
rect 10781 17085 10793 17088
rect 10827 17085 10839 17119
rect 10781 17079 10839 17085
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17116 12495 17119
rect 12618 17116 12624 17128
rect 12483 17088 12624 17116
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 11054 17048 11060 17060
rect 8128 17020 11060 17048
rect 11054 17008 11060 17020
rect 11112 17008 11118 17060
rect 14568 17048 14596 17147
rect 15010 17144 15016 17156
rect 15068 17144 15074 17196
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17184 15439 17187
rect 15657 17187 15715 17193
rect 15657 17184 15669 17187
rect 15427 17156 15669 17184
rect 15427 17153 15439 17156
rect 15381 17147 15439 17153
rect 15657 17153 15669 17156
rect 15703 17184 15715 17187
rect 16758 17184 16764 17196
rect 15703 17156 16764 17184
rect 15703 17153 15715 17156
rect 15657 17147 15715 17153
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17184 16911 17187
rect 17034 17184 17040 17196
rect 16899 17156 17040 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 17497 17187 17555 17193
rect 17497 17153 17509 17187
rect 17543 17184 17555 17187
rect 17586 17184 17592 17196
rect 17543 17156 17592 17184
rect 17543 17153 17555 17156
rect 17497 17147 17555 17153
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 18046 17184 18052 17196
rect 18007 17156 18052 17184
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 16298 17116 16304 17128
rect 16259 17088 16304 17116
rect 16298 17076 16304 17088
rect 16356 17076 16362 17128
rect 15378 17048 15384 17060
rect 14568 17020 15384 17048
rect 15378 17008 15384 17020
rect 15436 17008 15442 17060
rect 15841 17051 15899 17057
rect 15841 17017 15853 17051
rect 15887 17048 15899 17051
rect 17218 17048 17224 17060
rect 15887 17020 17224 17048
rect 15887 17017 15899 17020
rect 15841 17011 15899 17017
rect 17218 17008 17224 17020
rect 17276 17008 17282 17060
rect 17678 17048 17684 17060
rect 17639 17020 17684 17048
rect 17678 17008 17684 17020
rect 17736 17008 17742 17060
rect 10594 16980 10600 16992
rect 8036 16952 10600 16980
rect 10594 16940 10600 16952
rect 10652 16940 10658 16992
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 12069 16983 12127 16989
rect 12069 16980 12081 16983
rect 11940 16952 12081 16980
rect 11940 16940 11946 16952
rect 12069 16949 12081 16952
rect 12115 16949 12127 16983
rect 14826 16980 14832 16992
rect 14787 16952 14832 16980
rect 12069 16943 12127 16949
rect 14826 16940 14832 16952
rect 14884 16940 14890 16992
rect 16666 16980 16672 16992
rect 16627 16952 16672 16980
rect 16666 16940 16672 16952
rect 16724 16940 16730 16992
rect 1104 16890 18860 16912
rect 1104 16838 3915 16890
rect 3967 16838 3979 16890
rect 4031 16838 4043 16890
rect 4095 16838 4107 16890
rect 4159 16838 4171 16890
rect 4223 16838 9846 16890
rect 9898 16838 9910 16890
rect 9962 16838 9974 16890
rect 10026 16838 10038 16890
rect 10090 16838 10102 16890
rect 10154 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 15904 16890
rect 15956 16838 15968 16890
rect 16020 16838 16032 16890
rect 16084 16838 18860 16890
rect 1104 16816 18860 16838
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 2961 16779 3019 16785
rect 2961 16776 2973 16779
rect 2924 16748 2973 16776
rect 2924 16736 2930 16748
rect 2961 16745 2973 16748
rect 3007 16745 3019 16779
rect 2961 16739 3019 16745
rect 5997 16779 6055 16785
rect 5997 16745 6009 16779
rect 6043 16776 6055 16779
rect 6730 16776 6736 16788
rect 6043 16748 6736 16776
rect 6043 16745 6055 16748
rect 5997 16739 6055 16745
rect 6730 16736 6736 16748
rect 6788 16776 6794 16788
rect 8573 16779 8631 16785
rect 6788 16748 7696 16776
rect 6788 16736 6794 16748
rect 1857 16711 1915 16717
rect 1857 16677 1869 16711
rect 1903 16708 1915 16711
rect 2498 16708 2504 16720
rect 1903 16680 2504 16708
rect 1903 16677 1915 16680
rect 1857 16671 1915 16677
rect 2498 16668 2504 16680
rect 2556 16668 2562 16720
rect 3142 16708 3148 16720
rect 3103 16680 3148 16708
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 2406 16640 2412 16652
rect 2367 16612 2412 16640
rect 2406 16600 2412 16612
rect 2464 16600 2470 16652
rect 7668 16649 7696 16748
rect 8573 16745 8585 16779
rect 8619 16776 8631 16779
rect 9030 16776 9036 16788
rect 8619 16748 9036 16776
rect 8619 16745 8631 16748
rect 8573 16739 8631 16745
rect 9030 16736 9036 16748
rect 9088 16736 9094 16788
rect 9140 16748 12388 16776
rect 7742 16668 7748 16720
rect 7800 16708 7806 16720
rect 8113 16711 8171 16717
rect 8113 16708 8125 16711
rect 7800 16680 8125 16708
rect 7800 16668 7806 16680
rect 8113 16677 8125 16680
rect 8159 16677 8171 16711
rect 8113 16671 8171 16677
rect 9140 16652 9168 16748
rect 11606 16708 11612 16720
rect 11567 16680 11612 16708
rect 11606 16668 11612 16680
rect 11664 16668 11670 16720
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16609 7711 16643
rect 9122 16640 9128 16652
rect 9083 16612 9128 16640
rect 7653 16603 7711 16609
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 10318 16600 10324 16652
rect 10376 16640 10382 16652
rect 10962 16640 10968 16652
rect 10376 16612 10968 16640
rect 10376 16600 10382 16612
rect 10962 16600 10968 16612
rect 11020 16640 11026 16652
rect 11333 16643 11391 16649
rect 11333 16640 11345 16643
rect 11020 16612 11345 16640
rect 11020 16600 11026 16612
rect 11333 16609 11345 16612
rect 11379 16640 11391 16643
rect 12250 16640 12256 16652
rect 11379 16612 12256 16640
rect 11379 16609 11391 16612
rect 11333 16603 11391 16609
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 12360 16649 12388 16748
rect 14292 16748 16620 16776
rect 14292 16649 14320 16748
rect 16592 16652 16620 16748
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16640 12403 16643
rect 14277 16643 14335 16649
rect 12391 16612 12480 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 12452 16584 12480 16612
rect 14277 16609 14289 16643
rect 14323 16609 14335 16643
rect 16574 16640 16580 16652
rect 16487 16612 16580 16640
rect 14277 16603 14335 16609
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 14 16532 20 16584
rect 72 16572 78 16584
rect 2958 16572 2964 16584
rect 72 16544 2964 16572
rect 72 16532 78 16544
rect 2958 16532 2964 16544
rect 3016 16532 3022 16584
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4902 16575 4960 16581
rect 4902 16572 4914 16575
rect 4396 16544 4914 16572
rect 4396 16532 4402 16544
rect 4902 16541 4914 16544
rect 4948 16541 4960 16575
rect 5166 16572 5172 16584
rect 5127 16544 5172 16572
rect 4902 16535 4960 16541
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16572 5687 16575
rect 6362 16572 6368 16584
rect 5675 16544 6368 16572
rect 5675 16541 5687 16544
rect 5629 16535 5687 16541
rect 6362 16532 6368 16544
rect 6420 16532 6426 16584
rect 7377 16575 7435 16581
rect 7377 16541 7389 16575
rect 7423 16572 7435 16575
rect 7558 16572 7564 16584
rect 7423 16544 7564 16572
rect 7423 16541 7435 16544
rect 7377 16535 7435 16541
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 7659 16544 7757 16572
rect 1673 16507 1731 16513
rect 1673 16473 1685 16507
rect 1719 16473 1731 16507
rect 2222 16504 2228 16516
rect 2183 16476 2228 16504
rect 1673 16467 1731 16473
rect 1688 16436 1716 16467
rect 2222 16464 2228 16476
rect 2280 16464 2286 16516
rect 3326 16464 3332 16516
rect 3384 16504 3390 16516
rect 3421 16507 3479 16513
rect 3421 16504 3433 16507
rect 3384 16476 3433 16504
rect 3384 16464 3390 16476
rect 3421 16473 3433 16476
rect 3467 16473 3479 16507
rect 3421 16467 3479 16473
rect 7132 16507 7190 16513
rect 7132 16473 7144 16507
rect 7178 16504 7190 16507
rect 7466 16504 7472 16516
rect 7178 16476 7472 16504
rect 7178 16473 7190 16476
rect 7132 16467 7190 16473
rect 7466 16464 7472 16476
rect 7524 16464 7530 16516
rect 1946 16436 1952 16448
rect 1688 16408 1952 16436
rect 1946 16396 1952 16408
rect 2004 16436 2010 16448
rect 2774 16436 2780 16448
rect 2004 16408 2780 16436
rect 2004 16396 2010 16408
rect 2774 16396 2780 16408
rect 2832 16396 2838 16448
rect 3786 16436 3792 16448
rect 3747 16408 3792 16436
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 5445 16439 5503 16445
rect 5445 16405 5457 16439
rect 5491 16436 5503 16439
rect 5534 16436 5540 16448
rect 5491 16408 5540 16436
rect 5491 16405 5503 16408
rect 5445 16399 5503 16405
rect 5534 16396 5540 16408
rect 5592 16396 5598 16448
rect 6638 16396 6644 16448
rect 6696 16436 6702 16448
rect 7659 16436 7687 16544
rect 7745 16541 7757 16544
rect 7791 16541 7803 16575
rect 7926 16572 7932 16584
rect 7887 16544 7932 16572
rect 7745 16535 7803 16541
rect 7926 16532 7932 16544
rect 7984 16532 7990 16584
rect 10226 16532 10232 16584
rect 10284 16572 10290 16584
rect 11241 16575 11299 16581
rect 11241 16572 11253 16575
rect 10284 16544 11253 16572
rect 10284 16532 10290 16544
rect 11241 16541 11253 16544
rect 11287 16572 11299 16575
rect 11698 16572 11704 16584
rect 11287 16544 11704 16572
rect 11287 16541 11299 16544
rect 11241 16535 11299 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 11882 16572 11888 16584
rect 11843 16544 11888 16572
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 12434 16532 12440 16584
rect 12492 16532 12498 16584
rect 14544 16575 14602 16581
rect 14544 16541 14556 16575
rect 14590 16572 14602 16575
rect 14826 16572 14832 16584
rect 14590 16544 14832 16572
rect 14590 16541 14602 16544
rect 14544 16535 14602 16541
rect 14826 16532 14832 16544
rect 14884 16532 14890 16584
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 16833 16575 16891 16581
rect 16833 16572 16845 16575
rect 16724 16544 16845 16572
rect 16724 16532 16730 16544
rect 16833 16541 16845 16544
rect 16879 16541 16891 16575
rect 16833 16535 16891 16541
rect 9398 16513 9404 16516
rect 9392 16467 9404 16513
rect 9456 16504 9462 16516
rect 12590 16507 12648 16513
rect 12590 16504 12602 16507
rect 9456 16476 9492 16504
rect 12084 16476 12602 16504
rect 9398 16464 9404 16467
rect 9456 16464 9462 16476
rect 6696 16408 7687 16436
rect 10505 16439 10563 16445
rect 6696 16396 6702 16408
rect 10505 16405 10517 16439
rect 10551 16436 10563 16439
rect 11238 16436 11244 16448
rect 10551 16408 11244 16436
rect 10551 16405 10563 16408
rect 10505 16399 10563 16405
rect 11238 16396 11244 16408
rect 11296 16396 11302 16448
rect 12084 16445 12112 16476
rect 12590 16473 12602 16476
rect 12636 16473 12648 16507
rect 15930 16504 15936 16516
rect 15891 16476 15936 16504
rect 12590 16467 12648 16473
rect 15930 16464 15936 16476
rect 15988 16464 15994 16516
rect 16114 16464 16120 16516
rect 16172 16504 16178 16516
rect 16172 16476 17540 16504
rect 16172 16464 16178 16476
rect 17512 16448 17540 16476
rect 12069 16439 12127 16445
rect 12069 16405 12081 16439
rect 12115 16405 12127 16439
rect 12069 16399 12127 16405
rect 12158 16396 12164 16448
rect 12216 16436 12222 16448
rect 13446 16436 13452 16448
rect 12216 16408 13452 16436
rect 12216 16396 12222 16408
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 13722 16436 13728 16448
rect 13683 16408 13728 16436
rect 13722 16396 13728 16408
rect 13780 16396 13786 16448
rect 15470 16396 15476 16448
rect 15528 16436 15534 16448
rect 15657 16439 15715 16445
rect 15657 16436 15669 16439
rect 15528 16408 15669 16436
rect 15528 16396 15534 16408
rect 15657 16405 15669 16408
rect 15703 16405 15715 16439
rect 15657 16399 15715 16405
rect 16301 16439 16359 16445
rect 16301 16405 16313 16439
rect 16347 16436 16359 16439
rect 16850 16436 16856 16448
rect 16347 16408 16856 16436
rect 16347 16405 16359 16408
rect 16301 16399 16359 16405
rect 16850 16396 16856 16408
rect 16908 16396 16914 16448
rect 17494 16396 17500 16448
rect 17552 16436 17558 16448
rect 17957 16439 18015 16445
rect 17957 16436 17969 16439
rect 17552 16408 17969 16436
rect 17552 16396 17558 16408
rect 17957 16405 17969 16408
rect 18003 16405 18015 16439
rect 17957 16399 18015 16405
rect 1104 16346 18860 16368
rect 1104 16294 6880 16346
rect 6932 16294 6944 16346
rect 6996 16294 7008 16346
rect 7060 16294 7072 16346
rect 7124 16294 7136 16346
rect 7188 16294 12811 16346
rect 12863 16294 12875 16346
rect 12927 16294 12939 16346
rect 12991 16294 13003 16346
rect 13055 16294 13067 16346
rect 13119 16294 18860 16346
rect 1104 16272 18860 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 2222 16232 2228 16244
rect 2183 16204 2228 16232
rect 2222 16192 2228 16204
rect 2280 16192 2286 16244
rect 3510 16232 3516 16244
rect 3471 16204 3516 16232
rect 3510 16192 3516 16204
rect 3568 16192 3574 16244
rect 3694 16192 3700 16244
rect 3752 16232 3758 16244
rect 5626 16232 5632 16244
rect 3752 16204 5632 16232
rect 3752 16192 3758 16204
rect 5626 16192 5632 16204
rect 5684 16192 5690 16244
rect 6362 16232 6368 16244
rect 6323 16204 6368 16232
rect 6362 16192 6368 16204
rect 6420 16192 6426 16244
rect 9398 16232 9404 16244
rect 9359 16204 9404 16232
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 10226 16232 10232 16244
rect 10187 16204 10232 16232
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 10597 16235 10655 16241
rect 10597 16201 10609 16235
rect 10643 16201 10655 16235
rect 10597 16195 10655 16201
rect 3602 16164 3608 16176
rect 3563 16136 3608 16164
rect 3602 16124 3608 16136
rect 3660 16124 3666 16176
rect 3881 16167 3939 16173
rect 3881 16133 3893 16167
rect 3927 16164 3939 16167
rect 6546 16164 6552 16176
rect 3927 16136 6408 16164
rect 6507 16136 6552 16164
rect 3927 16133 3939 16136
rect 3881 16127 3939 16133
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 2774 16056 2780 16108
rect 2832 16096 2838 16108
rect 2961 16099 3019 16105
rect 2832 16068 2877 16096
rect 2832 16056 2838 16068
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16096 3111 16099
rect 3326 16096 3332 16108
rect 3099 16068 3332 16096
rect 3099 16065 3111 16068
rect 3053 16059 3111 16065
rect 1762 15920 1768 15972
rect 1820 15960 1826 15972
rect 2777 15963 2835 15969
rect 2777 15960 2789 15963
rect 1820 15932 2789 15960
rect 1820 15920 1826 15932
rect 2777 15929 2789 15932
rect 2823 15929 2835 15963
rect 2976 15960 3004 16059
rect 3326 16056 3332 16068
rect 3384 16096 3390 16108
rect 4246 16096 4252 16108
rect 3384 16068 4252 16096
rect 3384 16056 3390 16068
rect 4246 16056 4252 16068
rect 4304 16096 4310 16108
rect 4433 16099 4491 16105
rect 4433 16096 4445 16099
rect 4304 16068 4445 16096
rect 4304 16056 4310 16068
rect 4433 16065 4445 16068
rect 4479 16096 4491 16099
rect 5537 16099 5595 16105
rect 5537 16096 5549 16099
rect 4479 16068 5549 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 5537 16065 5549 16068
rect 5583 16065 5595 16099
rect 5537 16059 5595 16065
rect 5626 16056 5632 16108
rect 5684 16096 5690 16108
rect 6380 16096 6408 16136
rect 6546 16124 6552 16136
rect 6604 16124 6610 16176
rect 6730 16124 6736 16176
rect 6788 16164 6794 16176
rect 10612 16164 10640 16195
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 12584 16204 13124 16232
rect 12584 16192 12590 16204
rect 6788 16136 7420 16164
rect 6788 16124 6794 16136
rect 6638 16096 6644 16108
rect 5684 16068 5729 16096
rect 6380 16068 6644 16096
rect 5684 16056 5690 16068
rect 6638 16056 6644 16068
rect 6696 16096 6702 16108
rect 6917 16099 6975 16105
rect 6917 16096 6929 16099
rect 6696 16068 6929 16096
rect 6696 16056 6702 16068
rect 6917 16065 6929 16068
rect 6963 16065 6975 16099
rect 7190 16096 7196 16108
rect 7151 16068 7196 16096
rect 6917 16059 6975 16065
rect 7190 16056 7196 16068
rect 7248 16056 7254 16108
rect 7392 16105 7420 16136
rect 9600 16136 10640 16164
rect 10781 16167 10839 16173
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 7558 16056 7564 16108
rect 7616 16096 7622 16108
rect 8018 16105 8024 16108
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7616 16068 7757 16096
rect 7616 16056 7622 16068
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 8012 16059 8024 16105
rect 8076 16096 8082 16108
rect 9600 16105 9628 16136
rect 10781 16133 10793 16167
rect 10827 16133 10839 16167
rect 10781 16127 10839 16133
rect 9585 16099 9643 16105
rect 8076 16068 8112 16096
rect 8018 16056 8024 16059
rect 8076 16056 8082 16068
rect 9585 16065 9597 16099
rect 9631 16065 9643 16099
rect 10045 16099 10103 16105
rect 10045 16096 10057 16099
rect 9585 16059 9643 16065
rect 9784 16068 10057 16096
rect 3510 15988 3516 16040
rect 3568 16028 3574 16040
rect 3786 16028 3792 16040
rect 3568 16000 3792 16028
rect 3568 15988 3574 16000
rect 3786 15988 3792 16000
rect 3844 16028 3850 16040
rect 4157 16031 4215 16037
rect 4157 16028 4169 16031
rect 3844 16000 4169 16028
rect 3844 15988 3850 16000
rect 4157 15997 4169 16000
rect 4203 15997 4215 16031
rect 4157 15991 4215 15997
rect 5353 16031 5411 16037
rect 5353 15997 5365 16031
rect 5399 15997 5411 16031
rect 5353 15991 5411 15997
rect 3329 15963 3387 15969
rect 3329 15960 3341 15963
rect 2976 15932 3341 15960
rect 2777 15923 2835 15929
rect 3329 15929 3341 15932
rect 3375 15960 3387 15963
rect 3418 15960 3424 15972
rect 3375 15932 3424 15960
rect 3375 15929 3387 15932
rect 3329 15923 3387 15929
rect 3418 15920 3424 15932
rect 3476 15920 3482 15972
rect 5258 15852 5264 15904
rect 5316 15892 5322 15904
rect 5368 15892 5396 15991
rect 5442 15988 5448 16040
rect 5500 16028 5506 16040
rect 5500 16000 5545 16028
rect 5500 15988 5506 16000
rect 5813 15963 5871 15969
rect 5813 15929 5825 15963
rect 5859 15960 5871 15963
rect 9125 15963 9183 15969
rect 5859 15932 6592 15960
rect 5859 15929 5871 15932
rect 5813 15923 5871 15929
rect 6564 15901 6592 15932
rect 9125 15929 9137 15963
rect 9171 15960 9183 15963
rect 9214 15960 9220 15972
rect 9171 15932 9220 15960
rect 9171 15929 9183 15932
rect 9125 15923 9183 15929
rect 9214 15920 9220 15932
rect 9272 15920 9278 15972
rect 9784 15960 9812 16068
rect 10045 16065 10057 16068
rect 10091 16065 10103 16099
rect 10318 16096 10324 16108
rect 10279 16068 10324 16096
rect 10045 16059 10103 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 9861 16031 9919 16037
rect 9861 15997 9873 16031
rect 9907 16028 9919 16031
rect 10796 16028 10824 16127
rect 12710 16124 12716 16176
rect 12768 16164 12774 16176
rect 12989 16167 13047 16173
rect 12989 16164 13001 16167
rect 12768 16136 13001 16164
rect 12768 16124 12774 16136
rect 12989 16133 13001 16136
rect 13035 16133 13047 16167
rect 13096 16164 13124 16204
rect 13446 16192 13452 16244
rect 13504 16232 13510 16244
rect 14829 16235 14887 16241
rect 13504 16204 13860 16232
rect 13504 16192 13510 16204
rect 13832 16173 13860 16204
rect 14829 16201 14841 16235
rect 14875 16232 14887 16235
rect 15010 16232 15016 16244
rect 14875 16204 15016 16232
rect 14875 16201 14887 16204
rect 14829 16195 14887 16201
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 15286 16192 15292 16244
rect 15344 16232 15350 16244
rect 15673 16235 15731 16241
rect 15673 16232 15685 16235
rect 15344 16204 15685 16232
rect 15344 16192 15350 16204
rect 15673 16201 15685 16204
rect 15719 16201 15731 16235
rect 15841 16235 15899 16241
rect 15841 16232 15853 16235
rect 15673 16195 15731 16201
rect 15764 16204 15853 16232
rect 13601 16167 13659 16173
rect 13601 16164 13613 16167
rect 13096 16136 13613 16164
rect 12989 16127 13047 16133
rect 13601 16133 13613 16136
rect 13647 16133 13659 16167
rect 13601 16127 13659 16133
rect 13817 16167 13875 16173
rect 13817 16133 13829 16167
rect 13863 16133 13875 16167
rect 13817 16127 13875 16133
rect 14645 16167 14703 16173
rect 14645 16133 14657 16167
rect 14691 16164 14703 16167
rect 15194 16164 15200 16176
rect 14691 16136 15200 16164
rect 14691 16133 14703 16136
rect 14645 16127 14703 16133
rect 15194 16124 15200 16136
rect 15252 16124 15258 16176
rect 15470 16164 15476 16176
rect 15431 16136 15476 16164
rect 15470 16124 15476 16136
rect 15528 16124 15534 16176
rect 15764 16164 15792 16204
rect 15841 16201 15853 16204
rect 15887 16232 15899 16235
rect 15930 16232 15936 16244
rect 15887 16204 15936 16232
rect 15887 16201 15899 16204
rect 15841 16195 15899 16201
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 17034 16232 17040 16244
rect 16995 16204 17040 16232
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 16666 16164 16672 16176
rect 15764 16136 16436 16164
rect 16627 16136 16672 16164
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 10928 16068 11529 16096
rect 10928 16056 10934 16068
rect 11517 16065 11529 16068
rect 11563 16096 11575 16099
rect 13262 16096 13268 16108
rect 11563 16068 13268 16096
rect 11563 16065 11575 16068
rect 11517 16059 11575 16065
rect 13262 16056 13268 16068
rect 13320 16096 13326 16108
rect 13722 16096 13728 16108
rect 13320 16068 13728 16096
rect 13320 16056 13326 16068
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 14277 16099 14335 16105
rect 14277 16065 14289 16099
rect 14323 16096 14335 16099
rect 15764 16096 15792 16136
rect 14323 16068 15792 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 16206 16056 16212 16108
rect 16264 16096 16270 16108
rect 16301 16099 16359 16105
rect 16301 16096 16313 16099
rect 16264 16068 16313 16096
rect 16264 16056 16270 16068
rect 16301 16065 16313 16068
rect 16347 16065 16359 16099
rect 16408 16096 16436 16136
rect 16666 16124 16672 16136
rect 16724 16124 16730 16176
rect 16885 16167 16943 16173
rect 16885 16133 16897 16167
rect 16931 16164 16943 16167
rect 17405 16167 17463 16173
rect 17405 16164 17417 16167
rect 16931 16136 17417 16164
rect 16931 16133 16943 16136
rect 16885 16127 16943 16133
rect 17405 16133 17417 16136
rect 17451 16133 17463 16167
rect 17405 16127 17463 16133
rect 17313 16099 17371 16105
rect 17313 16096 17325 16099
rect 16408 16068 17325 16096
rect 16301 16059 16359 16065
rect 17313 16065 17325 16068
rect 17359 16065 17371 16099
rect 17494 16096 17500 16108
rect 17455 16068 17500 16096
rect 17313 16059 17371 16065
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 9907 16000 10824 16028
rect 9907 15997 9919 16000
rect 9861 15991 9919 15997
rect 11698 15988 11704 16040
rect 11756 16028 11762 16040
rect 11793 16031 11851 16037
rect 11793 16028 11805 16031
rect 11756 16000 11805 16028
rect 11756 15988 11762 16000
rect 11793 15997 11805 16000
rect 11839 16028 11851 16031
rect 12066 16028 12072 16040
rect 11839 16000 12072 16028
rect 11839 15997 11851 16000
rect 11793 15991 11851 15997
rect 12066 15988 12072 16000
rect 12124 16028 12130 16040
rect 12124 16000 13676 16028
rect 12124 15988 12130 16000
rect 11149 15963 11207 15969
rect 9784 15932 11100 15960
rect 5316 15864 5396 15892
rect 6549 15895 6607 15901
rect 5316 15852 5322 15864
rect 6549 15861 6561 15895
rect 6595 15861 6607 15895
rect 6549 15855 6607 15861
rect 7282 15852 7288 15904
rect 7340 15892 7346 15904
rect 7377 15895 7435 15901
rect 7377 15892 7389 15895
rect 7340 15864 7389 15892
rect 7340 15852 7346 15864
rect 7377 15861 7389 15864
rect 7423 15892 7435 15895
rect 7926 15892 7932 15904
rect 7423 15864 7932 15892
rect 7423 15861 7435 15864
rect 7377 15855 7435 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 11072 15892 11100 15932
rect 11149 15929 11161 15963
rect 11195 15960 11207 15963
rect 12618 15960 12624 15972
rect 11195 15932 12434 15960
rect 12579 15932 12624 15960
rect 11195 15929 11207 15932
rect 11149 15923 11207 15929
rect 12406 15904 12434 15932
rect 12618 15920 12624 15932
rect 12676 15920 12682 15972
rect 13449 15963 13507 15969
rect 13449 15960 13461 15963
rect 12912 15932 13461 15960
rect 11974 15892 11980 15904
rect 11072 15864 11980 15892
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 12342 15852 12348 15904
rect 12400 15892 12434 15904
rect 12912 15892 12940 15932
rect 13449 15929 13461 15932
rect 13495 15929 13507 15963
rect 13449 15923 13507 15929
rect 12400 15864 12940 15892
rect 12400 15852 12406 15864
rect 12986 15852 12992 15904
rect 13044 15892 13050 15904
rect 13173 15895 13231 15901
rect 13044 15864 13089 15892
rect 13044 15852 13050 15864
rect 13173 15861 13185 15895
rect 13219 15892 13231 15895
rect 13538 15892 13544 15904
rect 13219 15864 13544 15892
rect 13219 15861 13231 15864
rect 13173 15855 13231 15861
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 13648 15901 13676 16000
rect 17402 15988 17408 16040
rect 17460 16028 17466 16040
rect 17773 16031 17831 16037
rect 17773 16028 17785 16031
rect 17460 16000 17785 16028
rect 17460 15988 17466 16000
rect 17773 15997 17785 16000
rect 17819 15997 17831 16031
rect 17773 15991 17831 15997
rect 16117 15963 16175 15969
rect 16117 15960 16129 15963
rect 15672 15932 16129 15960
rect 15672 15904 15700 15932
rect 16117 15929 16129 15932
rect 16163 15929 16175 15963
rect 16117 15923 16175 15929
rect 13633 15895 13691 15901
rect 13633 15861 13645 15895
rect 13679 15861 13691 15895
rect 13633 15855 13691 15861
rect 13998 15852 14004 15904
rect 14056 15892 14062 15904
rect 14645 15895 14703 15901
rect 14645 15892 14657 15895
rect 14056 15864 14657 15892
rect 14056 15852 14062 15864
rect 14645 15861 14657 15864
rect 14691 15861 14703 15895
rect 15654 15892 15660 15904
rect 15615 15864 15660 15892
rect 14645 15855 14703 15861
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 16850 15892 16856 15904
rect 16811 15864 16856 15892
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 1104 15802 18860 15824
rect 1104 15750 3915 15802
rect 3967 15750 3979 15802
rect 4031 15750 4043 15802
rect 4095 15750 4107 15802
rect 4159 15750 4171 15802
rect 4223 15750 9846 15802
rect 9898 15750 9910 15802
rect 9962 15750 9974 15802
rect 10026 15750 10038 15802
rect 10090 15750 10102 15802
rect 10154 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 15904 15802
rect 15956 15750 15968 15802
rect 16020 15750 16032 15802
rect 16084 15750 18860 15802
rect 1104 15728 18860 15750
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 3237 15691 3295 15697
rect 3237 15688 3249 15691
rect 2832 15660 3249 15688
rect 2832 15648 2838 15660
rect 3237 15657 3249 15660
rect 3283 15657 3295 15691
rect 3237 15651 3295 15657
rect 3326 15648 3332 15700
rect 3384 15688 3390 15700
rect 3384 15660 3429 15688
rect 3384 15648 3390 15660
rect 3602 15648 3608 15700
rect 3660 15688 3666 15700
rect 5258 15688 5264 15700
rect 3660 15660 5264 15688
rect 3660 15648 3666 15660
rect 5258 15648 5264 15660
rect 5316 15688 5322 15700
rect 6641 15691 6699 15697
rect 6641 15688 6653 15691
rect 5316 15660 6653 15688
rect 5316 15648 5322 15660
rect 6641 15657 6653 15660
rect 6687 15688 6699 15691
rect 7190 15688 7196 15700
rect 6687 15660 7196 15688
rect 6687 15657 6699 15660
rect 6641 15651 6699 15657
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 10870 15688 10876 15700
rect 10831 15660 10876 15688
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 12345 15691 12403 15697
rect 12345 15657 12357 15691
rect 12391 15688 12403 15691
rect 12618 15688 12624 15700
rect 12391 15660 12624 15688
rect 12391 15657 12403 15660
rect 12345 15651 12403 15657
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 15194 15688 15200 15700
rect 15155 15660 15200 15688
rect 15194 15648 15200 15660
rect 15252 15648 15258 15700
rect 16206 15648 16212 15700
rect 16264 15688 16270 15700
rect 18325 15691 18383 15697
rect 18325 15688 18337 15691
rect 16264 15660 18337 15688
rect 16264 15648 16270 15660
rect 18325 15657 18337 15660
rect 18371 15657 18383 15691
rect 18325 15651 18383 15657
rect 2869 15623 2927 15629
rect 2869 15589 2881 15623
rect 2915 15620 2927 15623
rect 7377 15623 7435 15629
rect 2915 15592 3832 15620
rect 2915 15589 2927 15592
rect 2869 15583 2927 15589
rect 3804 15564 3832 15592
rect 7377 15589 7389 15623
rect 7423 15620 7435 15623
rect 7834 15620 7840 15632
rect 7423 15592 7840 15620
rect 7423 15589 7435 15592
rect 7377 15583 7435 15589
rect 7834 15580 7840 15592
rect 7892 15580 7898 15632
rect 8294 15620 8300 15632
rect 7944 15592 8300 15620
rect 3142 15552 3148 15564
rect 3055 15524 3148 15552
rect 3142 15512 3148 15524
rect 3200 15512 3206 15564
rect 3786 15552 3792 15564
rect 3699 15524 3792 15552
rect 3786 15512 3792 15524
rect 3844 15512 3850 15564
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 1489 15487 1547 15493
rect 1489 15453 1501 15487
rect 1535 15484 1547 15487
rect 1535 15456 1900 15484
rect 1535 15453 1547 15456
rect 1489 15447 1547 15453
rect 1872 15428 1900 15456
rect 1762 15425 1768 15428
rect 1756 15416 1768 15425
rect 1723 15388 1768 15416
rect 1756 15379 1768 15388
rect 1762 15376 1768 15379
rect 1820 15376 1826 15428
rect 1854 15376 1860 15428
rect 1912 15376 1918 15428
rect 3160 15416 3188 15512
rect 3418 15484 3424 15496
rect 3331 15456 3424 15484
rect 3418 15444 3424 15456
rect 3476 15484 3482 15496
rect 4080 15484 4108 15515
rect 5166 15512 5172 15564
rect 5224 15552 5230 15564
rect 5261 15555 5319 15561
rect 5261 15552 5273 15555
rect 5224 15524 5273 15552
rect 5224 15512 5230 15524
rect 5261 15521 5273 15524
rect 5307 15521 5319 15555
rect 7944 15552 7972 15592
rect 8294 15580 8300 15592
rect 8352 15580 8358 15632
rect 11238 15620 11244 15632
rect 11199 15592 11244 15620
rect 11238 15580 11244 15592
rect 11296 15580 11302 15632
rect 8478 15552 8484 15564
rect 5261 15515 5319 15521
rect 7116 15524 7972 15552
rect 8036 15524 8484 15552
rect 4338 15484 4344 15496
rect 3476 15456 4344 15484
rect 3476 15444 3482 15456
rect 4338 15444 4344 15456
rect 4396 15484 4402 15496
rect 5350 15484 5356 15496
rect 4396 15456 5356 15484
rect 4396 15444 4402 15456
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 5534 15493 5540 15496
rect 5528 15484 5540 15493
rect 5495 15456 5540 15484
rect 5528 15447 5540 15456
rect 5534 15444 5540 15447
rect 5592 15444 5598 15496
rect 7116 15493 7144 15524
rect 7101 15487 7159 15493
rect 7101 15453 7113 15487
rect 7147 15453 7159 15487
rect 7101 15447 7159 15453
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15484 7435 15487
rect 7650 15484 7656 15496
rect 7423 15456 7656 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 8036 15493 8064 15524
rect 8478 15512 8484 15524
rect 8536 15552 8542 15564
rect 8536 15524 10272 15552
rect 8536 15512 8542 15524
rect 8021 15487 8079 15493
rect 8021 15453 8033 15487
rect 8067 15453 8079 15487
rect 8021 15447 8079 15453
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 8352 15456 9505 15484
rect 8352 15444 8358 15456
rect 9493 15453 9505 15456
rect 9539 15484 9551 15487
rect 9582 15484 9588 15496
rect 9539 15456 9588 15484
rect 9539 15453 9551 15456
rect 9493 15447 9551 15453
rect 9582 15444 9588 15456
rect 9640 15444 9646 15496
rect 9766 15484 9772 15496
rect 9679 15456 9772 15484
rect 9766 15444 9772 15456
rect 9824 15484 9830 15496
rect 10244 15493 10272 15524
rect 11330 15512 11336 15564
rect 11388 15552 11394 15564
rect 11701 15555 11759 15561
rect 11701 15552 11713 15555
rect 11388 15524 11713 15552
rect 11388 15512 11394 15524
rect 11701 15521 11713 15524
rect 11747 15521 11759 15555
rect 12636 15552 12664 15648
rect 12986 15580 12992 15632
rect 13044 15620 13050 15632
rect 14323 15623 14381 15629
rect 14323 15620 14335 15623
rect 13044 15592 14335 15620
rect 13044 15580 13050 15592
rect 14323 15589 14335 15592
rect 14369 15620 14381 15623
rect 16666 15620 16672 15632
rect 14369 15592 16672 15620
rect 14369 15589 14381 15592
rect 14323 15583 14381 15589
rect 16666 15580 16672 15592
rect 16724 15580 16730 15632
rect 15286 15552 15292 15564
rect 12636 15524 15292 15552
rect 11701 15515 11759 15521
rect 15286 15512 15292 15524
rect 15344 15552 15350 15564
rect 15344 15524 15700 15552
rect 15344 15512 15350 15524
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 9824 15456 10057 15484
rect 9824 15444 9830 15456
rect 10045 15453 10057 15456
rect 10091 15453 10103 15487
rect 10045 15447 10103 15453
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10321 15487 10379 15493
rect 10321 15453 10333 15487
rect 10367 15453 10379 15487
rect 10321 15447 10379 15453
rect 4062 15416 4068 15428
rect 3160 15388 4068 15416
rect 4062 15376 4068 15388
rect 4120 15376 4126 15428
rect 7926 15416 7932 15428
rect 7839 15388 7932 15416
rect 7926 15376 7932 15388
rect 7984 15416 7990 15428
rect 8662 15416 8668 15428
rect 7984 15388 8668 15416
rect 7984 15376 7990 15388
rect 8662 15376 8668 15388
rect 8720 15416 8726 15428
rect 10336 15416 10364 15447
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11609 15487 11667 15493
rect 11609 15484 11621 15487
rect 11204 15456 11621 15484
rect 11204 15444 11210 15456
rect 11609 15453 11621 15456
rect 11655 15453 11667 15487
rect 12066 15484 12072 15496
rect 12027 15456 12072 15484
rect 11609 15447 11667 15453
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 12526 15484 12532 15496
rect 12406 15456 12532 15484
rect 8720 15388 10364 15416
rect 11885 15419 11943 15425
rect 8720 15376 8726 15388
rect 11885 15385 11897 15419
rect 11931 15416 11943 15419
rect 12406 15416 12434 15456
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 12805 15487 12863 15493
rect 12805 15453 12817 15487
rect 12851 15484 12863 15487
rect 12851 15456 13492 15484
rect 12851 15453 12863 15456
rect 12805 15447 12863 15453
rect 12989 15419 13047 15425
rect 12989 15416 13001 15419
rect 11931 15388 12434 15416
rect 12544 15388 13001 15416
rect 11931 15385 11943 15388
rect 11885 15379 11943 15385
rect 7193 15351 7251 15357
rect 7193 15317 7205 15351
rect 7239 15348 7251 15351
rect 7466 15348 7472 15360
rect 7239 15320 7472 15348
rect 7239 15317 7251 15320
rect 7193 15311 7251 15317
rect 7466 15308 7472 15320
rect 7524 15348 7530 15360
rect 7837 15351 7895 15357
rect 7837 15348 7849 15351
rect 7524 15320 7849 15348
rect 7524 15308 7530 15320
rect 7837 15317 7849 15320
rect 7883 15317 7895 15351
rect 8202 15348 8208 15360
rect 8163 15320 8208 15348
rect 7837 15311 7895 15317
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 10686 15348 10692 15360
rect 10647 15320 10692 15348
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 10873 15351 10931 15357
rect 10873 15317 10885 15351
rect 10919 15348 10931 15351
rect 11698 15348 11704 15360
rect 10919 15320 11704 15348
rect 10919 15317 10931 15320
rect 10873 15311 10931 15317
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 11974 15348 11980 15360
rect 11935 15320 11980 15348
rect 11974 15308 11980 15320
rect 12032 15348 12038 15360
rect 12544 15348 12572 15388
rect 12989 15385 13001 15388
rect 13035 15385 13047 15419
rect 13170 15416 13176 15428
rect 13131 15388 13176 15416
rect 12989 15379 13047 15385
rect 13170 15376 13176 15388
rect 13228 15376 13234 15428
rect 13464 15416 13492 15456
rect 13538 15444 13544 15496
rect 13596 15484 13602 15496
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 13596 15456 13645 15484
rect 13596 15444 13602 15456
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13998 15444 14004 15496
rect 14056 15484 14062 15496
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 14056 15456 14105 15484
rect 14056 15444 14062 15456
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 15381 15487 15439 15493
rect 15381 15453 15393 15487
rect 15427 15484 15439 15487
rect 15470 15484 15476 15496
rect 15427 15456 15476 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 15672 15493 15700 15524
rect 16574 15512 16580 15564
rect 16632 15552 16638 15564
rect 16945 15555 17003 15561
rect 16945 15552 16957 15555
rect 16632 15524 16957 15552
rect 16632 15512 16638 15524
rect 16945 15521 16957 15524
rect 16991 15521 17003 15555
rect 16945 15515 17003 15521
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15484 15715 15487
rect 16022 15484 16028 15496
rect 15703 15456 16028 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 16022 15444 16028 15456
rect 16080 15484 16086 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 16080 15456 16129 15484
rect 16080 15444 16086 15456
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 16117 15447 16175 15453
rect 15194 15416 15200 15428
rect 13464 15388 15200 15416
rect 15194 15376 15200 15388
rect 15252 15376 15258 15428
rect 16298 15416 16304 15428
rect 16259 15388 16304 15416
rect 16298 15376 16304 15388
rect 16356 15376 16362 15428
rect 17212 15419 17270 15425
rect 17212 15385 17224 15419
rect 17258 15416 17270 15419
rect 17310 15416 17316 15428
rect 17258 15388 17316 15416
rect 17258 15385 17270 15388
rect 17212 15379 17270 15385
rect 17310 15376 17316 15388
rect 17368 15376 17374 15428
rect 12032 15320 12572 15348
rect 12032 15308 12038 15320
rect 12618 15308 12624 15360
rect 12676 15348 12682 15360
rect 12897 15351 12955 15357
rect 12676 15320 12721 15348
rect 12676 15308 12682 15320
rect 12897 15317 12909 15351
rect 12943 15348 12955 15351
rect 13262 15348 13268 15360
rect 12943 15320 13268 15348
rect 12943 15317 12955 15320
rect 12897 15311 12955 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 13446 15348 13452 15360
rect 13407 15320 13452 15348
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 15565 15351 15623 15357
rect 15565 15317 15577 15351
rect 15611 15348 15623 15351
rect 15654 15348 15660 15360
rect 15611 15320 15660 15348
rect 15611 15317 15623 15320
rect 15565 15311 15623 15317
rect 15654 15308 15660 15320
rect 15712 15348 15718 15360
rect 16316 15348 16344 15376
rect 15712 15320 16344 15348
rect 16485 15351 16543 15357
rect 15712 15308 15718 15320
rect 16485 15317 16497 15351
rect 16531 15348 16543 15351
rect 16850 15348 16856 15360
rect 16531 15320 16856 15348
rect 16531 15317 16543 15320
rect 16485 15311 16543 15317
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 1104 15258 18860 15280
rect 1104 15206 6880 15258
rect 6932 15206 6944 15258
rect 6996 15206 7008 15258
rect 7060 15206 7072 15258
rect 7124 15206 7136 15258
rect 7188 15206 12811 15258
rect 12863 15206 12875 15258
rect 12927 15206 12939 15258
rect 12991 15206 13003 15258
rect 13055 15206 13067 15258
rect 13119 15206 18860 15258
rect 1104 15184 18860 15206
rect 3786 15104 3792 15156
rect 3844 15144 3850 15156
rect 4065 15147 4123 15153
rect 4065 15144 4077 15147
rect 3844 15116 4077 15144
rect 3844 15104 3850 15116
rect 4065 15113 4077 15116
rect 4111 15113 4123 15147
rect 4065 15107 4123 15113
rect 4249 15147 4307 15153
rect 4249 15113 4261 15147
rect 4295 15144 4307 15147
rect 7929 15147 7987 15153
rect 4295 15116 5028 15144
rect 4295 15113 4307 15116
rect 4249 15107 4307 15113
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 14968 1458 15020
rect 5000 15017 5028 15116
rect 7929 15113 7941 15147
rect 7975 15144 7987 15147
rect 8018 15144 8024 15156
rect 7975 15116 8024 15144
rect 7975 15113 7987 15116
rect 7929 15107 7987 15113
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 11701 15147 11759 15153
rect 11701 15113 11713 15147
rect 11747 15144 11759 15147
rect 11974 15144 11980 15156
rect 11747 15116 11980 15144
rect 11747 15113 11759 15116
rect 11701 15107 11759 15113
rect 11974 15104 11980 15116
rect 12032 15104 12038 15156
rect 12710 15144 12716 15156
rect 12671 15116 12716 15144
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 13170 15104 13176 15156
rect 13228 15144 13234 15156
rect 14553 15147 14611 15153
rect 14553 15144 14565 15147
rect 13228 15116 14565 15144
rect 13228 15104 13234 15116
rect 14553 15113 14565 15116
rect 14599 15113 14611 15147
rect 14553 15107 14611 15113
rect 5626 15076 5632 15088
rect 5368 15048 5632 15076
rect 5368 15017 5396 15048
rect 5626 15036 5632 15048
rect 5684 15036 5690 15088
rect 5721 15079 5779 15085
rect 5721 15045 5733 15079
rect 5767 15076 5779 15079
rect 10781 15079 10839 15085
rect 10781 15076 10793 15079
rect 5767 15048 8892 15076
rect 5767 15045 5779 15048
rect 5721 15039 5779 15045
rect 2124 15011 2182 15017
rect 2124 14977 2136 15011
rect 2170 15008 2182 15011
rect 4525 15011 4583 15017
rect 4525 15008 4537 15011
rect 2170 14980 4537 15008
rect 2170 14977 2182 14980
rect 2124 14971 2182 14977
rect 4525 14977 4537 14980
rect 4571 14977 4583 15011
rect 4525 14971 4583 14977
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 14977 4767 15011
rect 4709 14971 4767 14977
rect 4985 15011 5043 15017
rect 4985 14977 4997 15011
rect 5031 15008 5043 15011
rect 5353 15011 5411 15017
rect 5031 14980 5212 15008
rect 5031 14977 5043 14980
rect 4985 14971 5043 14977
rect 1854 14940 1860 14952
rect 1815 14912 1860 14940
rect 1854 14900 1860 14912
rect 1912 14900 1918 14952
rect 3694 14940 3700 14952
rect 3655 14912 3700 14940
rect 3694 14900 3700 14912
rect 3752 14900 3758 14952
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4724 14940 4752 14971
rect 4120 14912 5028 14940
rect 4120 14900 4126 14912
rect 3237 14875 3295 14881
rect 3237 14841 3249 14875
rect 3283 14872 3295 14875
rect 3712 14872 3740 14900
rect 3283 14844 3740 14872
rect 3283 14841 3295 14844
rect 3237 14835 3295 14841
rect 3878 14832 3884 14884
rect 3936 14832 3942 14884
rect 3896 14804 3924 14832
rect 4065 14807 4123 14813
rect 4065 14804 4077 14807
rect 3896 14776 4077 14804
rect 4065 14773 4077 14776
rect 4111 14773 4123 14807
rect 4890 14804 4896 14816
rect 4851 14776 4896 14804
rect 4065 14767 4123 14773
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 5000 14804 5028 14912
rect 5184 14872 5212 14980
rect 5353 14977 5365 15011
rect 5399 14977 5411 15011
rect 5353 14971 5411 14977
rect 6733 15011 6791 15017
rect 6733 14977 6745 15011
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7282 15008 7288 15020
rect 6963 14980 7288 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 5258 14900 5264 14952
rect 5316 14940 5322 14952
rect 5445 14943 5503 14949
rect 5445 14940 5457 14943
rect 5316 14912 5457 14940
rect 5316 14900 5322 14912
rect 5445 14909 5457 14912
rect 5491 14909 5503 14943
rect 5445 14903 5503 14909
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 6270 14940 6276 14952
rect 5592 14912 6276 14940
rect 5592 14900 5598 14912
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 6748 14872 6776 14971
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 15008 7435 15011
rect 7466 15008 7472 15020
rect 7423 14980 7472 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 7392 14940 7420 14971
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 7834 15008 7840 15020
rect 7795 14980 7840 15008
rect 7834 14968 7840 14980
rect 7892 14968 7898 15020
rect 7929 15011 7987 15017
rect 7929 14977 7941 15011
rect 7975 15008 7987 15011
rect 8202 15008 8208 15020
rect 7975 14980 8208 15008
rect 7975 14977 7987 14980
rect 7929 14971 7987 14977
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 8478 15008 8484 15020
rect 8439 14980 8484 15008
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 8662 15008 8668 15020
rect 8623 14980 8668 15008
rect 8662 14968 8668 14980
rect 8720 14968 8726 15020
rect 8864 15017 8892 15048
rect 9508 15048 10793 15076
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 14977 8815 15011
rect 8757 14971 8815 14977
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 15008 8907 15011
rect 9401 15011 9459 15017
rect 9401 15008 9413 15011
rect 8895 14980 9413 15008
rect 8895 14977 8907 14980
rect 8849 14971 8907 14977
rect 9401 14977 9413 14980
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 7650 14940 7656 14952
rect 7064 14912 7420 14940
rect 7611 14912 7656 14940
rect 7064 14900 7070 14912
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 8496 14872 8524 14968
rect 8772 14940 8800 14971
rect 9306 14940 9312 14952
rect 8772 14912 9312 14940
rect 9306 14900 9312 14912
rect 9364 14940 9370 14952
rect 9508 14940 9536 15048
rect 10781 15045 10793 15048
rect 10827 15045 10839 15079
rect 12342 15076 12348 15088
rect 12303 15048 12348 15076
rect 10781 15039 10839 15045
rect 12342 15036 12348 15048
rect 12400 15036 12406 15088
rect 12526 15036 12532 15088
rect 12584 15076 12590 15088
rect 13188 15076 13216 15104
rect 13446 15085 13452 15088
rect 13440 15076 13452 15085
rect 12584 15048 13216 15076
rect 13407 15048 13452 15076
rect 12584 15036 12590 15048
rect 13440 15039 13452 15048
rect 13446 15036 13452 15039
rect 13504 15036 13510 15088
rect 14568 15076 14596 15107
rect 15194 15104 15200 15156
rect 15252 15144 15258 15156
rect 15657 15147 15715 15153
rect 15657 15144 15669 15147
rect 15252 15116 15669 15144
rect 15252 15104 15258 15116
rect 15657 15113 15669 15116
rect 15703 15113 15715 15147
rect 15657 15107 15715 15113
rect 17037 15147 17095 15153
rect 17037 15113 17049 15147
rect 17083 15113 17095 15147
rect 17310 15144 17316 15156
rect 17271 15116 17316 15144
rect 17037 15107 17095 15113
rect 15013 15079 15071 15085
rect 15013 15076 15025 15079
rect 14568 15048 15025 15076
rect 15013 15045 15025 15048
rect 15059 15045 15071 15079
rect 15013 15039 15071 15045
rect 15381 15079 15439 15085
rect 15381 15045 15393 15079
rect 15427 15076 15439 15079
rect 15933 15079 15991 15085
rect 15933 15076 15945 15079
rect 15427 15048 15945 15076
rect 15427 15045 15439 15048
rect 15381 15039 15439 15045
rect 15933 15045 15945 15048
rect 15979 15076 15991 15079
rect 16114 15076 16120 15088
rect 15979 15048 16120 15076
rect 15979 15045 15991 15048
rect 15933 15039 15991 15045
rect 16114 15036 16120 15048
rect 16172 15036 16178 15088
rect 16666 15076 16672 15088
rect 16627 15048 16672 15076
rect 16666 15036 16672 15048
rect 16724 15036 16730 15088
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 16869 15079 16927 15085
rect 16869 15076 16881 15079
rect 16816 15048 16881 15076
rect 16816 15036 16822 15048
rect 16869 15045 16881 15048
rect 16915 15045 16927 15079
rect 16869 15039 16927 15045
rect 9582 14968 9588 15020
rect 9640 15008 9646 15020
rect 9640 14980 9812 15008
rect 9640 14968 9646 14980
rect 9674 14940 9680 14952
rect 9364 14912 9536 14940
rect 9635 14912 9680 14940
rect 9364 14900 9370 14912
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 9784 14940 9812 14980
rect 10226 14968 10232 15020
rect 10284 15008 10290 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 10284 14980 10517 15008
rect 10284 14968 10290 14980
rect 10505 14977 10517 14980
rect 10551 14977 10563 15011
rect 10505 14971 10563 14977
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 12066 15008 12072 15020
rect 10928 14980 10973 15008
rect 12027 14980 12072 15008
rect 10928 14968 10934 14980
rect 12066 14968 12072 14980
rect 12124 14968 12130 15020
rect 15289 15011 15347 15017
rect 15289 14977 15301 15011
rect 15335 15008 15347 15011
rect 15470 15008 15476 15020
rect 15335 14980 15476 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 15008 15715 15011
rect 16298 15008 16304 15020
rect 15703 14980 16304 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 16298 14968 16304 14980
rect 16356 14968 16362 15020
rect 17052 15008 17080 15107
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 17497 15011 17555 15017
rect 17497 15008 17509 15011
rect 17052 14980 17509 15008
rect 17497 14977 17509 14980
rect 17543 14977 17555 15011
rect 18322 15008 18328 15020
rect 18283 14980 18328 15008
rect 17497 14971 17555 14977
rect 18322 14968 18328 14980
rect 18380 14968 18386 15020
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 9784 14912 10701 14940
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12710 14940 12716 14952
rect 12492 14912 12716 14940
rect 12492 14900 12498 14912
rect 12710 14900 12716 14912
rect 12768 14940 12774 14952
rect 13173 14943 13231 14949
rect 13173 14940 13185 14943
rect 12768 14912 13185 14940
rect 12768 14900 12774 14912
rect 13173 14909 13185 14912
rect 13219 14909 13231 14943
rect 15488 14940 15516 14968
rect 15749 14943 15807 14949
rect 15749 14940 15761 14943
rect 15488 14912 15761 14940
rect 13173 14903 13231 14909
rect 15749 14909 15761 14912
rect 15795 14909 15807 14943
rect 15749 14903 15807 14909
rect 5184 14844 8524 14872
rect 9125 14875 9183 14881
rect 9125 14841 9137 14875
rect 9171 14872 9183 14875
rect 11330 14872 11336 14884
rect 9171 14844 11336 14872
rect 9171 14841 9183 14844
rect 9125 14835 9183 14841
rect 11330 14832 11336 14844
rect 11388 14832 11394 14884
rect 15013 14875 15071 14881
rect 15013 14872 15025 14875
rect 12406 14844 12848 14872
rect 6546 14804 6552 14816
rect 5000 14776 6552 14804
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 6638 14764 6644 14816
rect 6696 14804 6702 14816
rect 6825 14807 6883 14813
rect 6825 14804 6837 14807
rect 6696 14776 6837 14804
rect 6696 14764 6702 14776
rect 6825 14773 6837 14776
rect 6871 14773 6883 14807
rect 6825 14767 6883 14773
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 7064 14776 7297 14804
rect 7064 14764 7070 14776
rect 7285 14773 7297 14776
rect 7331 14773 7343 14807
rect 7285 14767 7343 14773
rect 8202 14764 8208 14816
rect 8260 14804 8266 14816
rect 9398 14804 9404 14816
rect 8260 14776 9404 14804
rect 8260 14764 8266 14776
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 10502 14804 10508 14816
rect 10463 14776 10508 14804
rect 10502 14764 10508 14776
rect 10560 14764 10566 14816
rect 10870 14764 10876 14816
rect 10928 14804 10934 14816
rect 11517 14807 11575 14813
rect 11517 14804 11529 14807
rect 10928 14776 11529 14804
rect 10928 14764 10934 14776
rect 11517 14773 11529 14776
rect 11563 14773 11575 14807
rect 11698 14804 11704 14816
rect 11659 14776 11704 14804
rect 11517 14767 11575 14773
rect 11698 14764 11704 14776
rect 11756 14804 11762 14816
rect 12406 14804 12434 14844
rect 11756 14776 12434 14804
rect 12820 14804 12848 14844
rect 14108 14844 15025 14872
rect 14108 14804 14136 14844
rect 15013 14841 15025 14844
rect 15059 14841 15071 14875
rect 15013 14835 15071 14841
rect 15197 14875 15255 14881
rect 15197 14841 15209 14875
rect 15243 14872 15255 14875
rect 16206 14872 16212 14884
rect 15243 14844 16212 14872
rect 15243 14841 15255 14844
rect 15197 14835 15255 14841
rect 16206 14832 16212 14844
rect 16264 14832 16270 14884
rect 16850 14804 16856 14816
rect 12820 14776 14136 14804
rect 16811 14776 16856 14804
rect 11756 14764 11762 14776
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 1104 14714 18860 14736
rect 1104 14662 3915 14714
rect 3967 14662 3979 14714
rect 4031 14662 4043 14714
rect 4095 14662 4107 14714
rect 4159 14662 4171 14714
rect 4223 14662 9846 14714
rect 9898 14662 9910 14714
rect 9962 14662 9974 14714
rect 10026 14662 10038 14714
rect 10090 14662 10102 14714
rect 10154 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 15904 14714
rect 15956 14662 15968 14714
rect 16020 14662 16032 14714
rect 16084 14662 18860 14714
rect 1104 14640 18860 14662
rect 3973 14603 4031 14609
rect 3973 14569 3985 14603
rect 4019 14600 4031 14603
rect 4890 14600 4896 14612
rect 4019 14572 4896 14600
rect 4019 14569 4031 14572
rect 3973 14563 4031 14569
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 5353 14603 5411 14609
rect 5353 14569 5365 14603
rect 5399 14600 5411 14603
rect 5718 14600 5724 14612
rect 5399 14572 5724 14600
rect 5399 14569 5411 14572
rect 5353 14563 5411 14569
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 6270 14600 6276 14612
rect 6231 14572 6276 14600
rect 6270 14560 6276 14572
rect 6328 14560 6334 14612
rect 6457 14603 6515 14609
rect 6457 14569 6469 14603
rect 6503 14600 6515 14603
rect 9306 14600 9312 14612
rect 6503 14572 9312 14600
rect 6503 14569 6515 14572
rect 6457 14563 6515 14569
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 10045 14603 10103 14609
rect 10045 14600 10057 14603
rect 9732 14572 10057 14600
rect 9732 14560 9738 14572
rect 10045 14569 10057 14572
rect 10091 14600 10103 14603
rect 10778 14600 10784 14612
rect 10091 14572 10784 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 10962 14600 10968 14612
rect 10923 14572 10968 14600
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 11793 14603 11851 14609
rect 11793 14569 11805 14603
rect 11839 14600 11851 14603
rect 11974 14600 11980 14612
rect 11839 14572 11980 14600
rect 11839 14569 11851 14572
rect 11793 14563 11851 14569
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 16209 14603 16267 14609
rect 16209 14569 16221 14603
rect 16255 14600 16267 14603
rect 16758 14600 16764 14612
rect 16255 14572 16764 14600
rect 16255 14569 16267 14572
rect 16209 14563 16267 14569
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 17862 14600 17868 14612
rect 17823 14572 17868 14600
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 6914 14532 6920 14544
rect 5644 14504 6920 14532
rect 3694 14424 3700 14476
rect 3752 14464 3758 14476
rect 3789 14467 3847 14473
rect 3789 14464 3801 14467
rect 3752 14436 3801 14464
rect 3752 14424 3758 14436
rect 3789 14433 3801 14436
rect 3835 14433 3847 14467
rect 3789 14427 3847 14433
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 4246 14396 4252 14408
rect 4207 14368 4252 14396
rect 4246 14356 4252 14368
rect 4304 14356 4310 14408
rect 5644 14405 5672 14504
rect 6914 14492 6920 14504
rect 6972 14492 6978 14544
rect 7009 14535 7067 14541
rect 7009 14501 7021 14535
rect 7055 14532 7067 14535
rect 7374 14532 7380 14544
rect 7055 14504 7380 14532
rect 7055 14501 7067 14504
rect 7009 14495 7067 14501
rect 7374 14492 7380 14504
rect 7432 14492 7438 14544
rect 8294 14532 8300 14544
rect 7576 14504 8300 14532
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 7576 14473 7604 14504
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 8938 14532 8944 14544
rect 8899 14504 8944 14532
rect 8938 14492 8944 14504
rect 8996 14492 9002 14544
rect 10134 14492 10140 14544
rect 10192 14532 10198 14544
rect 12618 14532 12624 14544
rect 10192 14504 12624 14532
rect 10192 14492 10198 14504
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 13998 14532 14004 14544
rect 12912 14504 14004 14532
rect 7470 14467 7528 14473
rect 7470 14464 7482 14467
rect 7340 14436 7482 14464
rect 7340 14424 7346 14436
rect 7470 14433 7482 14436
rect 7516 14433 7528 14467
rect 7470 14427 7528 14433
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14433 7619 14467
rect 7561 14427 7619 14433
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 10870 14464 10876 14476
rect 9171 14436 10876 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 12912 14464 12940 14504
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 14093 14535 14151 14541
rect 14093 14501 14105 14535
rect 14139 14501 14151 14535
rect 14093 14495 14151 14501
rect 14108 14464 14136 14495
rect 11072 14436 12940 14464
rect 13004 14436 14136 14464
rect 14737 14467 14795 14473
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 4157 14331 4215 14337
rect 4157 14297 4169 14331
rect 4203 14328 4215 14331
rect 4338 14328 4344 14340
rect 4203 14300 4344 14328
rect 4203 14297 4215 14300
rect 4157 14291 4215 14297
rect 4338 14288 4344 14300
rect 4396 14288 4402 14340
rect 4982 14328 4988 14340
rect 4943 14300 4988 14328
rect 4982 14288 4988 14300
rect 5040 14288 5046 14340
rect 5399 14331 5457 14337
rect 5399 14297 5411 14331
rect 5445 14328 5457 14331
rect 5534 14328 5540 14340
rect 5445 14300 5540 14328
rect 5445 14297 5457 14300
rect 5399 14291 5457 14297
rect 5534 14288 5540 14300
rect 5592 14288 5598 14340
rect 5644 14328 5672 14359
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 5905 14399 5963 14405
rect 5905 14396 5917 14399
rect 5776 14368 5917 14396
rect 5776 14356 5782 14368
rect 5905 14365 5917 14368
rect 5951 14365 5963 14399
rect 6730 14396 6736 14408
rect 6691 14368 6736 14396
rect 5905 14359 5963 14365
rect 6730 14356 6736 14368
rect 6788 14356 6794 14408
rect 7006 14396 7012 14408
rect 6967 14368 7012 14396
rect 7006 14356 7012 14368
rect 7064 14356 7070 14408
rect 7653 14399 7711 14405
rect 7653 14396 7665 14399
rect 7576 14368 7665 14396
rect 5810 14328 5816 14340
rect 5644 14300 5816 14328
rect 5810 14288 5816 14300
rect 5868 14288 5874 14340
rect 5994 14288 6000 14340
rect 6052 14328 6058 14340
rect 6917 14331 6975 14337
rect 6917 14328 6929 14331
rect 6052 14300 6929 14328
rect 6052 14288 6058 14300
rect 6917 14297 6929 14300
rect 6963 14328 6975 14331
rect 7098 14328 7104 14340
rect 6963 14300 7104 14328
rect 6963 14297 6975 14300
rect 6917 14291 6975 14297
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 5000 14260 5028 14288
rect 5258 14260 5264 14272
rect 5000 14232 5264 14260
rect 5258 14220 5264 14232
rect 5316 14260 5322 14272
rect 6273 14263 6331 14269
rect 6273 14260 6285 14263
rect 5316 14232 6285 14260
rect 5316 14220 5322 14232
rect 6273 14229 6285 14232
rect 6319 14229 6331 14263
rect 6273 14223 6331 14229
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 7340 14232 7385 14260
rect 7340 14220 7346 14232
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 7576 14260 7604 14368
rect 7653 14365 7665 14368
rect 7699 14365 7711 14399
rect 7653 14359 7711 14365
rect 7742 14356 7748 14408
rect 7800 14396 7806 14408
rect 9217 14399 9275 14405
rect 7800 14368 7845 14396
rect 7800 14356 7806 14368
rect 9217 14365 9229 14399
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 8294 14328 8300 14340
rect 8255 14300 8300 14328
rect 8294 14288 8300 14300
rect 8352 14288 8358 14340
rect 8478 14288 8484 14340
rect 8536 14328 8542 14340
rect 9030 14328 9036 14340
rect 8536 14300 9036 14328
rect 8536 14288 8542 14300
rect 9030 14288 9036 14300
rect 9088 14288 9094 14340
rect 7926 14260 7932 14272
rect 7524 14232 7932 14260
rect 7524 14220 7530 14232
rect 7926 14220 7932 14232
rect 7984 14220 7990 14272
rect 8110 14260 8116 14272
rect 8071 14232 8116 14260
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 8312 14260 8340 14288
rect 9232 14260 9260 14359
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 11072 14396 11100 14436
rect 9640 14368 11100 14396
rect 9640 14356 9646 14368
rect 11238 14356 11244 14408
rect 11296 14396 11302 14408
rect 11609 14399 11667 14405
rect 11609 14396 11621 14399
rect 11296 14368 11621 14396
rect 11296 14356 11302 14368
rect 11609 14365 11621 14368
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 12526 14356 12532 14408
rect 12584 14396 12590 14408
rect 13004 14405 13032 14436
rect 14737 14433 14749 14467
rect 14783 14464 14795 14467
rect 16577 14467 16635 14473
rect 16577 14464 16589 14467
rect 14783 14436 15240 14464
rect 14783 14433 14795 14436
rect 14737 14427 14795 14433
rect 12713 14399 12771 14405
rect 12713 14396 12725 14399
rect 12584 14368 12725 14396
rect 12584 14356 12590 14368
rect 12713 14365 12725 14368
rect 12759 14365 12771 14399
rect 12713 14359 12771 14365
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14365 12955 14399
rect 12897 14359 12955 14365
rect 12989 14399 13047 14405
rect 12989 14365 13001 14399
rect 13035 14365 13047 14399
rect 12989 14359 13047 14365
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13262 14396 13268 14408
rect 13127 14368 13268 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 9766 14288 9772 14340
rect 9824 14328 9830 14340
rect 9861 14331 9919 14337
rect 9861 14328 9873 14331
rect 9824 14300 9873 14328
rect 9824 14288 9830 14300
rect 9861 14297 9873 14300
rect 9907 14297 9919 14331
rect 9861 14291 9919 14297
rect 10077 14331 10135 14337
rect 10077 14297 10089 14331
rect 10123 14328 10135 14331
rect 10686 14328 10692 14340
rect 10123 14300 10692 14328
rect 10123 14297 10135 14300
rect 10077 14291 10135 14297
rect 10686 14288 10692 14300
rect 10744 14288 10750 14340
rect 11146 14328 11152 14340
rect 11107 14300 11152 14328
rect 11146 14288 11152 14300
rect 11204 14288 11210 14340
rect 11330 14328 11336 14340
rect 11291 14300 11336 14328
rect 11330 14288 11336 14300
rect 11388 14288 11394 14340
rect 12434 14288 12440 14340
rect 12492 14328 12498 14340
rect 12912 14328 12940 14359
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 14090 14356 14096 14408
rect 14148 14396 14154 14408
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 14148 14368 14565 14396
rect 14148 14356 14154 14368
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 15120 14328 15148 14359
rect 12492 14300 12940 14328
rect 13188 14300 15148 14328
rect 12492 14288 12498 14300
rect 8312 14232 9260 14260
rect 9306 14220 9312 14272
rect 9364 14260 9370 14272
rect 9585 14263 9643 14269
rect 9585 14260 9597 14263
rect 9364 14232 9597 14260
rect 9364 14220 9370 14232
rect 9585 14229 9597 14232
rect 9631 14229 9643 14263
rect 9585 14223 9643 14229
rect 9674 14220 9680 14272
rect 9732 14260 9738 14272
rect 10226 14260 10232 14272
rect 9732 14232 10232 14260
rect 9732 14220 9738 14232
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 11164 14260 11192 14288
rect 13188 14260 13216 14300
rect 13354 14260 13360 14272
rect 11164 14232 13216 14260
rect 13315 14232 13360 14260
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 14458 14260 14464 14272
rect 14419 14232 14464 14260
rect 14458 14220 14464 14232
rect 14516 14220 14522 14272
rect 15212 14260 15240 14436
rect 15764 14436 16589 14464
rect 15289 14399 15347 14405
rect 15289 14365 15301 14399
rect 15335 14365 15347 14399
rect 15289 14359 15347 14365
rect 15304 14328 15332 14359
rect 15562 14356 15568 14408
rect 15620 14396 15626 14408
rect 15764 14405 15792 14436
rect 16577 14433 16589 14436
rect 16623 14433 16635 14467
rect 16577 14427 16635 14433
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15620 14368 15761 14396
rect 15620 14356 15626 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 16114 14396 16120 14408
rect 16075 14368 16120 14396
rect 15749 14359 15807 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 16298 14396 16304 14408
rect 16259 14368 16304 14396
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 18322 14396 18328 14408
rect 18283 14368 18328 14396
rect 18322 14356 18328 14368
rect 18380 14356 18386 14408
rect 18230 14328 18236 14340
rect 15304 14300 18236 14328
rect 18230 14288 18236 14300
rect 18288 14288 18294 14340
rect 15289 14263 15347 14269
rect 15289 14260 15301 14263
rect 15212 14232 15301 14260
rect 15289 14229 15301 14232
rect 15335 14260 15347 14263
rect 15378 14260 15384 14272
rect 15335 14232 15384 14260
rect 15335 14229 15347 14232
rect 15289 14223 15347 14229
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 15562 14260 15568 14272
rect 15523 14232 15568 14260
rect 15562 14220 15568 14232
rect 15620 14220 15626 14272
rect 1104 14170 18860 14192
rect 1104 14118 6880 14170
rect 6932 14118 6944 14170
rect 6996 14118 7008 14170
rect 7060 14118 7072 14170
rect 7124 14118 7136 14170
rect 7188 14118 12811 14170
rect 12863 14118 12875 14170
rect 12927 14118 12939 14170
rect 12991 14118 13003 14170
rect 13055 14118 13067 14170
rect 13119 14118 18860 14170
rect 1104 14096 18860 14118
rect 5813 14059 5871 14065
rect 5813 14025 5825 14059
rect 5859 14056 5871 14059
rect 5994 14056 6000 14068
rect 5859 14028 6000 14056
rect 5859 14025 5871 14028
rect 5813 14019 5871 14025
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 7374 14016 7380 14068
rect 7432 14056 7438 14068
rect 9519 14059 9577 14065
rect 9519 14056 9531 14059
rect 7432 14028 7788 14056
rect 7432 14016 7438 14028
rect 5166 13988 5172 14000
rect 3344 13960 5172 13988
rect 3344 13929 3372 13960
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 6086 13948 6092 14000
rect 6144 13988 6150 14000
rect 6609 13991 6667 13997
rect 6609 13988 6621 13991
rect 6144 13960 6621 13988
rect 6144 13948 6150 13960
rect 6609 13957 6621 13960
rect 6655 13957 6667 13991
rect 6609 13951 6667 13957
rect 6825 13991 6883 13997
rect 6825 13957 6837 13991
rect 6871 13988 6883 13991
rect 7760 13988 7788 14028
rect 8772 14028 9531 14056
rect 6871 13960 7420 13988
rect 7760 13960 8708 13988
rect 6871 13957 6883 13960
rect 6825 13951 6883 13957
rect 3602 13929 3608 13932
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 3596 13883 3608 13929
rect 3660 13920 3666 13932
rect 3660 13892 3696 13920
rect 3602 13880 3608 13883
rect 3660 13880 3666 13892
rect 4522 13880 4528 13932
rect 4580 13920 4586 13932
rect 4982 13920 4988 13932
rect 4580 13892 4988 13920
rect 4580 13880 4586 13892
rect 4982 13880 4988 13892
rect 5040 13920 5046 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 5040 13892 5273 13920
rect 5040 13880 5046 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 5629 13923 5687 13929
rect 5629 13889 5641 13923
rect 5675 13920 5687 13923
rect 5718 13920 5724 13932
rect 5675 13892 5724 13920
rect 5675 13889 5687 13892
rect 5629 13883 5687 13889
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 4338 13812 4344 13864
rect 4396 13852 4402 13864
rect 7101 13855 7159 13861
rect 7101 13852 7113 13855
rect 4396 13824 7113 13852
rect 4396 13812 4402 13824
rect 7101 13821 7113 13824
rect 7147 13821 7159 13855
rect 7392 13852 7420 13960
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 7561 13923 7619 13929
rect 7561 13920 7573 13923
rect 7524 13892 7573 13920
rect 7524 13880 7530 13892
rect 7561 13889 7573 13892
rect 7607 13889 7619 13923
rect 7742 13920 7748 13932
rect 7703 13892 7748 13920
rect 7561 13883 7619 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 7926 13920 7932 13932
rect 7883 13892 7932 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 8680 13929 8708 13960
rect 8772 13929 8800 14028
rect 9519 14025 9531 14028
rect 9565 14056 9577 14059
rect 9953 14059 10011 14065
rect 9953 14056 9965 14059
rect 9565 14028 9965 14056
rect 9565 14025 9577 14028
rect 9519 14019 9577 14025
rect 9953 14025 9965 14028
rect 9999 14025 10011 14059
rect 11146 14056 11152 14068
rect 9953 14019 10011 14025
rect 10704 14028 11152 14056
rect 8846 13948 8852 14000
rect 8904 13988 8910 14000
rect 9309 13991 9367 13997
rect 9309 13988 9321 13991
rect 8904 13960 9321 13988
rect 8904 13948 8910 13960
rect 9309 13957 9321 13960
rect 9355 13957 9367 13991
rect 9309 13951 9367 13957
rect 9398 13948 9404 14000
rect 9456 13988 9462 14000
rect 10704 13988 10732 14028
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 13262 14056 13268 14068
rect 12084 14028 13268 14056
rect 9456 13960 10732 13988
rect 9456 13948 9462 13960
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13889 8723 13923
rect 8665 13883 8723 13889
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13920 9091 13923
rect 9674 13920 9680 13932
rect 9079 13892 9680 13920
rect 9079 13889 9091 13892
rect 9033 13883 9091 13889
rect 8846 13852 8852 13864
rect 7392 13824 8852 13852
rect 7101 13815 7159 13821
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 5258 13744 5264 13796
rect 5316 13784 5322 13796
rect 8956 13784 8984 13883
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 9968 13929 9996 13960
rect 10778 13948 10784 14000
rect 10836 13988 10842 14000
rect 10873 13991 10931 13997
rect 10873 13988 10885 13991
rect 10836 13960 10885 13988
rect 10836 13948 10842 13960
rect 10873 13957 10885 13960
rect 10919 13988 10931 13991
rect 12084 13988 12112 14028
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 14516 14028 14749 14056
rect 14516 14016 14522 14028
rect 14737 14025 14749 14028
rect 14783 14056 14795 14059
rect 15194 14056 15200 14068
rect 14783 14028 15200 14056
rect 14783 14025 14795 14028
rect 14737 14019 14795 14025
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 16666 14016 16672 14068
rect 16724 14056 16730 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 16724 14028 18061 14056
rect 16724 14016 16730 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 10919 13960 12112 13988
rect 10919 13957 10931 13960
rect 10873 13951 10931 13957
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13889 10011 13923
rect 10134 13920 10140 13932
rect 10095 13892 10140 13920
rect 9953 13883 10011 13889
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 12084 13929 12112 13960
rect 12342 13948 12348 14000
rect 12400 13988 12406 14000
rect 12980 13991 13038 13997
rect 12400 13960 12940 13988
rect 12400 13948 12406 13960
rect 12069 13923 12127 13929
rect 12069 13889 12081 13923
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12176 13852 12204 13883
rect 12250 13880 12256 13932
rect 12308 13920 12314 13932
rect 12452 13929 12480 13960
rect 12437 13923 12495 13929
rect 12308 13892 12353 13920
rect 12308 13880 12314 13892
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 12710 13920 12716 13932
rect 12483 13892 12517 13920
rect 12671 13892 12716 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 12912 13920 12940 13960
rect 12980 13957 12992 13991
rect 13026 13988 13038 13991
rect 13354 13988 13360 14000
rect 13026 13960 13360 13988
rect 13026 13957 13038 13960
rect 12980 13951 13038 13957
rect 13354 13948 13360 13960
rect 13412 13948 13418 14000
rect 14642 13920 14648 13932
rect 12912 13892 14648 13920
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 15850 13923 15908 13929
rect 15850 13920 15862 13923
rect 15344 13892 15862 13920
rect 15344 13880 15350 13892
rect 15850 13889 15862 13892
rect 15896 13889 15908 13923
rect 15850 13883 15908 13889
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 16574 13920 16580 13932
rect 16163 13892 16580 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16574 13880 16580 13892
rect 16632 13920 16638 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16632 13892 16681 13920
rect 16632 13880 16638 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 16758 13880 16764 13932
rect 16816 13920 16822 13932
rect 16925 13923 16983 13929
rect 16925 13920 16937 13923
rect 16816 13892 16937 13920
rect 16816 13880 16822 13892
rect 16925 13889 16937 13892
rect 16971 13889 16983 13923
rect 16925 13883 16983 13889
rect 12618 13852 12624 13864
rect 12176 13824 12624 13852
rect 12618 13812 12624 13824
rect 12676 13812 12682 13864
rect 10502 13784 10508 13796
rect 5316 13756 8984 13784
rect 9508 13756 10508 13784
rect 5316 13744 5322 13756
rect 4706 13716 4712 13728
rect 4619 13688 4712 13716
rect 4706 13676 4712 13688
rect 4764 13716 4770 13728
rect 5534 13716 5540 13728
rect 4764 13688 5540 13716
rect 4764 13676 4770 13688
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 6457 13719 6515 13725
rect 6457 13685 6469 13719
rect 6503 13716 6515 13719
rect 6546 13716 6552 13728
rect 6503 13688 6552 13716
rect 6503 13685 6515 13688
rect 6457 13679 6515 13685
rect 6546 13676 6552 13688
rect 6604 13676 6610 13728
rect 6638 13676 6644 13728
rect 6696 13716 6702 13728
rect 7926 13716 7932 13728
rect 6696 13688 7932 13716
rect 6696 13676 6702 13688
rect 7926 13676 7932 13688
rect 7984 13676 7990 13728
rect 8202 13676 8208 13728
rect 8260 13716 8266 13728
rect 9508 13725 9536 13756
rect 10502 13744 10508 13756
rect 10560 13744 10566 13796
rect 10686 13784 10692 13796
rect 10647 13756 10692 13784
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 8481 13719 8539 13725
rect 8481 13716 8493 13719
rect 8260 13688 8493 13716
rect 8260 13676 8266 13688
rect 8481 13685 8493 13688
rect 8527 13685 8539 13719
rect 8481 13679 8539 13685
rect 9493 13719 9551 13725
rect 9493 13685 9505 13719
rect 9539 13685 9551 13719
rect 9493 13679 9551 13685
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 9677 13719 9735 13725
rect 9677 13716 9689 13719
rect 9640 13688 9689 13716
rect 9640 13676 9646 13688
rect 9677 13685 9689 13688
rect 9723 13685 9735 13719
rect 11790 13716 11796 13728
rect 11751 13688 11796 13716
rect 9677 13679 9735 13685
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 14090 13716 14096 13728
rect 14051 13688 14096 13716
rect 14090 13676 14096 13688
rect 14148 13676 14154 13728
rect 1104 13626 18860 13648
rect 1104 13574 3915 13626
rect 3967 13574 3979 13626
rect 4031 13574 4043 13626
rect 4095 13574 4107 13626
rect 4159 13574 4171 13626
rect 4223 13574 9846 13626
rect 9898 13574 9910 13626
rect 9962 13574 9974 13626
rect 10026 13574 10038 13626
rect 10090 13574 10102 13626
rect 10154 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 15904 13626
rect 15956 13574 15968 13626
rect 16020 13574 16032 13626
rect 16084 13574 18860 13626
rect 1104 13552 18860 13574
rect 3602 13472 3608 13524
rect 3660 13512 3666 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3660 13484 3801 13512
rect 3660 13472 3666 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 5258 13512 5264 13524
rect 3789 13475 3847 13481
rect 4172 13484 5028 13512
rect 5219 13484 5264 13512
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 1912 13280 2053 13308
rect 1912 13268 1918 13280
rect 2041 13277 2053 13280
rect 2087 13308 2099 13311
rect 3786 13308 3792 13320
rect 2087 13280 3792 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4172 13308 4200 13484
rect 4893 13447 4951 13453
rect 4893 13413 4905 13447
rect 4939 13413 4951 13447
rect 5000 13444 5028 13484
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5350 13472 5356 13524
rect 5408 13512 5414 13524
rect 5721 13515 5779 13521
rect 5721 13512 5733 13515
rect 5408 13484 5733 13512
rect 5408 13472 5414 13484
rect 5721 13481 5733 13484
rect 5767 13481 5779 13515
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 5721 13475 5779 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 7009 13515 7067 13521
rect 7009 13481 7021 13515
rect 7055 13512 7067 13515
rect 7374 13512 7380 13524
rect 7055 13484 7380 13512
rect 7055 13481 7067 13484
rect 7009 13475 7067 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 8202 13512 8208 13524
rect 8163 13484 8208 13512
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 9125 13515 9183 13521
rect 9125 13481 9137 13515
rect 9171 13512 9183 13515
rect 11882 13512 11888 13524
rect 9171 13484 11888 13512
rect 9171 13481 9183 13484
rect 9125 13475 9183 13481
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 18230 13472 18236 13524
rect 18288 13512 18294 13524
rect 18325 13515 18383 13521
rect 18325 13512 18337 13515
rect 18288 13484 18337 13512
rect 18288 13472 18294 13484
rect 18325 13481 18337 13484
rect 18371 13481 18383 13515
rect 18325 13475 18383 13481
rect 8389 13447 8447 13453
rect 8389 13444 8401 13447
rect 5000 13416 8401 13444
rect 4893 13407 4951 13413
rect 8389 13413 8401 13416
rect 8435 13413 8447 13447
rect 8389 13407 8447 13413
rect 4908 13376 4936 13407
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 11238 13444 11244 13456
rect 11112 13416 11244 13444
rect 11112 13404 11118 13416
rect 11238 13404 11244 13416
rect 11296 13404 11302 13456
rect 12710 13404 12716 13456
rect 12768 13444 12774 13456
rect 13173 13447 13231 13453
rect 13173 13444 13185 13447
rect 12768 13416 13185 13444
rect 12768 13404 12774 13416
rect 13173 13413 13185 13416
rect 13219 13413 13231 13447
rect 15378 13444 15384 13456
rect 13173 13407 13231 13413
rect 14384 13416 15384 13444
rect 4908 13348 5488 13376
rect 5460 13320 5488 13348
rect 4019 13280 4200 13308
rect 4249 13311 4307 13317
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4249 13277 4261 13311
rect 4295 13308 4307 13311
rect 4522 13308 4528 13320
rect 4295 13280 4528 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 2308 13243 2366 13249
rect 2308 13209 2320 13243
rect 2354 13240 2366 13243
rect 2590 13240 2596 13252
rect 2354 13212 2596 13240
rect 2354 13209 2366 13212
rect 2308 13203 2366 13209
rect 2590 13200 2596 13212
rect 2648 13200 2654 13252
rect 4264 13240 4292 13271
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4706 13308 4712 13320
rect 4667 13280 4712 13308
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 5350 13308 5356 13320
rect 5311 13280 5356 13308
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 5721 13311 5779 13317
rect 5721 13308 5733 13311
rect 5500 13280 5733 13308
rect 5500 13268 5506 13280
rect 5721 13277 5733 13280
rect 5767 13277 5779 13311
rect 5721 13271 5779 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 7834 13308 7840 13320
rect 7795 13280 7840 13308
rect 5813 13271 5871 13277
rect 3436 13212 4292 13240
rect 5169 13243 5227 13249
rect 3436 13181 3464 13212
rect 5169 13209 5181 13243
rect 5215 13240 5227 13243
rect 5258 13240 5264 13252
rect 5215 13212 5264 13240
rect 5215 13209 5227 13212
rect 5169 13203 5227 13209
rect 5258 13200 5264 13212
rect 5316 13240 5322 13252
rect 5828 13240 5856 13271
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 7984 13280 8953 13308
rect 7984 13268 7990 13280
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 9088 13280 9137 13308
rect 9088 13268 9094 13280
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 9861 13311 9919 13317
rect 9861 13277 9873 13311
rect 9907 13308 9919 13311
rect 11422 13308 11428 13320
rect 9907 13280 11428 13308
rect 9907 13277 9919 13280
rect 9861 13271 9919 13277
rect 11422 13268 11428 13280
rect 11480 13308 11486 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 11480 13280 11529 13308
rect 11480 13268 11486 13280
rect 11517 13277 11529 13280
rect 11563 13308 11575 13311
rect 12728 13308 12756 13404
rect 11563 13280 12756 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 14384 13252 14412 13416
rect 15378 13404 15384 13416
rect 15436 13444 15442 13456
rect 15436 13416 15516 13444
rect 15436 13404 15442 13416
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 15488 13385 15516 13416
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 15252 13348 15301 13376
rect 15252 13336 15258 13348
rect 15289 13345 15301 13348
rect 15335 13345 15347 13379
rect 15289 13339 15347 13345
rect 15473 13379 15531 13385
rect 15473 13345 15485 13379
rect 15519 13345 15531 13379
rect 16482 13376 16488 13388
rect 16443 13348 16488 13376
rect 15473 13339 15531 13345
rect 16482 13336 16488 13348
rect 16540 13336 16546 13388
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 16942 13376 16948 13388
rect 16632 13348 16948 13376
rect 16632 13336 16638 13348
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 16393 13311 16451 13317
rect 16393 13308 16405 13311
rect 15212 13280 16405 13308
rect 5316 13212 5856 13240
rect 5316 13200 5322 13212
rect 6730 13200 6736 13252
rect 6788 13240 6794 13252
rect 7193 13243 7251 13249
rect 7193 13240 7205 13243
rect 6788 13212 7205 13240
rect 6788 13200 6794 13212
rect 7193 13209 7205 13212
rect 7239 13240 7251 13243
rect 7239 13212 8064 13240
rect 7239 13209 7251 13212
rect 7193 13203 7251 13209
rect 3421 13175 3479 13181
rect 3421 13141 3433 13175
rect 3467 13141 3479 13175
rect 3421 13135 3479 13141
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 4433 13175 4491 13181
rect 4433 13172 4445 13175
rect 4304 13144 4445 13172
rect 4304 13132 4310 13144
rect 4433 13141 4445 13144
rect 4479 13141 4491 13175
rect 4433 13135 4491 13141
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 6825 13175 6883 13181
rect 6825 13172 6837 13175
rect 5592 13144 6837 13172
rect 5592 13132 5598 13144
rect 6825 13141 6837 13144
rect 6871 13141 6883 13175
rect 6825 13135 6883 13141
rect 6993 13175 7051 13181
rect 6993 13141 7005 13175
rect 7039 13172 7051 13175
rect 7282 13172 7288 13184
rect 7039 13144 7288 13172
rect 7039 13141 7051 13144
rect 6993 13135 7051 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 8036 13172 8064 13212
rect 8110 13200 8116 13252
rect 8168 13240 8174 13252
rect 8205 13243 8263 13249
rect 8205 13240 8217 13243
rect 8168 13212 8217 13240
rect 8168 13200 8174 13212
rect 8205 13209 8217 13212
rect 8251 13209 8263 13243
rect 8205 13203 8263 13209
rect 10128 13243 10186 13249
rect 10128 13209 10140 13243
rect 10174 13240 10186 13243
rect 10410 13240 10416 13252
rect 10174 13212 10416 13240
rect 10174 13209 10186 13212
rect 10128 13203 10186 13209
rect 10410 13200 10416 13212
rect 10468 13200 10474 13252
rect 11790 13249 11796 13252
rect 11784 13240 11796 13249
rect 11751 13212 11796 13240
rect 11784 13203 11796 13212
rect 11790 13200 11796 13203
rect 11848 13200 11854 13252
rect 13357 13243 13415 13249
rect 13357 13209 13369 13243
rect 13403 13240 13415 13243
rect 13446 13240 13452 13252
rect 13403 13212 13452 13240
rect 13403 13209 13415 13212
rect 13357 13203 13415 13209
rect 13446 13200 13452 13212
rect 13504 13200 13510 13252
rect 14366 13240 14372 13252
rect 14327 13212 14372 13240
rect 14366 13200 14372 13212
rect 14424 13200 14430 13252
rect 15212 13249 15240 13280
rect 16393 13277 16405 13280
rect 16439 13308 16451 13311
rect 16666 13308 16672 13320
rect 16439 13280 16672 13308
rect 16439 13277 16451 13280
rect 16393 13271 16451 13277
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 15197 13243 15255 13249
rect 14476 13212 15148 13240
rect 9214 13172 9220 13184
rect 8036 13144 9220 13172
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 12897 13175 12955 13181
rect 12897 13141 12909 13175
rect 12943 13172 12955 13175
rect 13170 13172 13176 13184
rect 12943 13144 13176 13172
rect 12943 13141 12955 13144
rect 12897 13135 12955 13141
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 14476 13181 14504 13212
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 13780 13144 14473 13172
rect 13780 13132 13786 13144
rect 14461 13141 14473 13144
rect 14507 13141 14519 13175
rect 14461 13135 14519 13141
rect 14829 13175 14887 13181
rect 14829 13141 14841 13175
rect 14875 13172 14887 13175
rect 15010 13172 15016 13184
rect 14875 13144 15016 13172
rect 14875 13141 14887 13144
rect 14829 13135 14887 13141
rect 15010 13132 15016 13144
rect 15068 13132 15074 13184
rect 15120 13172 15148 13212
rect 15197 13209 15209 13243
rect 15243 13209 15255 13243
rect 16482 13240 16488 13252
rect 15197 13203 15255 13209
rect 15764 13212 16488 13240
rect 15764 13172 15792 13212
rect 16482 13200 16488 13212
rect 16540 13200 16546 13252
rect 16850 13200 16856 13252
rect 16908 13240 16914 13252
rect 17190 13243 17248 13249
rect 17190 13240 17202 13243
rect 16908 13212 17202 13240
rect 16908 13200 16914 13212
rect 17190 13209 17202 13212
rect 17236 13209 17248 13243
rect 17190 13203 17248 13209
rect 15930 13172 15936 13184
rect 15120 13144 15792 13172
rect 15891 13144 15936 13172
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 16301 13175 16359 13181
rect 16301 13141 16313 13175
rect 16347 13172 16359 13175
rect 17034 13172 17040 13184
rect 16347 13144 17040 13172
rect 16347 13141 16359 13144
rect 16301 13135 16359 13141
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 1104 13082 18860 13104
rect 1104 13030 6880 13082
rect 6932 13030 6944 13082
rect 6996 13030 7008 13082
rect 7060 13030 7072 13082
rect 7124 13030 7136 13082
rect 7188 13030 12811 13082
rect 12863 13030 12875 13082
rect 12927 13030 12939 13082
rect 12991 13030 13003 13082
rect 13055 13030 13067 13082
rect 13119 13030 18860 13082
rect 1104 13008 18860 13030
rect 2590 12968 2596 12980
rect 2551 12940 2596 12968
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 3786 12928 3792 12980
rect 3844 12968 3850 12980
rect 4341 12971 4399 12977
rect 4341 12968 4353 12971
rect 3844 12940 4353 12968
rect 3844 12928 3850 12940
rect 4341 12937 4353 12940
rect 4387 12968 4399 12971
rect 5166 12968 5172 12980
rect 4387 12940 5172 12968
rect 4387 12937 4399 12940
rect 4341 12931 4399 12937
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 5813 12971 5871 12977
rect 5813 12937 5825 12971
rect 5859 12968 5871 12971
rect 10410 12968 10416 12980
rect 5859 12940 9352 12968
rect 10371 12940 10416 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 4433 12903 4491 12909
rect 4433 12869 4445 12903
rect 4479 12900 4491 12903
rect 5626 12900 5632 12912
rect 4479 12872 5632 12900
rect 4479 12869 4491 12872
rect 4433 12863 4491 12869
rect 5626 12860 5632 12872
rect 5684 12860 5690 12912
rect 7558 12860 7564 12912
rect 7616 12900 7622 12912
rect 7616 12872 8248 12900
rect 7616 12860 7622 12872
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12801 2283 12835
rect 2225 12795 2283 12801
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12832 3295 12835
rect 4801 12835 4859 12841
rect 4801 12832 4813 12835
rect 3283 12804 4813 12832
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 4801 12801 4813 12804
rect 4847 12801 4859 12835
rect 4982 12832 4988 12844
rect 4943 12804 4988 12832
rect 4801 12795 4859 12801
rect 2240 12696 2268 12795
rect 2792 12764 2820 12795
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 5534 12832 5540 12844
rect 5092 12804 5540 12832
rect 5092 12764 5120 12804
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 5776 12804 6561 12832
rect 5776 12792 5782 12804
rect 6549 12801 6561 12804
rect 6595 12832 6607 12835
rect 6595 12804 6868 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 2792 12736 5120 12764
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12733 5227 12767
rect 5169 12727 5227 12733
rect 3694 12696 3700 12708
rect 2240 12668 3700 12696
rect 3694 12656 3700 12668
rect 3752 12656 3758 12708
rect 5184 12696 5212 12727
rect 5258 12724 5264 12776
rect 5316 12764 5322 12776
rect 5629 12767 5687 12773
rect 5629 12764 5641 12767
rect 5316 12736 5641 12764
rect 5316 12724 5322 12736
rect 5629 12733 5641 12736
rect 5675 12733 5687 12767
rect 5629 12727 5687 12733
rect 5997 12767 6055 12773
rect 5997 12733 6009 12767
rect 6043 12764 6055 12767
rect 6043 12736 6408 12764
rect 6043 12733 6055 12736
rect 5997 12727 6055 12733
rect 5350 12696 5356 12708
rect 5184 12668 5356 12696
rect 5350 12656 5356 12668
rect 5408 12696 5414 12708
rect 5718 12696 5724 12708
rect 5408 12668 5724 12696
rect 5408 12656 5414 12668
rect 5718 12656 5724 12668
rect 5776 12696 5782 12708
rect 6012 12696 6040 12727
rect 6380 12705 6408 12736
rect 6840 12705 6868 12804
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 8220 12841 8248 12872
rect 9324 12844 9352 12940
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 11885 12971 11943 12977
rect 11885 12937 11897 12971
rect 11931 12968 11943 12971
rect 13170 12968 13176 12980
rect 11931 12940 13176 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 13170 12928 13176 12940
rect 13228 12928 13234 12980
rect 15197 12971 15255 12977
rect 14568 12940 15148 12968
rect 9861 12903 9919 12909
rect 9861 12869 9873 12903
rect 9907 12900 9919 12903
rect 12342 12900 12348 12912
rect 9907 12872 12348 12900
rect 9907 12869 9919 12872
rect 9861 12863 9919 12869
rect 12342 12860 12348 12872
rect 12400 12860 12406 12912
rect 13081 12903 13139 12909
rect 13081 12869 13093 12903
rect 13127 12900 13139 12903
rect 14090 12900 14096 12912
rect 13127 12872 14096 12900
rect 13127 12869 13139 12872
rect 13081 12863 13139 12869
rect 14090 12860 14096 12872
rect 14148 12860 14154 12912
rect 7938 12835 7996 12841
rect 7938 12832 7950 12835
rect 7248 12804 7950 12832
rect 7248 12792 7254 12804
rect 7938 12801 7950 12804
rect 7984 12801 7996 12835
rect 7938 12795 7996 12801
rect 8205 12835 8263 12841
rect 8205 12801 8217 12835
rect 8251 12801 8263 12835
rect 9306 12832 9312 12844
rect 9219 12804 9312 12832
rect 8205 12795 8263 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12801 9735 12835
rect 10686 12832 10692 12844
rect 10647 12804 10692 12832
rect 9677 12795 9735 12801
rect 9030 12764 9036 12776
rect 8991 12736 9036 12764
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 9214 12724 9220 12776
rect 9272 12764 9278 12776
rect 9692 12764 9720 12795
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 9272 12736 9720 12764
rect 10796 12764 10824 12795
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 11054 12832 11060 12844
rect 10928 12804 10973 12832
rect 11015 12804 11060 12832
rect 10928 12792 10934 12804
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 11238 12792 11244 12844
rect 11296 12832 11302 12844
rect 11977 12835 12035 12841
rect 11977 12832 11989 12835
rect 11296 12804 11989 12832
rect 11296 12792 11302 12804
rect 11977 12801 11989 12804
rect 12023 12801 12035 12835
rect 11977 12795 12035 12801
rect 12526 12792 12532 12844
rect 12584 12832 12590 12844
rect 14568 12841 14596 12940
rect 15010 12900 15016 12912
rect 14844 12872 15016 12900
rect 14844 12841 14872 12872
rect 15010 12860 15016 12872
rect 15068 12860 15074 12912
rect 14553 12835 14611 12841
rect 14553 12832 14565 12835
rect 12584 12804 14565 12832
rect 12584 12792 12590 12804
rect 14553 12801 14565 12804
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12801 14795 12835
rect 14737 12795 14795 12801
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 12161 12767 12219 12773
rect 10796 12736 11560 12764
rect 9272 12724 9278 12736
rect 11532 12705 11560 12736
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 13357 12767 13415 12773
rect 12207 12736 13308 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 5776 12668 6040 12696
rect 6365 12699 6423 12705
rect 5776 12656 5782 12668
rect 6365 12665 6377 12699
rect 6411 12665 6423 12699
rect 6365 12659 6423 12665
rect 6825 12699 6883 12705
rect 6825 12665 6837 12699
rect 6871 12665 6883 12699
rect 6825 12659 6883 12665
rect 11517 12699 11575 12705
rect 11517 12665 11529 12699
rect 11563 12665 11575 12699
rect 11517 12659 11575 12665
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 12713 12699 12771 12705
rect 12713 12696 12725 12699
rect 12676 12668 12725 12696
rect 12676 12656 12682 12668
rect 12713 12665 12725 12668
rect 12759 12665 12771 12699
rect 13280 12696 13308 12736
rect 13357 12733 13369 12767
rect 13403 12764 13415 12767
rect 14366 12764 14372 12776
rect 13403 12736 14372 12764
rect 13403 12733 13415 12736
rect 13357 12727 13415 12733
rect 14366 12724 14372 12736
rect 14424 12724 14430 12776
rect 14752 12708 14780 12795
rect 14918 12792 14924 12844
rect 14976 12832 14982 12844
rect 15120 12832 15148 12940
rect 15197 12937 15209 12971
rect 15243 12968 15255 12971
rect 15286 12968 15292 12980
rect 15243 12940 15292 12968
rect 15243 12937 15255 12940
rect 15197 12931 15255 12937
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 16301 12971 16359 12977
rect 16301 12937 16313 12971
rect 16347 12968 16359 12971
rect 16758 12968 16764 12980
rect 16347 12940 16764 12968
rect 16347 12937 16359 12940
rect 16301 12931 16359 12937
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17129 12971 17187 12977
rect 17129 12968 17141 12971
rect 17092 12940 17141 12968
rect 17092 12928 17098 12940
rect 17129 12937 17141 12940
rect 17175 12937 17187 12971
rect 18230 12968 18236 12980
rect 18191 12940 18236 12968
rect 17129 12931 17187 12937
rect 18230 12928 18236 12940
rect 18288 12928 18294 12980
rect 15654 12832 15660 12844
rect 14976 12804 15021 12832
rect 15120 12804 15660 12832
rect 14976 12792 14982 12804
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 15820 12838 15878 12844
rect 15820 12804 15832 12838
rect 15866 12804 15878 12838
rect 15952 12838 16010 12844
rect 15952 12835 15964 12838
rect 15820 12798 15878 12804
rect 15935 12804 15964 12835
rect 15998 12804 16010 12838
rect 15935 12798 16010 12804
rect 16045 12835 16103 12841
rect 16045 12801 16057 12835
rect 16091 12832 16103 12835
rect 16390 12832 16396 12844
rect 16091 12804 16396 12832
rect 16091 12801 16103 12804
rect 15378 12724 15384 12776
rect 15436 12764 15442 12776
rect 15835 12764 15863 12798
rect 15436 12736 15863 12764
rect 15436 12724 15442 12736
rect 15935 12708 15963 12798
rect 16045 12795 16103 12801
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17770 12832 17776 12844
rect 17083 12804 17776 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 18046 12832 18052 12844
rect 18007 12804 18052 12832
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 16482 12724 16488 12776
rect 16540 12764 16546 12776
rect 17221 12767 17279 12773
rect 17221 12764 17233 12767
rect 16540 12736 17233 12764
rect 16540 12724 16546 12736
rect 17221 12733 17233 12736
rect 17267 12733 17279 12767
rect 17221 12727 17279 12733
rect 13722 12696 13728 12708
rect 13280 12668 13728 12696
rect 12713 12659 12771 12665
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 14734 12656 14740 12708
rect 14792 12656 14798 12708
rect 15930 12656 15936 12708
rect 15988 12656 15994 12708
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 2041 12631 2099 12637
rect 2041 12628 2053 12631
rect 2004 12600 2053 12628
rect 2004 12588 2010 12600
rect 2041 12597 2053 12600
rect 2087 12597 2099 12631
rect 3050 12628 3056 12640
rect 3011 12600 3056 12628
rect 2041 12591 2099 12597
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 4246 12588 4252 12640
rect 4304 12628 4310 12640
rect 5258 12628 5264 12640
rect 4304 12600 5264 12628
rect 4304 12588 4310 12600
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5442 12628 5448 12640
rect 5403 12600 5448 12628
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 5534 12588 5540 12640
rect 5592 12628 5598 12640
rect 5810 12628 5816 12640
rect 5592 12600 5816 12628
rect 5592 12588 5598 12600
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 16666 12628 16672 12640
rect 16627 12600 16672 12628
rect 16666 12588 16672 12600
rect 16724 12588 16730 12640
rect 1104 12538 18860 12560
rect 1104 12486 3915 12538
rect 3967 12486 3979 12538
rect 4031 12486 4043 12538
rect 4095 12486 4107 12538
rect 4159 12486 4171 12538
rect 4223 12486 9846 12538
rect 9898 12486 9910 12538
rect 9962 12486 9974 12538
rect 10026 12486 10038 12538
rect 10090 12486 10102 12538
rect 10154 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 15904 12538
rect 15956 12486 15968 12538
rect 16020 12486 16032 12538
rect 16084 12486 18860 12538
rect 1104 12464 18860 12486
rect 3694 12384 3700 12436
rect 3752 12424 3758 12436
rect 4801 12427 4859 12433
rect 4801 12424 4813 12427
rect 3752 12396 4813 12424
rect 3752 12384 3758 12396
rect 4801 12393 4813 12396
rect 4847 12393 4859 12427
rect 4801 12387 4859 12393
rect 5350 12384 5356 12436
rect 5408 12424 5414 12436
rect 5534 12424 5540 12436
rect 5408 12396 5540 12424
rect 5408 12384 5414 12396
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 5718 12424 5724 12436
rect 5679 12396 5724 12424
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 6270 12424 6276 12436
rect 6231 12396 6276 12424
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 7190 12424 7196 12436
rect 7151 12396 7196 12424
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 7558 12384 7564 12436
rect 7616 12424 7622 12436
rect 7653 12427 7711 12433
rect 7653 12424 7665 12427
rect 7616 12396 7665 12424
rect 7616 12384 7622 12396
rect 7653 12393 7665 12396
rect 7699 12393 7711 12427
rect 7653 12387 7711 12393
rect 10597 12427 10655 12433
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 10870 12424 10876 12436
rect 10643 12396 10876 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11885 12427 11943 12433
rect 11885 12393 11897 12427
rect 11931 12424 11943 12427
rect 12434 12424 12440 12436
rect 11931 12396 12440 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 14734 12424 14740 12436
rect 14695 12396 14740 12424
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 15378 12424 15384 12436
rect 15339 12396 15384 12424
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 17126 12384 17132 12436
rect 17184 12424 17190 12436
rect 18325 12427 18383 12433
rect 18325 12424 18337 12427
rect 17184 12396 18337 12424
rect 17184 12384 17190 12396
rect 18325 12393 18337 12396
rect 18371 12393 18383 12427
rect 18325 12387 18383 12393
rect 4522 12356 4528 12368
rect 4356 12328 4528 12356
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 1762 12220 1768 12232
rect 1719 12192 1768 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 1762 12180 1768 12192
rect 1820 12180 1826 12232
rect 1946 12229 1952 12232
rect 1940 12220 1952 12229
rect 1907 12192 1952 12220
rect 1940 12183 1952 12192
rect 1946 12180 1952 12183
rect 2004 12180 2010 12232
rect 4246 12220 4252 12232
rect 4207 12192 4252 12220
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 4356 12229 4384 12328
rect 4522 12316 4528 12328
rect 4580 12356 4586 12368
rect 6730 12356 6736 12368
rect 4580 12328 6736 12356
rect 4580 12316 4586 12328
rect 6730 12316 6736 12328
rect 6788 12316 6794 12368
rect 9030 12356 9036 12368
rect 7024 12328 9036 12356
rect 5258 12248 5264 12300
rect 5316 12288 5322 12300
rect 7024 12297 7052 12328
rect 9030 12316 9036 12328
rect 9088 12316 9094 12368
rect 11241 12359 11299 12365
rect 11241 12325 11253 12359
rect 11287 12356 11299 12359
rect 12250 12356 12256 12368
rect 11287 12328 12256 12356
rect 11287 12325 11299 12328
rect 11241 12319 11299 12325
rect 12250 12316 12256 12328
rect 12308 12316 12314 12368
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 5316 12260 5733 12288
rect 5316 12248 5322 12260
rect 5721 12257 5733 12260
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12257 7067 12291
rect 7282 12288 7288 12300
rect 7009 12251 7067 12257
rect 7116 12260 7288 12288
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12189 4399 12223
rect 4341 12183 4399 12189
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12220 5043 12223
rect 5074 12220 5080 12232
rect 5031 12192 5080 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 5169 12223 5227 12229
rect 5169 12189 5181 12223
rect 5215 12220 5227 12223
rect 5442 12220 5448 12232
rect 5215 12192 5448 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 5552 12192 6469 12220
rect 4525 12155 4583 12161
rect 4525 12121 4537 12155
rect 4571 12152 4583 12155
rect 5552 12152 5580 12192
rect 6457 12189 6469 12192
rect 6503 12189 6515 12223
rect 6457 12183 6515 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 7116 12220 7144 12260
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 8846 12248 8852 12300
rect 8904 12288 8910 12300
rect 8941 12291 8999 12297
rect 8941 12288 8953 12291
rect 8904 12260 8953 12288
rect 8904 12248 8910 12260
rect 8941 12257 8953 12260
rect 8987 12257 8999 12291
rect 9214 12288 9220 12300
rect 9175 12260 9220 12288
rect 8941 12251 8999 12257
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 12437 12291 12495 12297
rect 10244 12260 12296 12288
rect 6871 12192 7144 12220
rect 7193 12223 7251 12229
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 7650 12220 7656 12232
rect 7239 12192 7656 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7650 12180 7656 12192
rect 7708 12180 7714 12232
rect 4571 12124 5580 12152
rect 4571 12121 4583 12124
rect 4525 12115 4583 12121
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 5810 12152 5816 12164
rect 5684 12124 5816 12152
rect 5684 12112 5690 12124
rect 5810 12112 5816 12124
rect 5868 12152 5874 12164
rect 7561 12155 7619 12161
rect 7561 12152 7573 12155
rect 5868 12124 7573 12152
rect 5868 12112 5874 12124
rect 7561 12121 7573 12124
rect 7607 12121 7619 12155
rect 7561 12115 7619 12121
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 10244 12161 10272 12260
rect 10873 12223 10931 12229
rect 10873 12220 10885 12223
rect 10796 12192 10885 12220
rect 10229 12155 10287 12161
rect 10229 12152 10241 12155
rect 9088 12124 10241 12152
rect 9088 12112 9094 12124
rect 10229 12121 10241 12124
rect 10275 12121 10287 12155
rect 10229 12115 10287 12121
rect 10318 12112 10324 12164
rect 10376 12152 10382 12164
rect 10413 12155 10471 12161
rect 10413 12152 10425 12155
rect 10376 12124 10425 12152
rect 10376 12112 10382 12124
rect 10413 12121 10425 12124
rect 10459 12121 10471 12155
rect 10413 12115 10471 12121
rect 3053 12087 3111 12093
rect 3053 12053 3065 12087
rect 3099 12084 3111 12087
rect 3694 12084 3700 12096
rect 3099 12056 3700 12084
rect 3099 12053 3111 12056
rect 3053 12047 3111 12053
rect 3694 12044 3700 12056
rect 3752 12044 3758 12096
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 5997 12087 6055 12093
rect 5997 12084 6009 12087
rect 5592 12056 6009 12084
rect 5592 12044 5598 12056
rect 5997 12053 6009 12056
rect 6043 12084 6055 12087
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 6043 12056 6929 12084
rect 6043 12053 6055 12056
rect 5997 12047 6055 12053
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 6917 12047 6975 12053
rect 9306 12044 9312 12096
rect 9364 12084 9370 12096
rect 10796 12084 10824 12192
rect 10873 12189 10885 12192
rect 10919 12220 10931 12223
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 10919 12192 11529 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 11517 12189 11529 12192
rect 11563 12220 11575 12223
rect 11563 12192 11836 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 11057 12155 11115 12161
rect 11057 12121 11069 12155
rect 11103 12152 11115 12155
rect 11103 12124 11468 12152
rect 11103 12121 11115 12124
rect 11057 12115 11115 12121
rect 9364 12056 10824 12084
rect 11440 12084 11468 12124
rect 11606 12112 11612 12164
rect 11664 12152 11670 12164
rect 11701 12155 11759 12161
rect 11701 12152 11713 12155
rect 11664 12124 11713 12152
rect 11664 12112 11670 12124
rect 11701 12121 11713 12124
rect 11747 12121 11759 12155
rect 11808 12152 11836 12192
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12161 12223 12219 12229
rect 12161 12220 12173 12223
rect 12124 12192 12173 12220
rect 12124 12180 12130 12192
rect 12161 12189 12173 12192
rect 12207 12189 12219 12223
rect 12268 12220 12296 12260
rect 12437 12257 12449 12291
rect 12483 12288 12495 12291
rect 12526 12288 12532 12300
rect 12483 12260 12532 12288
rect 12483 12257 12495 12260
rect 12437 12251 12495 12257
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 16666 12288 16672 12300
rect 16316 12260 16672 12288
rect 12618 12220 12624 12232
rect 12268 12192 12624 12220
rect 12161 12183 12219 12189
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 13262 12180 13268 12232
rect 13320 12220 13326 12232
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 13320 12192 13461 12220
rect 13320 12180 13326 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13722 12220 13728 12232
rect 13683 12192 13728 12220
rect 13449 12183 13507 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 14384 12192 15025 12220
rect 14384 12161 14412 12192
rect 15013 12189 15025 12192
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 15654 12180 15660 12232
rect 15712 12220 15718 12232
rect 16025 12223 16083 12229
rect 16025 12220 16037 12223
rect 15712 12192 16037 12220
rect 15712 12180 15718 12192
rect 16025 12189 16037 12192
rect 16071 12189 16083 12223
rect 16206 12220 16212 12232
rect 16167 12192 16212 12220
rect 16025 12183 16083 12189
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 16316 12229 16344 12260
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12189 16359 12223
rect 16301 12183 16359 12189
rect 16390 12180 16396 12232
rect 16448 12220 16454 12232
rect 16448 12192 16493 12220
rect 16448 12180 16454 12192
rect 16758 12180 16764 12232
rect 16816 12220 16822 12232
rect 16942 12220 16948 12232
rect 16816 12192 16948 12220
rect 16816 12180 16822 12192
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 14369 12155 14427 12161
rect 14369 12152 14381 12155
rect 11808 12124 14381 12152
rect 11701 12115 11759 12121
rect 14369 12121 14381 12124
rect 14415 12121 14427 12155
rect 14369 12115 14427 12121
rect 14553 12155 14611 12161
rect 14553 12121 14565 12155
rect 14599 12152 14611 12155
rect 14734 12152 14740 12164
rect 14599 12124 14740 12152
rect 14599 12121 14611 12124
rect 14553 12115 14611 12121
rect 14734 12112 14740 12124
rect 14792 12112 14798 12164
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12152 15255 12155
rect 15286 12152 15292 12164
rect 15243 12124 15292 12152
rect 15243 12121 15255 12124
rect 15197 12115 15255 12121
rect 15286 12112 15292 12124
rect 15344 12112 15350 12164
rect 16669 12155 16727 12161
rect 16669 12121 16681 12155
rect 16715 12152 16727 12155
rect 17190 12155 17248 12161
rect 17190 12152 17202 12155
rect 16715 12124 17202 12152
rect 16715 12121 16727 12124
rect 16669 12115 16727 12121
rect 17190 12121 17202 12124
rect 17236 12121 17248 12155
rect 17190 12115 17248 12121
rect 12710 12084 12716 12096
rect 11440 12056 12716 12084
rect 9364 12044 9370 12056
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 13228 12056 13277 12084
rect 13228 12044 13234 12056
rect 13265 12053 13277 12056
rect 13311 12053 13323 12087
rect 13265 12047 13323 12053
rect 13633 12087 13691 12093
rect 13633 12053 13645 12087
rect 13679 12084 13691 12087
rect 14458 12084 14464 12096
rect 13679 12056 14464 12084
rect 13679 12053 13691 12056
rect 13633 12047 13691 12053
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 1104 11994 18860 12016
rect 1104 11942 6880 11994
rect 6932 11942 6944 11994
rect 6996 11942 7008 11994
rect 7060 11942 7072 11994
rect 7124 11942 7136 11994
rect 7188 11942 12811 11994
rect 12863 11942 12875 11994
rect 12927 11942 12939 11994
rect 12991 11942 13003 11994
rect 13055 11942 13067 11994
rect 13119 11942 18860 11994
rect 1104 11920 18860 11942
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 5810 11880 5816 11892
rect 5767 11852 5816 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 5902 11840 5908 11892
rect 5960 11880 5966 11892
rect 8757 11883 8815 11889
rect 5960 11852 7972 11880
rect 5960 11840 5966 11852
rect 2124 11815 2182 11821
rect 2124 11781 2136 11815
rect 2170 11812 2182 11815
rect 3050 11812 3056 11824
rect 2170 11784 3056 11812
rect 2170 11781 2182 11784
rect 2124 11775 2182 11781
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 4056 11815 4114 11821
rect 4056 11781 4068 11815
rect 4102 11812 4114 11815
rect 6270 11812 6276 11824
rect 4102 11784 6276 11812
rect 4102 11781 4114 11784
rect 4056 11775 4114 11781
rect 6270 11772 6276 11784
rect 6328 11772 6334 11824
rect 7009 11815 7067 11821
rect 7009 11781 7021 11815
rect 7055 11812 7067 11815
rect 7644 11815 7702 11821
rect 7644 11812 7656 11815
rect 7055 11784 7656 11812
rect 7055 11781 7067 11784
rect 7009 11775 7067 11781
rect 7644 11781 7656 11784
rect 7690 11812 7702 11815
rect 7834 11812 7840 11824
rect 7690 11784 7840 11812
rect 7690 11781 7702 11784
rect 7644 11775 7702 11781
rect 7834 11772 7840 11784
rect 7892 11772 7898 11824
rect 7944 11812 7972 11852
rect 8757 11849 8769 11883
rect 8803 11880 8815 11883
rect 13722 11880 13728 11892
rect 8803 11852 13728 11880
rect 8803 11849 8815 11852
rect 8757 11843 8815 11849
rect 13722 11840 13728 11852
rect 13780 11840 13786 11892
rect 13440 11815 13498 11821
rect 7944 11784 9628 11812
rect 9600 11756 9628 11784
rect 13440 11781 13452 11815
rect 13486 11812 13498 11815
rect 13538 11812 13544 11824
rect 13486 11784 13544 11812
rect 13486 11781 13498 11784
rect 13440 11775 13498 11781
rect 13538 11772 13544 11784
rect 13596 11772 13602 11824
rect 14918 11772 14924 11824
rect 14976 11812 14982 11824
rect 16301 11815 16359 11821
rect 14976 11784 16068 11812
rect 14976 11772 14982 11784
rect 1854 11744 1860 11756
rect 1815 11716 1860 11744
rect 1854 11704 1860 11716
rect 1912 11704 1918 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6546 11744 6552 11756
rect 5859 11716 6552 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 6730 11744 6736 11756
rect 6691 11716 6736 11744
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11744 7435 11747
rect 7466 11744 7472 11756
rect 7423 11716 7472 11744
rect 7423 11713 7435 11716
rect 7377 11707 7435 11713
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 9033 11747 9091 11753
rect 9033 11713 9045 11747
rect 9079 11744 9091 11747
rect 9122 11744 9128 11756
rect 9079 11716 9128 11744
rect 9079 11713 9091 11716
rect 9033 11707 9091 11713
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 9306 11753 9312 11756
rect 9300 11707 9312 11753
rect 9364 11744 9370 11756
rect 9364 11716 9400 11744
rect 9306 11704 9312 11707
rect 9364 11704 9370 11716
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 9640 11716 10701 11744
rect 9640 11704 9646 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11713 10931 11747
rect 10873 11707 10931 11713
rect 3786 11676 3792 11688
rect 3747 11648 3792 11676
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6144 11648 6837 11676
rect 6144 11636 6150 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11645 7067 11679
rect 10888 11676 10916 11707
rect 10962 11704 10968 11756
rect 11020 11744 11026 11756
rect 11773 11747 11831 11753
rect 11773 11744 11785 11747
rect 11020 11716 11785 11744
rect 11020 11704 11026 11716
rect 11773 11713 11785 11716
rect 11819 11713 11831 11747
rect 11773 11707 11831 11713
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 15010 11744 15016 11756
rect 12676 11716 15016 11744
rect 12676 11704 12682 11716
rect 15010 11704 15016 11716
rect 15068 11704 15074 11756
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11713 15255 11747
rect 15654 11744 15660 11756
rect 15615 11716 15660 11744
rect 15197 11707 15255 11713
rect 11330 11676 11336 11688
rect 10888 11648 11336 11676
rect 7009 11639 7067 11645
rect 1394 11608 1400 11620
rect 1355 11580 1400 11608
rect 1394 11568 1400 11580
rect 1452 11568 1458 11620
rect 4982 11568 4988 11620
rect 5040 11608 5046 11620
rect 5040 11580 6592 11608
rect 5040 11568 5046 11580
rect 3234 11540 3240 11552
rect 3195 11512 3240 11540
rect 3234 11500 3240 11512
rect 3292 11500 3298 11552
rect 5166 11540 5172 11552
rect 5127 11512 5172 11540
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 6564 11540 6592 11580
rect 6638 11568 6644 11620
rect 6696 11608 6702 11620
rect 7024 11608 7052 11639
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11480 11648 11529 11676
rect 11480 11636 11486 11648
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 6696 11580 7052 11608
rect 6696 11568 6702 11580
rect 7558 11540 7564 11552
rect 6564 11512 7564 11540
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 10413 11543 10471 11549
rect 10413 11540 10425 11543
rect 10376 11512 10425 11540
rect 10376 11500 10382 11512
rect 10413 11509 10425 11512
rect 10459 11509 10471 11543
rect 10413 11503 10471 11509
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 10836 11512 11069 11540
rect 10836 11500 10842 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 11057 11503 11115 11509
rect 12710 11500 12716 11552
rect 12768 11540 12774 11552
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12768 11512 12909 11540
rect 12768 11500 12774 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 13188 11540 13216 11639
rect 14642 11636 14648 11688
rect 14700 11676 14706 11688
rect 15212 11676 15240 11707
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 16040 11753 16068 11784
rect 16301 11781 16313 11815
rect 16347 11812 16359 11815
rect 17006 11815 17064 11821
rect 17006 11812 17018 11815
rect 16347 11784 17018 11812
rect 16347 11781 16359 11784
rect 16301 11775 16359 11781
rect 17006 11781 17018 11784
rect 17052 11781 17064 11815
rect 17006 11775 17064 11781
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11744 16083 11747
rect 16390 11744 16396 11756
rect 16071 11716 16396 11744
rect 16071 11713 16083 11716
rect 16025 11707 16083 11713
rect 14700 11648 15240 11676
rect 15381 11679 15439 11685
rect 14700 11636 14706 11648
rect 15381 11645 15393 11679
rect 15427 11676 15439 11679
rect 15856 11676 15884 11707
rect 15427 11648 15884 11676
rect 15948 11676 15976 11707
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 16114 11676 16120 11688
rect 15948 11648 16120 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 16758 11676 16764 11688
rect 16719 11648 16764 11676
rect 16758 11636 16764 11648
rect 16816 11636 16822 11688
rect 14274 11540 14280 11552
rect 13188 11512 14280 11540
rect 12897 11503 12955 11509
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 14458 11500 14464 11552
rect 14516 11540 14522 11552
rect 14553 11543 14611 11549
rect 14553 11540 14565 11543
rect 14516 11512 14565 11540
rect 14516 11500 14522 11512
rect 14553 11509 14565 11512
rect 14599 11540 14611 11543
rect 16298 11540 16304 11552
rect 14599 11512 16304 11540
rect 14599 11509 14611 11512
rect 14553 11503 14611 11509
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 17770 11540 17776 11552
rect 16632 11512 17776 11540
rect 16632 11500 16638 11512
rect 17770 11500 17776 11512
rect 17828 11540 17834 11552
rect 18141 11543 18199 11549
rect 18141 11540 18153 11543
rect 17828 11512 18153 11540
rect 17828 11500 17834 11512
rect 18141 11509 18153 11512
rect 18187 11509 18199 11543
rect 18141 11503 18199 11509
rect 1104 11450 18860 11472
rect 1104 11398 3915 11450
rect 3967 11398 3979 11450
rect 4031 11398 4043 11450
rect 4095 11398 4107 11450
rect 4159 11398 4171 11450
rect 4223 11398 9846 11450
rect 9898 11398 9910 11450
rect 9962 11398 9974 11450
rect 10026 11398 10038 11450
rect 10090 11398 10102 11450
rect 10154 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 15904 11450
rect 15956 11398 15968 11450
rect 16020 11398 16032 11450
rect 16084 11398 18860 11450
rect 1104 11376 18860 11398
rect 3234 11296 3240 11348
rect 3292 11336 3298 11348
rect 3973 11339 4031 11345
rect 3973 11336 3985 11339
rect 3292 11308 3985 11336
rect 3292 11296 3298 11308
rect 3973 11305 3985 11308
rect 4019 11305 4031 11339
rect 3973 11299 4031 11305
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 5902 11336 5908 11348
rect 4663 11308 5908 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 3421 11271 3479 11277
rect 3421 11237 3433 11271
rect 3467 11268 3479 11271
rect 4154 11268 4160 11280
rect 3467 11240 4160 11268
rect 3467 11237 3479 11240
rect 3421 11231 3479 11237
rect 4154 11228 4160 11240
rect 4212 11228 4218 11280
rect 4632 11268 4660 11299
rect 5902 11296 5908 11308
rect 5960 11296 5966 11348
rect 5994 11296 6000 11348
rect 6052 11336 6058 11348
rect 6730 11336 6736 11348
rect 6052 11308 6736 11336
rect 6052 11296 6058 11308
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 9306 11336 9312 11348
rect 8619 11308 9312 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 10962 11336 10968 11348
rect 10923 11308 10968 11336
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 11330 11296 11336 11348
rect 11388 11336 11394 11348
rect 12161 11339 12219 11345
rect 12161 11336 12173 11339
rect 11388 11308 12173 11336
rect 11388 11296 11394 11308
rect 12161 11305 12173 11308
rect 12207 11305 12219 11339
rect 16114 11336 16120 11348
rect 16075 11308 16120 11336
rect 12161 11299 12219 11305
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 5166 11268 5172 11280
rect 4356 11240 4660 11268
rect 5127 11240 5172 11268
rect 2130 11160 2136 11212
rect 2188 11200 2194 11212
rect 2593 11203 2651 11209
rect 2593 11200 2605 11203
rect 2188 11172 2605 11200
rect 2188 11160 2194 11172
rect 2593 11169 2605 11172
rect 2639 11200 2651 11203
rect 4356 11200 4384 11240
rect 5166 11228 5172 11240
rect 5224 11228 5230 11280
rect 5261 11271 5319 11277
rect 5261 11237 5273 11271
rect 5307 11237 5319 11271
rect 5261 11231 5319 11237
rect 5276 11200 5304 11231
rect 7466 11228 7472 11280
rect 7524 11268 7530 11280
rect 7745 11271 7803 11277
rect 7745 11268 7757 11271
rect 7524 11240 7757 11268
rect 7524 11228 7530 11240
rect 7745 11237 7757 11240
rect 7791 11268 7803 11271
rect 8846 11268 8852 11280
rect 7791 11240 8852 11268
rect 7791 11237 7803 11240
rect 7745 11231 7803 11237
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 9585 11271 9643 11277
rect 9585 11237 9597 11271
rect 9631 11237 9643 11271
rect 9585 11231 9643 11237
rect 15841 11271 15899 11277
rect 15841 11237 15853 11271
rect 15887 11268 15899 11271
rect 16206 11268 16212 11280
rect 15887 11240 16212 11268
rect 15887 11237 15899 11240
rect 15841 11231 15899 11237
rect 2639 11172 4384 11200
rect 4448 11172 5304 11200
rect 2639 11169 2651 11172
rect 2593 11163 2651 11169
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2406 11132 2412 11144
rect 2367 11104 2412 11132
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3283 11104 3924 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3694 11024 3700 11076
rect 3752 11064 3758 11076
rect 3789 11067 3847 11073
rect 3789 11064 3801 11067
rect 3752 11036 3801 11064
rect 3752 11024 3758 11036
rect 3789 11033 3801 11036
rect 3835 11033 3847 11067
rect 3789 11027 3847 11033
rect 2225 10999 2283 11005
rect 2225 10965 2237 10999
rect 2271 10996 2283 10999
rect 2314 10996 2320 11008
rect 2271 10968 2320 10996
rect 2271 10965 2283 10968
rect 2225 10959 2283 10965
rect 2314 10956 2320 10968
rect 2372 10956 2378 11008
rect 3896 10996 3924 11104
rect 4005 11067 4063 11073
rect 4005 11033 4017 11067
rect 4051 11064 4063 11067
rect 4448 11064 4476 11172
rect 5350 11160 5356 11212
rect 5408 11200 5414 11212
rect 5408 11172 6132 11200
rect 5408 11160 5414 11172
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 5261 11135 5319 11141
rect 4571 11104 5212 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 4982 11064 4988 11076
rect 4051 11036 4476 11064
rect 4943 11036 4988 11064
rect 4051 11033 4063 11036
rect 4005 11027 4063 11033
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 5184 11064 5212 11104
rect 5261 11101 5273 11135
rect 5307 11132 5319 11135
rect 5368 11132 5396 11160
rect 5534 11132 5540 11144
rect 5307 11104 5396 11132
rect 5495 11104 5540 11132
rect 5307 11101 5319 11104
rect 5261 11095 5319 11101
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11132 5779 11135
rect 5994 11132 6000 11144
rect 5767 11104 6000 11132
rect 5767 11101 5779 11104
rect 5721 11095 5779 11101
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 6104 11132 6132 11172
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 9600 11200 9628 11231
rect 16206 11228 16212 11240
rect 16264 11228 16270 11280
rect 7616 11172 7880 11200
rect 7616 11160 7622 11172
rect 6730 11132 6736 11144
rect 6104 11104 6736 11132
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11132 7435 11135
rect 7650 11132 7656 11144
rect 7423 11104 7656 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 7852 11141 7880 11172
rect 9140 11172 9628 11200
rect 10229 11203 10287 11209
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11132 7895 11135
rect 8110 11132 8116 11144
rect 7883 11104 8116 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 9140 11141 9168 11172
rect 10229 11169 10241 11203
rect 10275 11200 10287 11203
rect 12158 11200 12164 11212
rect 10275 11172 12164 11200
rect 10275 11169 10287 11172
rect 10229 11163 10287 11169
rect 12158 11160 12164 11172
rect 12216 11200 12222 11212
rect 12713 11203 12771 11209
rect 12713 11200 12725 11203
rect 12216 11172 12725 11200
rect 12216 11160 12222 11172
rect 12713 11169 12725 11172
rect 12759 11169 12771 11203
rect 12713 11163 12771 11169
rect 16482 11160 16488 11212
rect 16540 11200 16546 11212
rect 16669 11203 16727 11209
rect 16669 11200 16681 11203
rect 16540 11172 16681 11200
rect 16540 11160 16546 11172
rect 16669 11169 16681 11172
rect 16715 11169 16727 11203
rect 16669 11163 16727 11169
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11132 8447 11135
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8435 11104 8953 11132
rect 8435 11101 8447 11104
rect 8389 11095 8447 11101
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9582 11132 9588 11144
rect 9355 11104 9588 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9824 11104 9965 11132
rect 9824 11092 9830 11104
rect 9953 11101 9965 11104
rect 9999 11132 10011 11135
rect 10594 11132 10600 11144
rect 9999 11104 10600 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 10778 11132 10784 11144
rect 10739 11104 10784 11132
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 15562 11132 15568 11144
rect 12575 11104 15568 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 16574 11132 16580 11144
rect 16535 11104 16580 11132
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 17865 11135 17923 11141
rect 17865 11101 17877 11135
rect 17911 11132 17923 11135
rect 18322 11132 18328 11144
rect 17911 11104 18328 11132
rect 17911 11101 17923 11104
rect 17865 11095 17923 11101
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 5629 11067 5687 11073
rect 5184 11036 5580 11064
rect 5552 11008 5580 11036
rect 5629 11033 5641 11067
rect 5675 11064 5687 11067
rect 7132 11067 7190 11073
rect 5675 11036 7052 11064
rect 5675 11033 5687 11036
rect 5629 11027 5687 11033
rect 4157 10999 4215 11005
rect 4157 10996 4169 10999
rect 3896 10968 4169 10996
rect 4157 10965 4169 10968
rect 4203 10965 4215 10999
rect 4157 10959 4215 10965
rect 5534 10956 5540 11008
rect 5592 10956 5598 11008
rect 7024 10996 7052 11036
rect 7132 11033 7144 11067
rect 7178 11064 7190 11067
rect 7558 11064 7564 11076
rect 7178 11036 7564 11064
rect 7178 11033 7190 11036
rect 7132 11027 7190 11033
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 10045 11067 10103 11073
rect 10045 11033 10057 11067
rect 10091 11064 10103 11067
rect 10318 11064 10324 11076
rect 10091 11036 10324 11064
rect 10091 11033 10103 11036
rect 10045 11027 10103 11033
rect 10318 11024 10324 11036
rect 10376 11024 10382 11076
rect 11146 11024 11152 11076
rect 11204 11064 11210 11076
rect 11333 11067 11391 11073
rect 11333 11064 11345 11067
rect 11204 11036 11345 11064
rect 11204 11024 11210 11036
rect 11333 11033 11345 11036
rect 11379 11064 11391 11067
rect 12066 11064 12072 11076
rect 11379 11036 12072 11064
rect 11379 11033 11391 11036
rect 11333 11027 11391 11033
rect 12066 11024 12072 11036
rect 12124 11024 12130 11076
rect 12621 11067 12679 11073
rect 12621 11033 12633 11067
rect 12667 11064 12679 11067
rect 12710 11064 12716 11076
rect 12667 11036 12716 11064
rect 12667 11033 12679 11036
rect 12621 11027 12679 11033
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 13262 11064 13268 11076
rect 13223 11036 13268 11064
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 13446 11064 13452 11076
rect 13407 11036 13452 11064
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 13998 11024 14004 11076
rect 14056 11064 14062 11076
rect 14550 11064 14556 11076
rect 14056 11036 14556 11064
rect 14056 11024 14062 11036
rect 14550 11024 14556 11036
rect 14608 11064 14614 11076
rect 14737 11067 14795 11073
rect 14737 11064 14749 11067
rect 14608 11036 14749 11064
rect 14608 11024 14614 11036
rect 14737 11033 14749 11036
rect 14783 11033 14795 11067
rect 14918 11064 14924 11076
rect 14879 11036 14924 11064
rect 14737 11027 14795 11033
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 15010 11024 15016 11076
rect 15068 11064 15074 11076
rect 15473 11067 15531 11073
rect 15473 11064 15485 11067
rect 15068 11036 15485 11064
rect 15068 11024 15074 11036
rect 15473 11033 15485 11036
rect 15519 11033 15531 11067
rect 15654 11064 15660 11076
rect 15615 11036 15660 11064
rect 15473 11027 15531 11033
rect 15654 11024 15660 11036
rect 15712 11024 15718 11076
rect 16298 11024 16304 11076
rect 16356 11064 16362 11076
rect 16485 11067 16543 11073
rect 16485 11064 16497 11067
rect 16356 11036 16497 11064
rect 16356 11024 16362 11036
rect 16485 11033 16497 11036
rect 16531 11033 16543 11067
rect 16485 11027 16543 11033
rect 17497 11067 17555 11073
rect 17497 11033 17509 11067
rect 17543 11064 17555 11067
rect 17586 11064 17592 11076
rect 17543 11036 17592 11064
rect 17543 11033 17555 11036
rect 17497 11027 17555 11033
rect 17586 11024 17592 11036
rect 17644 11024 17650 11076
rect 7282 10996 7288 11008
rect 7024 10968 7288 10996
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 10962 10956 10968 11008
rect 11020 10996 11026 11008
rect 11425 10999 11483 11005
rect 11425 10996 11437 10999
rect 11020 10968 11437 10996
rect 11020 10956 11026 10968
rect 11425 10965 11437 10968
rect 11471 10996 11483 10999
rect 12250 10996 12256 11008
rect 11471 10968 12256 10996
rect 11471 10965 11483 10968
rect 11425 10959 11483 10965
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 17862 10956 17868 11008
rect 17920 10996 17926 11008
rect 18141 10999 18199 11005
rect 18141 10996 18153 10999
rect 17920 10968 18153 10996
rect 17920 10956 17926 10968
rect 18141 10965 18153 10968
rect 18187 10965 18199 10999
rect 18141 10959 18199 10965
rect 1104 10906 18860 10928
rect 1104 10854 6880 10906
rect 6932 10854 6944 10906
rect 6996 10854 7008 10906
rect 7060 10854 7072 10906
rect 7124 10854 7136 10906
rect 7188 10854 12811 10906
rect 12863 10854 12875 10906
rect 12927 10854 12939 10906
rect 12991 10854 13003 10906
rect 13055 10854 13067 10906
rect 13119 10854 18860 10906
rect 1104 10832 18860 10854
rect 5074 10752 5080 10804
rect 5132 10792 5138 10804
rect 5721 10795 5779 10801
rect 5721 10792 5733 10795
rect 5132 10764 5733 10792
rect 5132 10752 5138 10764
rect 5721 10761 5733 10764
rect 5767 10792 5779 10795
rect 9766 10792 9772 10804
rect 5767 10764 8524 10792
rect 9727 10764 9772 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 3786 10684 3792 10736
rect 3844 10724 3850 10736
rect 5994 10724 6000 10736
rect 3844 10696 6000 10724
rect 3844 10684 3850 10696
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 1854 10656 1860 10668
rect 1811 10628 1860 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 1854 10616 1860 10628
rect 1912 10616 1918 10668
rect 2038 10665 2044 10668
rect 2032 10619 2044 10665
rect 2096 10656 2102 10668
rect 3896 10665 3924 10696
rect 5994 10684 6000 10696
rect 6052 10684 6058 10736
rect 6917 10727 6975 10733
rect 6917 10693 6929 10727
rect 6963 10724 6975 10727
rect 7466 10724 7472 10736
rect 6963 10696 7472 10724
rect 6963 10693 6975 10696
rect 6917 10687 6975 10693
rect 7466 10684 7472 10696
rect 7524 10684 7530 10736
rect 7561 10727 7619 10733
rect 7561 10693 7573 10727
rect 7607 10724 7619 10727
rect 7742 10724 7748 10736
rect 7607 10696 7748 10724
rect 7607 10693 7619 10696
rect 7561 10687 7619 10693
rect 7742 10684 7748 10696
rect 7800 10724 7806 10736
rect 8496 10724 8524 10764
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 11146 10792 11152 10804
rect 9876 10764 11152 10792
rect 9876 10724 9904 10764
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 13170 10752 13176 10804
rect 13228 10752 13234 10804
rect 14274 10752 14280 10804
rect 14332 10792 14338 10804
rect 16117 10795 16175 10801
rect 16117 10792 16129 10795
rect 14332 10764 16129 10792
rect 14332 10752 14338 10764
rect 16117 10761 16129 10764
rect 16163 10761 16175 10795
rect 16117 10755 16175 10761
rect 7800 10696 8064 10724
rect 8496 10696 9904 10724
rect 7800 10684 7806 10696
rect 4154 10665 4160 10668
rect 3881 10659 3939 10665
rect 2096 10628 2132 10656
rect 2038 10616 2044 10619
rect 2096 10616 2102 10628
rect 3881 10625 3893 10659
rect 3927 10625 3939 10659
rect 4148 10656 4160 10665
rect 4115 10628 4160 10656
rect 3881 10619 3939 10625
rect 4148 10619 4160 10628
rect 4154 10616 4160 10619
rect 4212 10616 4218 10668
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5592 10628 5641 10656
rect 5592 10616 5598 10628
rect 5629 10625 5641 10628
rect 5675 10656 5687 10659
rect 7282 10656 7288 10668
rect 5675 10628 6684 10656
rect 7243 10628 7288 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 6656 10532 6684 10628
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10625 7435 10659
rect 7834 10656 7840 10668
rect 7795 10628 7840 10656
rect 7377 10619 7435 10625
rect 7392 10588 7420 10619
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 8036 10665 8064 10696
rect 10686 10684 10692 10736
rect 10744 10724 10750 10736
rect 10965 10727 11023 10733
rect 10965 10724 10977 10727
rect 10744 10696 10977 10724
rect 10744 10684 10750 10696
rect 10965 10693 10977 10696
rect 11011 10693 11023 10727
rect 10965 10687 11023 10693
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 11977 10727 12035 10733
rect 11977 10724 11989 10727
rect 11388 10696 11989 10724
rect 11388 10684 11394 10696
rect 11977 10693 11989 10696
rect 12023 10693 12035 10727
rect 13188 10724 13216 10752
rect 11977 10687 12035 10693
rect 13004 10696 13216 10724
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 9674 10656 9680 10668
rect 9635 10628 9680 10656
rect 8021 10619 8079 10625
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10284 10628 10609 10656
rect 10284 10616 10290 10628
rect 10597 10625 10609 10628
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 11882 10656 11888 10668
rect 11572 10628 11888 10656
rect 11572 10616 11578 10628
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 7466 10588 7472 10600
rect 7392 10560 7472 10588
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9824 10560 9873 10588
rect 9824 10548 9830 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 11974 10548 11980 10600
rect 12032 10588 12038 10600
rect 12176 10588 12204 10619
rect 12250 10616 12256 10668
rect 12308 10656 12314 10668
rect 13004 10665 13032 10696
rect 13446 10684 13452 10736
rect 13504 10724 13510 10736
rect 16025 10727 16083 10733
rect 16025 10724 16037 10727
rect 13504 10696 16037 10724
rect 13504 10684 13510 10696
rect 16025 10693 16037 10696
rect 16071 10693 16083 10727
rect 16025 10687 16083 10693
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12308 10628 12817 10656
rect 12308 10616 12314 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 14090 10656 14096 10668
rect 13219 10628 14096 10656
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 12032 10560 12204 10588
rect 12032 10548 12038 10560
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 13096 10588 13124 10619
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 14274 10656 14280 10668
rect 14235 10628 14280 10656
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 14550 10665 14556 10668
rect 14544 10619 14556 10665
rect 14608 10656 14614 10668
rect 16132 10656 16160 10755
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 14608 10628 14644 10656
rect 16132 10628 16681 10656
rect 14550 10616 14556 10619
rect 14608 10616 14614 10628
rect 16669 10625 16681 10628
rect 16715 10656 16727 10659
rect 16758 10656 16764 10668
rect 16715 10628 16764 10656
rect 16715 10625 16727 10628
rect 16669 10619 16727 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 16942 10665 16948 10668
rect 16936 10619 16948 10665
rect 17000 10656 17006 10668
rect 17000 10628 17036 10656
rect 16942 10616 16948 10619
rect 17000 10616 17006 10628
rect 12676 10560 13124 10588
rect 13449 10591 13507 10597
rect 12676 10548 12682 10560
rect 13449 10557 13461 10591
rect 13495 10588 13507 10591
rect 13538 10588 13544 10600
rect 13495 10560 13544 10588
rect 13495 10557 13507 10560
rect 13449 10551 13507 10557
rect 13538 10548 13544 10560
rect 13596 10548 13602 10600
rect 6638 10480 6644 10532
rect 6696 10520 6702 10532
rect 6733 10523 6791 10529
rect 6733 10520 6745 10523
rect 6696 10492 6745 10520
rect 6696 10480 6702 10492
rect 6733 10489 6745 10492
rect 6779 10489 6791 10523
rect 7558 10520 7564 10532
rect 7519 10492 7564 10520
rect 6733 10483 6791 10489
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 11149 10523 11207 10529
rect 11149 10489 11161 10523
rect 11195 10520 11207 10523
rect 13262 10520 13268 10532
rect 11195 10492 13268 10520
rect 11195 10489 11207 10492
rect 11149 10483 11207 10489
rect 13262 10480 13268 10492
rect 13320 10480 13326 10532
rect 15470 10480 15476 10532
rect 15528 10520 15534 10532
rect 15654 10520 15660 10532
rect 15528 10492 15660 10520
rect 15528 10480 15534 10492
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 3145 10455 3203 10461
rect 3145 10452 3157 10455
rect 2924 10424 3157 10452
rect 2924 10412 2930 10424
rect 3145 10421 3157 10424
rect 3191 10421 3203 10455
rect 5258 10452 5264 10464
rect 5219 10424 5264 10452
rect 3145 10415 3203 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 7837 10455 7895 10461
rect 7837 10421 7849 10455
rect 7883 10452 7895 10455
rect 7926 10452 7932 10464
rect 7883 10424 7932 10452
rect 7883 10421 7895 10424
rect 7837 10415 7895 10421
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 9309 10455 9367 10461
rect 9309 10421 9321 10455
rect 9355 10452 9367 10455
rect 9582 10452 9588 10464
rect 9355 10424 9588 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 10410 10452 10416 10464
rect 10371 10424 10416 10452
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 12161 10455 12219 10461
rect 12161 10421 12173 10455
rect 12207 10452 12219 10455
rect 12250 10452 12256 10464
rect 12207 10424 12256 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 14001 10455 14059 10461
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 15378 10452 15384 10464
rect 14047 10424 15384 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 16206 10412 16212 10464
rect 16264 10452 16270 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 16264 10424 18061 10452
rect 16264 10412 16270 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 1104 10362 18860 10384
rect 1104 10310 3915 10362
rect 3967 10310 3979 10362
rect 4031 10310 4043 10362
rect 4095 10310 4107 10362
rect 4159 10310 4171 10362
rect 4223 10310 9846 10362
rect 9898 10310 9910 10362
rect 9962 10310 9974 10362
rect 10026 10310 10038 10362
rect 10090 10310 10102 10362
rect 10154 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 15904 10362
rect 15956 10310 15968 10362
rect 16020 10310 16032 10362
rect 16084 10310 18860 10362
rect 1104 10288 18860 10310
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 2133 10251 2191 10257
rect 2133 10248 2145 10251
rect 2096 10220 2145 10248
rect 2096 10208 2102 10220
rect 2133 10217 2145 10220
rect 2179 10217 2191 10251
rect 2133 10211 2191 10217
rect 2406 10208 2412 10260
rect 2464 10248 2470 10260
rect 2685 10251 2743 10257
rect 2685 10248 2697 10251
rect 2464 10220 2697 10248
rect 2464 10208 2470 10220
rect 2685 10217 2697 10220
rect 2731 10217 2743 10251
rect 5350 10248 5356 10260
rect 5263 10220 5356 10248
rect 2685 10211 2743 10217
rect 5350 10208 5356 10220
rect 5408 10248 5414 10260
rect 14182 10248 14188 10260
rect 5408 10220 14188 10248
rect 5408 10208 5414 10220
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 18325 10251 18383 10257
rect 18325 10248 18337 10251
rect 18104 10220 18337 10248
rect 18104 10208 18110 10220
rect 18325 10217 18337 10220
rect 18371 10217 18383 10251
rect 18325 10211 18383 10217
rect 7742 10140 7748 10192
rect 7800 10180 7806 10192
rect 7929 10183 7987 10189
rect 7929 10180 7941 10183
rect 7800 10152 7941 10180
rect 7800 10140 7806 10152
rect 7929 10149 7941 10152
rect 7975 10149 7987 10183
rect 7929 10143 7987 10149
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 3329 10115 3387 10121
rect 3329 10112 3341 10115
rect 3200 10084 3341 10112
rect 3200 10072 3206 10084
rect 3329 10081 3341 10084
rect 3375 10112 3387 10115
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 3375 10084 3985 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 3973 10081 3985 10084
rect 4019 10081 4031 10115
rect 3973 10075 4031 10081
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10112 10563 10115
rect 11422 10112 11428 10124
rect 10551 10084 11428 10112
rect 10551 10081 10563 10084
rect 10505 10075 10563 10081
rect 11422 10072 11428 10084
rect 11480 10112 11486 10124
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 11480 10084 12265 10112
rect 11480 10072 11486 10084
rect 12253 10081 12265 10084
rect 12299 10081 12311 10115
rect 16114 10112 16120 10124
rect 16075 10084 16120 10112
rect 12253 10075 12311 10081
rect 16114 10072 16120 10084
rect 16172 10072 16178 10124
rect 16758 10072 16764 10124
rect 16816 10112 16822 10124
rect 16945 10115 17003 10121
rect 16945 10112 16957 10115
rect 16816 10084 16957 10112
rect 16816 10072 16822 10084
rect 16945 10081 16957 10084
rect 16991 10081 17003 10115
rect 16945 10075 17003 10081
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2314 10044 2320 10056
rect 2275 10016 2320 10044
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 3050 10044 3056 10056
rect 3011 10016 3056 10044
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4338 10044 4344 10056
rect 4203 10016 4344 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4522 10044 4528 10056
rect 4483 10016 4528 10044
rect 4522 10004 4528 10016
rect 4580 10044 4586 10056
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 4580 10016 5457 10044
rect 4580 10004 4586 10016
rect 5445 10013 5457 10016
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5592 10016 6009 10044
rect 5592 10004 5598 10016
rect 5997 10013 6009 10016
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10044 6331 10047
rect 7650 10044 7656 10056
rect 6319 10016 7656 10044
rect 6319 10013 6331 10016
rect 6273 10007 6331 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 8110 10044 8116 10056
rect 8071 10016 8116 10044
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 10249 10047 10307 10053
rect 10249 10013 10261 10047
rect 10295 10044 10307 10047
rect 10410 10044 10416 10056
rect 10295 10016 10416 10044
rect 10295 10013 10307 10016
rect 10249 10007 10307 10013
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 11330 10044 11336 10056
rect 11291 10016 11336 10044
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11514 10044 11520 10056
rect 11475 10016 11520 10044
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 11793 10047 11851 10053
rect 11793 10044 11805 10047
rect 11756 10016 11805 10044
rect 11756 10004 11762 10016
rect 11793 10013 11805 10016
rect 11839 10013 11851 10047
rect 11793 10007 11851 10013
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12032 10016 13584 10044
rect 12032 10004 12038 10016
rect 2866 9936 2872 9988
rect 2924 9976 2930 9988
rect 3145 9979 3203 9985
rect 3145 9976 3157 9979
rect 2924 9948 3157 9976
rect 2924 9936 2930 9948
rect 3145 9945 3157 9948
rect 3191 9945 3203 9979
rect 4356 9976 4384 10004
rect 4614 9976 4620 9988
rect 4356 9948 4620 9976
rect 3145 9939 3203 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 6540 9979 6598 9985
rect 6540 9945 6552 9979
rect 6586 9976 6598 9979
rect 6730 9976 6736 9988
rect 6586 9948 6736 9976
rect 6586 9945 6598 9948
rect 6540 9939 6598 9945
rect 6730 9936 6736 9948
rect 6788 9936 6794 9988
rect 8573 9979 8631 9985
rect 8573 9945 8585 9979
rect 8619 9976 8631 9979
rect 9306 9976 9312 9988
rect 8619 9948 9312 9976
rect 8619 9945 8631 9948
rect 8573 9939 8631 9945
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 10778 9936 10784 9988
rect 10836 9976 10842 9988
rect 10965 9979 11023 9985
rect 10965 9976 10977 9979
rect 10836 9948 10977 9976
rect 10836 9936 10842 9948
rect 10965 9945 10977 9948
rect 11011 9945 11023 9979
rect 10965 9939 11023 9945
rect 12342 9936 12348 9988
rect 12400 9976 12406 9988
rect 12498 9979 12556 9985
rect 12498 9976 12510 9979
rect 12400 9948 12510 9976
rect 12400 9936 12406 9948
rect 12498 9945 12510 9948
rect 12544 9945 12556 9979
rect 12498 9939 12556 9945
rect 4706 9908 4712 9920
rect 4667 9880 4712 9908
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 5776 9880 5825 9908
rect 5776 9868 5782 9880
rect 5813 9877 5825 9880
rect 5859 9877 5871 9911
rect 5813 9871 5871 9877
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 7653 9911 7711 9917
rect 7653 9908 7665 9911
rect 7616 9880 7665 9908
rect 7616 9868 7622 9880
rect 7653 9877 7665 9880
rect 7699 9877 7711 9911
rect 7653 9871 7711 9877
rect 9125 9911 9183 9917
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9674 9908 9680 9920
rect 9171 9880 9680 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9674 9868 9680 9880
rect 9732 9908 9738 9920
rect 10686 9908 10692 9920
rect 9732 9880 10692 9908
rect 9732 9868 9738 9880
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 10870 9908 10876 9920
rect 10831 9880 10876 9908
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11977 9911 12035 9917
rect 11977 9877 11989 9911
rect 12023 9908 12035 9911
rect 12618 9908 12624 9920
rect 12023 9880 12624 9908
rect 12023 9877 12035 9880
rect 11977 9871 12035 9877
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 13556 9908 13584 10016
rect 14274 10004 14280 10056
rect 14332 10044 14338 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 14332 10016 15485 10044
rect 14332 10004 14338 10016
rect 15473 10013 15485 10016
rect 15519 10013 15531 10047
rect 15473 10007 15531 10013
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10044 16359 10047
rect 17770 10044 17776 10056
rect 16347 10016 17776 10044
rect 16347 10013 16359 10016
rect 16301 10007 16359 10013
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 13814 9936 13820 9988
rect 13872 9976 13878 9988
rect 15206 9979 15264 9985
rect 15206 9976 15218 9979
rect 13872 9948 15218 9976
rect 13872 9936 13878 9948
rect 15206 9945 15218 9948
rect 15252 9945 15264 9979
rect 15206 9939 15264 9945
rect 17212 9979 17270 9985
rect 17212 9945 17224 9979
rect 17258 9976 17270 9979
rect 17310 9976 17316 9988
rect 17258 9948 17316 9976
rect 17258 9945 17270 9948
rect 17212 9939 17270 9945
rect 17310 9936 17316 9948
rect 17368 9936 17374 9988
rect 13633 9911 13691 9917
rect 13633 9908 13645 9911
rect 13556 9880 13645 9908
rect 13633 9877 13645 9880
rect 13679 9908 13691 9911
rect 13906 9908 13912 9920
rect 13679 9880 13912 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 14090 9908 14096 9920
rect 14003 9880 14096 9908
rect 14090 9868 14096 9880
rect 14148 9908 14154 9920
rect 14458 9908 14464 9920
rect 14148 9880 14464 9908
rect 14148 9868 14154 9880
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 15286 9868 15292 9920
rect 15344 9908 15350 9920
rect 15654 9908 15660 9920
rect 15344 9880 15660 9908
rect 15344 9868 15350 9880
rect 15654 9868 15660 9880
rect 15712 9908 15718 9920
rect 16206 9908 16212 9920
rect 15712 9880 16212 9908
rect 15712 9868 15718 9880
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 16669 9911 16727 9917
rect 16669 9877 16681 9911
rect 16715 9908 16727 9911
rect 16850 9908 16856 9920
rect 16715 9880 16856 9908
rect 16715 9877 16727 9880
rect 16669 9871 16727 9877
rect 16850 9868 16856 9880
rect 16908 9868 16914 9920
rect 1104 9818 18860 9840
rect 1104 9766 6880 9818
rect 6932 9766 6944 9818
rect 6996 9766 7008 9818
rect 7060 9766 7072 9818
rect 7124 9766 7136 9818
rect 7188 9766 12811 9818
rect 12863 9766 12875 9818
rect 12927 9766 12939 9818
rect 12991 9766 13003 9818
rect 13055 9766 13067 9818
rect 13119 9766 18860 9818
rect 1104 9744 18860 9766
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6788 9676 6837 9704
rect 6788 9664 6794 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 7558 9704 7564 9716
rect 6825 9667 6883 9673
rect 7208 9676 7564 9704
rect 4341 9639 4399 9645
rect 4341 9605 4353 9639
rect 4387 9636 4399 9639
rect 5534 9636 5540 9648
rect 4387 9608 5540 9636
rect 4387 9605 4399 9608
rect 4341 9599 4399 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 7208 9636 7236 9676
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 9674 9704 9680 9716
rect 8168 9676 9680 9704
rect 8168 9664 8174 9676
rect 9674 9664 9680 9676
rect 9732 9704 9738 9716
rect 10778 9704 10784 9716
rect 9732 9676 10784 9704
rect 9732 9664 9738 9676
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 10870 9664 10876 9716
rect 10928 9704 10934 9716
rect 13630 9704 13636 9716
rect 10928 9676 13636 9704
rect 10928 9664 10934 9676
rect 13630 9664 13636 9676
rect 13688 9704 13694 9716
rect 13688 9676 13860 9704
rect 13688 9664 13694 9676
rect 7742 9636 7748 9648
rect 7116 9608 7236 9636
rect 7392 9608 7748 9636
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2314 9568 2320 9580
rect 2275 9540 2320 9568
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2547 9540 2973 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2961 9537 2973 9540
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4246 9568 4252 9580
rect 4203 9540 4252 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 5718 9528 5724 9580
rect 5776 9577 5782 9580
rect 5776 9568 5788 9577
rect 5994 9568 6000 9580
rect 5776 9540 5821 9568
rect 5955 9540 6000 9568
rect 5776 9531 5788 9540
rect 5776 9528 5782 9531
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 7116 9577 7144 9608
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9537 7159 9571
rect 7282 9568 7288 9580
rect 7243 9540 7288 9568
rect 7101 9531 7159 9537
rect 3973 9503 4031 9509
rect 3973 9469 3985 9503
rect 4019 9500 4031 9503
rect 4706 9500 4712 9512
rect 4019 9472 4712 9500
rect 4019 9469 4031 9472
rect 3973 9463 4031 9469
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 7024 9500 7052 9531
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 7392 9577 7420 9608
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 10796 9646 10833 9664
rect 10805 9636 10833 9646
rect 12526 9636 12532 9648
rect 10805 9608 12532 9636
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 12618 9596 12624 9648
rect 12676 9645 12682 9648
rect 12676 9636 12688 9645
rect 12676 9608 12721 9636
rect 12676 9599 12688 9608
rect 12676 9596 12682 9599
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7650 9568 7656 9580
rect 7611 9540 7656 9568
rect 7377 9531 7435 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7926 9577 7932 9580
rect 7920 9568 7932 9577
rect 7887 9540 7932 9568
rect 7920 9531 7932 9540
rect 7926 9528 7932 9531
rect 7984 9528 7990 9580
rect 9306 9568 9312 9580
rect 9267 9540 9312 9568
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 13832 9577 13860 9676
rect 14550 9664 14556 9716
rect 14608 9704 14614 9716
rect 14645 9707 14703 9713
rect 14645 9704 14657 9707
rect 14608 9676 14657 9704
rect 14608 9664 14614 9676
rect 14645 9673 14657 9676
rect 14691 9673 14703 9707
rect 14645 9667 14703 9673
rect 14918 9664 14924 9716
rect 14976 9664 14982 9716
rect 17310 9704 17316 9716
rect 15396 9676 15792 9704
rect 17271 9676 17316 9704
rect 14936 9636 14964 9664
rect 15396 9636 15424 9676
rect 14936 9608 15424 9636
rect 15764 9636 15792 9676
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 16758 9636 16764 9648
rect 15764 9608 16764 9636
rect 13173 9571 13231 9577
rect 13173 9537 13185 9571
rect 13219 9568 13231 9571
rect 13633 9571 13691 9577
rect 13633 9568 13645 9571
rect 13219 9540 13645 9568
rect 13219 9537 13231 9540
rect 13173 9531 13231 9537
rect 13633 9537 13645 9540
rect 13679 9537 13691 9571
rect 13633 9531 13691 9537
rect 13817 9571 13875 9577
rect 13817 9537 13829 9571
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 14090 9568 14096 9580
rect 14047 9540 14096 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 14182 9528 14188 9580
rect 14240 9568 14246 9580
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 14240 9540 14289 9568
rect 14240 9528 14246 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9568 14887 9571
rect 14936 9568 14964 9608
rect 16758 9596 16764 9608
rect 16816 9636 16822 9648
rect 16816 9608 17448 9636
rect 16816 9596 16822 9608
rect 17420 9580 17448 9608
rect 17586 9596 17592 9648
rect 17644 9636 17650 9648
rect 18230 9636 18236 9648
rect 17644 9608 18236 9636
rect 17644 9596 17650 9608
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 14875 9540 14964 9568
rect 14875 9537 14887 9540
rect 14829 9531 14887 9537
rect 15562 9528 15568 9580
rect 15620 9568 15626 9580
rect 15620 9540 15665 9568
rect 15620 9528 15626 9540
rect 15746 9528 15752 9580
rect 15804 9568 15810 9580
rect 16117 9571 16175 9577
rect 15804 9540 15849 9568
rect 15804 9528 15810 9540
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16163 9540 16681 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16850 9568 16856 9580
rect 16811 9540 16856 9568
rect 16669 9531 16727 9537
rect 16850 9528 16856 9540
rect 16908 9528 16914 9580
rect 17402 9528 17408 9580
rect 17460 9568 17466 9580
rect 17497 9571 17555 9577
rect 17497 9568 17509 9571
rect 17460 9540 17509 9568
rect 17460 9528 17466 9540
rect 17497 9537 17509 9540
rect 17543 9537 17555 9571
rect 17497 9531 17555 9537
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18049 9571 18107 9577
rect 18049 9568 18061 9571
rect 18012 9540 18061 9568
rect 18012 9528 18018 9540
rect 18049 9537 18061 9540
rect 18095 9537 18107 9571
rect 18049 9531 18107 9537
rect 7466 9500 7472 9512
rect 7024 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 14918 9500 14924 9512
rect 12943 9472 14924 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 15105 9503 15163 9509
rect 15105 9469 15117 9503
rect 15151 9500 15163 9503
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 15151 9472 15393 9500
rect 15151 9469 15163 9472
rect 15105 9463 15163 9469
rect 15381 9469 15393 9472
rect 15427 9469 15439 9503
rect 17034 9500 17040 9512
rect 16995 9472 17040 9500
rect 15381 9463 15439 9469
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 17770 9500 17776 9512
rect 17731 9472 17776 9500
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 13357 9435 13415 9441
rect 13357 9401 13369 9435
rect 13403 9432 13415 9435
rect 13814 9432 13820 9444
rect 13403 9404 13820 9432
rect 13403 9401 13415 9404
rect 13357 9395 13415 9401
rect 13814 9392 13820 9404
rect 13872 9392 13878 9444
rect 16301 9435 16359 9441
rect 16301 9401 16313 9435
rect 16347 9432 16359 9435
rect 16942 9432 16948 9444
rect 16347 9404 16948 9432
rect 16347 9401 16359 9404
rect 16301 9395 16359 9401
rect 16942 9392 16948 9404
rect 17000 9392 17006 9444
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 2832 9336 2877 9364
rect 2832 9324 2838 9336
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 4617 9367 4675 9373
rect 4617 9364 4629 9367
rect 4488 9336 4629 9364
rect 4488 9324 4494 9336
rect 4617 9333 4629 9336
rect 4663 9333 4675 9367
rect 4617 9327 4675 9333
rect 9033 9367 9091 9373
rect 9033 9333 9045 9367
rect 9079 9364 9091 9367
rect 10410 9364 10416 9376
rect 9079 9336 10416 9364
rect 9079 9333 9091 9336
rect 9033 9327 9091 9333
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 10594 9364 10600 9376
rect 10555 9336 10600 9364
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 11388 9336 11529 9364
rect 11388 9324 11394 9336
rect 11517 9333 11529 9336
rect 11563 9364 11575 9367
rect 13078 9364 13084 9376
rect 11563 9336 13084 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 15010 9364 15016 9376
rect 14971 9336 15016 9364
rect 15010 9324 15016 9336
rect 15068 9324 15074 9376
rect 17678 9364 17684 9376
rect 17639 9336 17684 9364
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 1104 9274 18860 9296
rect 1104 9222 3915 9274
rect 3967 9222 3979 9274
rect 4031 9222 4043 9274
rect 4095 9222 4107 9274
rect 4159 9222 4171 9274
rect 4223 9222 9846 9274
rect 9898 9222 9910 9274
rect 9962 9222 9974 9274
rect 10026 9222 10038 9274
rect 10090 9222 10102 9274
rect 10154 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 15904 9274
rect 15956 9222 15968 9274
rect 16020 9222 16032 9274
rect 16084 9222 18860 9274
rect 1104 9200 18860 9222
rect 4065 9163 4123 9169
rect 4065 9129 4077 9163
rect 4111 9160 4123 9163
rect 4246 9160 4252 9172
rect 4111 9132 4252 9160
rect 4111 9129 4123 9132
rect 4065 9123 4123 9129
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 7834 9120 7840 9172
rect 7892 9160 7898 9172
rect 7929 9163 7987 9169
rect 7929 9160 7941 9163
rect 7892 9132 7941 9160
rect 7892 9120 7898 9132
rect 7929 9129 7941 9132
rect 7975 9129 7987 9163
rect 9122 9160 9128 9172
rect 9083 9132 9128 9160
rect 7929 9123 7987 9129
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 9953 9163 10011 9169
rect 9953 9129 9965 9163
rect 9999 9160 10011 9163
rect 10226 9160 10232 9172
rect 9999 9132 10232 9160
rect 9999 9129 10011 9132
rect 9953 9123 10011 9129
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 10410 9120 10416 9172
rect 10468 9160 10474 9172
rect 10965 9163 11023 9169
rect 10965 9160 10977 9163
rect 10468 9132 10977 9160
rect 10468 9120 10474 9132
rect 10965 9129 10977 9132
rect 11011 9160 11023 9163
rect 11146 9160 11152 9172
rect 11011 9132 11152 9160
rect 11011 9129 11023 9132
rect 10965 9123 11023 9129
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 11514 9160 11520 9172
rect 11475 9132 11520 9160
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 12253 9163 12311 9169
rect 11848 9132 12204 9160
rect 11848 9120 11854 9132
rect 12176 9104 12204 9132
rect 12253 9129 12265 9163
rect 12299 9160 12311 9163
rect 12342 9160 12348 9172
rect 12299 9132 12348 9160
rect 12299 9129 12311 9132
rect 12253 9123 12311 9129
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 14090 9160 14096 9172
rect 14051 9132 14096 9160
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 14182 9120 14188 9172
rect 14240 9160 14246 9172
rect 15841 9163 15899 9169
rect 15841 9160 15853 9163
rect 14240 9132 15853 9160
rect 14240 9120 14246 9132
rect 15841 9129 15853 9132
rect 15887 9129 15899 9163
rect 17770 9160 17776 9172
rect 17731 9132 17776 9160
rect 15841 9123 15899 9129
rect 6546 9092 6552 9104
rect 6507 9064 6552 9092
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 11974 9092 11980 9104
rect 11072 9064 11980 9092
rect 4706 9024 4712 9036
rect 4619 8996 4712 9024
rect 4706 8984 4712 8996
rect 4764 9024 4770 9036
rect 5077 9027 5135 9033
rect 5077 9024 5089 9027
rect 4764 8996 5089 9024
rect 4764 8984 4770 8996
rect 5077 8993 5089 8996
rect 5123 8993 5135 9027
rect 10594 9024 10600 9036
rect 5077 8987 5135 8993
rect 6748 8996 10600 9024
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 1848 8959 1906 8965
rect 1848 8925 1860 8959
rect 1894 8956 1906 8959
rect 2774 8956 2780 8968
rect 1894 8928 2780 8956
rect 1894 8925 1906 8928
rect 1848 8919 1906 8925
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 5442 8956 5448 8968
rect 3283 8928 5448 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 6086 8956 6092 8968
rect 6047 8928 6092 8956
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6748 8965 6776 8996
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 11072 9033 11100 9064
rect 11974 9052 11980 9064
rect 12032 9052 12038 9104
rect 12158 9052 12164 9104
rect 12216 9092 12222 9104
rect 12216 9064 14780 9092
rect 12216 9052 12222 9064
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 8993 11115 9027
rect 11057 8987 11115 8993
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 11655 9027 11713 9033
rect 11296 8996 11468 9024
rect 11296 8984 11302 8996
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8925 6791 8959
rect 7558 8956 7564 8968
rect 7471 8928 7564 8956
rect 6733 8919 6791 8925
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 8110 8956 8116 8968
rect 8071 8928 8116 8956
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 8260 8928 8309 8956
rect 8260 8916 8266 8928
rect 8297 8925 8309 8928
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 8754 8956 8760 8968
rect 8435 8928 8760 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 2866 8848 2872 8900
rect 2924 8888 2930 8900
rect 4525 8891 4583 8897
rect 4525 8888 4537 8891
rect 2924 8860 4537 8888
rect 2924 8848 2930 8860
rect 4525 8857 4537 8860
rect 4571 8857 4583 8891
rect 5258 8888 5264 8900
rect 5219 8860 5264 8888
rect 4525 8851 4583 8857
rect 5258 8848 5264 8860
rect 5316 8848 5322 8900
rect 7576 8888 7604 8916
rect 8404 8888 8432 8919
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 9582 8956 9588 8968
rect 9543 8928 9588 8956
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 9732 8928 9781 8956
rect 9732 8916 9738 8928
rect 9769 8925 9781 8928
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 10962 8956 10968 8968
rect 10827 8928 10968 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11333 8959 11391 8965
rect 11333 8925 11345 8959
rect 11379 8925 11391 8959
rect 11440 8956 11468 8996
rect 11655 8993 11667 9027
rect 11701 9024 11713 9027
rect 12526 9024 12532 9036
rect 11701 8996 12532 9024
rect 11701 8993 11713 8996
rect 11655 8987 11713 8993
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 13078 9024 13084 9036
rect 12820 8996 13084 9024
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 11440 8928 11805 8956
rect 11333 8919 11391 8925
rect 11793 8925 11805 8928
rect 11839 8956 11851 8959
rect 11882 8956 11888 8968
rect 11839 8928 11888 8956
rect 11839 8925 11851 8928
rect 11793 8919 11851 8925
rect 7576 8860 8432 8888
rect 9309 8891 9367 8897
rect 9309 8857 9321 8891
rect 9355 8888 9367 8891
rect 9490 8888 9496 8900
rect 9355 8860 9496 8888
rect 9355 8857 9367 8860
rect 9309 8851 9367 8857
rect 9490 8848 9496 8860
rect 9548 8848 9554 8900
rect 11054 8888 11060 8900
rect 10428 8860 11060 8888
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 2961 8823 3019 8829
rect 2961 8820 2973 8823
rect 2832 8792 2973 8820
rect 2832 8780 2838 8792
rect 2961 8789 2973 8792
rect 3007 8789 3019 8823
rect 3418 8820 3424 8832
rect 3379 8792 3424 8820
rect 2961 8783 3019 8789
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 4430 8820 4436 8832
rect 4391 8792 4436 8820
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8820 6331 8823
rect 6454 8820 6460 8832
rect 6319 8792 6460 8820
rect 6319 8789 6331 8792
rect 6273 8783 6331 8789
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 7561 8823 7619 8829
rect 7561 8789 7573 8823
rect 7607 8820 7619 8823
rect 8386 8820 8392 8832
rect 7607 8792 8392 8820
rect 7607 8789 7619 8792
rect 7561 8783 7619 8789
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8536 8792 8953 8820
rect 8536 8780 8542 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 9109 8823 9167 8829
rect 9109 8789 9121 8823
rect 9155 8820 9167 8823
rect 10428 8820 10456 8860
rect 11054 8848 11060 8860
rect 11112 8848 11118 8900
rect 10594 8820 10600 8832
rect 9155 8792 10456 8820
rect 10555 8792 10600 8820
rect 9155 8789 9167 8792
rect 9109 8783 9167 8789
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 11348 8820 11376 8919
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 12069 8959 12127 8965
rect 12069 8925 12081 8959
rect 12115 8925 12127 8959
rect 12250 8956 12256 8968
rect 12211 8928 12256 8956
rect 12069 8919 12127 8925
rect 11425 8891 11483 8897
rect 11425 8857 11437 8891
rect 11471 8888 11483 8891
rect 11698 8888 11704 8900
rect 11471 8860 11704 8888
rect 11471 8857 11483 8860
rect 11425 8851 11483 8857
rect 11698 8848 11704 8860
rect 11756 8888 11762 8900
rect 12084 8888 12112 8919
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 12820 8965 12848 8996
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 14752 9033 14780 9064
rect 14737 9027 14795 9033
rect 14737 8993 14749 9027
rect 14783 9024 14795 9027
rect 15856 9024 15884 9123
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 16209 9027 16267 9033
rect 16209 9024 16221 9027
rect 14783 8996 15700 9024
rect 15856 8996 16221 9024
rect 14783 8993 14795 8996
rect 14737 8987 14795 8993
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8925 12863 8959
rect 12986 8956 12992 8968
rect 12947 8928 12992 8956
rect 12805 8919 12863 8925
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8956 13231 8959
rect 13446 8956 13452 8968
rect 13219 8928 13452 8956
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 15562 8956 15568 8968
rect 15523 8928 15568 8956
rect 15562 8916 15568 8928
rect 15620 8916 15626 8968
rect 15672 8956 15700 8996
rect 16209 8993 16221 8996
rect 16255 9024 16267 9027
rect 17034 9024 17040 9036
rect 16255 8996 17040 9024
rect 16255 8993 16267 8996
rect 16209 8987 16267 8993
rect 17034 8984 17040 8996
rect 17092 8984 17098 9036
rect 16114 8956 16120 8968
rect 15672 8928 16120 8956
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16390 8956 16396 8968
rect 16351 8928 16396 8956
rect 16390 8916 16396 8928
rect 16448 8916 16454 8968
rect 16577 8959 16635 8965
rect 16577 8925 16589 8959
rect 16623 8956 16635 8959
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16623 8928 16865 8956
rect 16623 8925 16635 8928
rect 16577 8919 16635 8925
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 17494 8956 17500 8968
rect 17455 8928 17500 8956
rect 16853 8919 16911 8925
rect 17494 8916 17500 8928
rect 17552 8916 17558 8968
rect 17954 8956 17960 8968
rect 17915 8928 17960 8956
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 18046 8916 18052 8968
rect 18104 8956 18110 8968
rect 18104 8928 18149 8956
rect 18104 8916 18110 8928
rect 11756 8860 12112 8888
rect 12176 8860 12434 8888
rect 11756 8848 11762 8860
rect 12176 8820 12204 8860
rect 11348 8792 12204 8820
rect 12406 8820 12434 8860
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 13081 8891 13139 8897
rect 13081 8888 13093 8891
rect 12768 8860 13093 8888
rect 12768 8848 12774 8860
rect 13081 8857 13093 8860
rect 13127 8857 13139 8891
rect 13725 8891 13783 8897
rect 13081 8851 13139 8857
rect 13188 8860 13676 8888
rect 13188 8820 13216 8860
rect 12406 8792 13216 8820
rect 13357 8823 13415 8829
rect 13357 8789 13369 8823
rect 13403 8820 13415 8823
rect 13538 8820 13544 8832
rect 13403 8792 13544 8820
rect 13403 8789 13415 8792
rect 13357 8783 13415 8789
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 13648 8820 13676 8860
rect 13725 8857 13737 8891
rect 13771 8888 13783 8891
rect 16482 8888 16488 8900
rect 13771 8860 16488 8888
rect 13771 8857 13783 8860
rect 13725 8851 13783 8857
rect 16482 8848 16488 8860
rect 16540 8848 16546 8900
rect 13998 8820 14004 8832
rect 13648 8792 14004 8820
rect 13998 8780 14004 8792
rect 14056 8780 14062 8832
rect 14182 8780 14188 8832
rect 14240 8820 14246 8832
rect 14461 8823 14519 8829
rect 14461 8820 14473 8823
rect 14240 8792 14473 8820
rect 14240 8780 14246 8792
rect 14461 8789 14473 8792
rect 14507 8789 14519 8823
rect 14461 8783 14519 8789
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 14608 8792 14653 8820
rect 14608 8780 14614 8792
rect 15194 8780 15200 8832
rect 15252 8820 15258 8832
rect 15381 8823 15439 8829
rect 15381 8820 15393 8823
rect 15252 8792 15393 8820
rect 15252 8780 15258 8792
rect 15381 8789 15393 8792
rect 15427 8789 15439 8823
rect 15381 8783 15439 8789
rect 15562 8780 15568 8832
rect 15620 8820 15626 8832
rect 16206 8820 16212 8832
rect 15620 8792 16212 8820
rect 15620 8780 15626 8792
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 17034 8820 17040 8832
rect 16995 8792 17040 8820
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 1104 8730 18860 8752
rect 1104 8678 6880 8730
rect 6932 8678 6944 8730
rect 6996 8678 7008 8730
rect 7060 8678 7072 8730
rect 7124 8678 7136 8730
rect 7188 8678 12811 8730
rect 12863 8678 12875 8730
rect 12927 8678 12939 8730
rect 12991 8678 13003 8730
rect 13055 8678 13067 8730
rect 13119 8678 18860 8730
rect 1104 8656 18860 8678
rect 1486 8616 1492 8628
rect 1447 8588 1492 8616
rect 1486 8576 1492 8588
rect 1544 8576 1550 8628
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2501 8619 2559 8625
rect 2501 8616 2513 8619
rect 2372 8588 2513 8616
rect 2372 8576 2378 8588
rect 2501 8585 2513 8588
rect 2547 8585 2559 8619
rect 2866 8616 2872 8628
rect 2827 8588 2872 8616
rect 2501 8579 2559 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 5166 8616 5172 8628
rect 5127 8588 5172 8616
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5442 8616 5448 8628
rect 5403 8588 5448 8616
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 7742 8616 7748 8628
rect 6288 8588 7748 8616
rect 3418 8508 3424 8560
rect 3476 8548 3482 8560
rect 4034 8551 4092 8557
rect 4034 8548 4046 8551
rect 3476 8520 4046 8548
rect 3476 8508 3482 8520
rect 4034 8517 4046 8520
rect 4080 8517 4092 8551
rect 4034 8511 4092 8517
rect 4798 8508 4804 8560
rect 4856 8548 4862 8560
rect 4856 8520 5764 8548
rect 4856 8508 4862 8520
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1719 8452 2053 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 5626 8480 5632 8492
rect 2179 8452 5488 8480
rect 5587 8452 5632 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2832 8384 2973 8412
rect 2832 8372 2838 8384
rect 2961 8381 2973 8384
rect 3007 8381 3019 8415
rect 3142 8412 3148 8424
rect 3103 8384 3148 8412
rect 2961 8375 3019 8381
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8381 3847 8415
rect 5460 8412 5488 8452
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5736 8489 5764 8520
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 6288 8412 6316 8588
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 8849 8619 8907 8625
rect 8849 8616 8861 8619
rect 8168 8588 8861 8616
rect 8168 8576 8174 8588
rect 8849 8585 8861 8588
rect 8895 8585 8907 8619
rect 10870 8616 10876 8628
rect 8849 8579 8907 8585
rect 9048 8588 10876 8616
rect 7282 8548 7288 8560
rect 6380 8520 7288 8548
rect 6380 8489 6408 8520
rect 7282 8508 7288 8520
rect 7340 8508 7346 8560
rect 8386 8548 8392 8560
rect 8347 8520 8392 8548
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 6621 8483 6679 8489
rect 6621 8480 6633 8483
rect 6512 8452 6633 8480
rect 6512 8440 6518 8452
rect 6621 8449 6633 8452
rect 6667 8449 6679 8483
rect 6621 8443 6679 8449
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 8202 8480 8208 8492
rect 7524 8452 8208 8480
rect 7524 8440 7530 8452
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 9048 8489 9076 8588
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11609 8619 11667 8625
rect 11609 8585 11621 8619
rect 11655 8616 11667 8619
rect 11698 8616 11704 8628
rect 11655 8588 11704 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 12618 8616 12624 8628
rect 11808 8588 12624 8616
rect 10226 8508 10232 8560
rect 10284 8548 10290 8560
rect 10502 8548 10508 8560
rect 10284 8520 10508 8548
rect 10284 8508 10290 8520
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 10594 8508 10600 8560
rect 10652 8548 10658 8560
rect 10790 8551 10848 8557
rect 10790 8548 10802 8551
rect 10652 8520 10802 8548
rect 10652 8508 10658 8520
rect 10790 8517 10802 8520
rect 10836 8517 10848 8551
rect 10790 8511 10848 8517
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 11808 8489 11836 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 14090 8616 14096 8628
rect 13096 8588 14096 8616
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 9180 8452 9225 8480
rect 10060 8452 11805 8480
rect 9180 8440 9186 8452
rect 5460 8384 6316 8412
rect 9217 8415 9275 8421
rect 3789 8375 3847 8381
rect 9217 8381 9229 8415
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8412 9367 8415
rect 9674 8412 9680 8424
rect 9355 8384 9680 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 1578 8304 1584 8356
rect 1636 8344 1642 8356
rect 3804 8344 3832 8375
rect 8573 8347 8631 8353
rect 1636 8316 3832 8344
rect 5092 8316 5304 8344
rect 1636 8304 1642 8316
rect 2222 8236 2228 8288
rect 2280 8276 2286 8288
rect 5092 8276 5120 8316
rect 2280 8248 5120 8276
rect 5276 8276 5304 8316
rect 8573 8313 8585 8347
rect 8619 8344 8631 8347
rect 9232 8344 9260 8375
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 9490 8344 9496 8356
rect 8619 8316 9076 8344
rect 9232 8316 9496 8344
rect 8619 8313 8631 8316
rect 8573 8307 8631 8313
rect 7374 8276 7380 8288
rect 5276 8248 7380 8276
rect 2280 8236 2286 8248
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 9048 8276 9076 8316
rect 9490 8304 9496 8316
rect 9548 8304 9554 8356
rect 10060 8344 10088 8452
rect 11793 8449 11805 8452
rect 11839 8449 11851 8483
rect 12066 8480 12072 8492
rect 12027 8452 12072 8480
rect 11793 8443 11851 8449
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 12250 8489 12256 8492
rect 12248 8480 12256 8489
rect 12211 8452 12256 8480
rect 12248 8443 12256 8452
rect 12250 8440 12256 8443
rect 12308 8440 12314 8492
rect 12348 8486 12406 8492
rect 12348 8452 12360 8486
rect 12394 8452 12406 8486
rect 12348 8446 12406 8452
rect 12483 8483 12541 8489
rect 12483 8449 12495 8483
rect 12529 8480 12541 8483
rect 12710 8480 12716 8492
rect 12529 8452 12716 8480
rect 12529 8449 12541 8452
rect 11057 8415 11115 8421
rect 11057 8381 11069 8415
rect 11103 8381 11115 8415
rect 12360 8412 12388 8446
rect 12483 8443 12541 8449
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12986 8480 12992 8492
rect 12947 8452 12992 8480
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13096 8480 13124 8588
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 17678 8616 17684 8628
rect 14844 8588 17684 8616
rect 13538 8508 13544 8560
rect 13596 8548 13602 8560
rect 14844 8548 14872 8588
rect 17678 8576 17684 8588
rect 17736 8576 17742 8628
rect 17034 8557 17040 8560
rect 17028 8548 17040 8557
rect 13596 8520 14136 8548
rect 13596 8508 13602 8520
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 13096 8452 13185 8480
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 13280 8412 13308 8443
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 13909 8483 13967 8489
rect 13412 8452 13457 8480
rect 13412 8440 13418 8452
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 13998 8480 14004 8492
rect 13955 8452 14004 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 14108 8489 14136 8520
rect 14752 8520 14872 8548
rect 14936 8520 16804 8548
rect 16995 8520 17040 8548
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8449 14151 8483
rect 14274 8480 14280 8492
rect 14235 8452 14280 8480
rect 14093 8443 14151 8449
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 14458 8480 14464 8492
rect 14419 8452 14464 8480
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 14752 8480 14780 8520
rect 14936 8492 14964 8520
rect 16776 8492 16804 8520
rect 17028 8511 17040 8520
rect 17034 8508 17040 8511
rect 17092 8508 17098 8560
rect 14918 8480 14924 8492
rect 14568 8452 14780 8480
rect 14879 8452 14924 8480
rect 12360 8384 13308 8412
rect 11057 8375 11115 8381
rect 9600 8316 10088 8344
rect 9600 8276 9628 8316
rect 9048 8248 9628 8276
rect 9677 8279 9735 8285
rect 9677 8245 9689 8279
rect 9723 8276 9735 8279
rect 10410 8276 10416 8288
rect 9723 8248 10416 8276
rect 9723 8245 9735 8248
rect 9677 8239 9735 8245
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 11072 8276 11100 8375
rect 12544 8356 12572 8384
rect 12526 8304 12532 8356
rect 12584 8304 12590 8356
rect 12713 8347 12771 8353
rect 12713 8313 12725 8347
rect 12759 8344 12771 8347
rect 13280 8344 13308 8384
rect 13814 8372 13820 8424
rect 13872 8412 13878 8424
rect 14185 8415 14243 8421
rect 14185 8412 14197 8415
rect 13872 8384 14197 8412
rect 13872 8372 13878 8384
rect 14185 8381 14197 8384
rect 14231 8381 14243 8415
rect 14185 8375 14243 8381
rect 13354 8344 13360 8356
rect 12759 8316 13032 8344
rect 13280 8316 13360 8344
rect 12759 8313 12771 8316
rect 12713 8307 12771 8313
rect 12158 8276 12164 8288
rect 11072 8248 12164 8276
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 13004 8276 13032 8316
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 13633 8347 13691 8353
rect 13633 8313 13645 8347
rect 13679 8344 13691 8347
rect 14568 8344 14596 8452
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 15177 8483 15235 8489
rect 15177 8480 15189 8483
rect 15028 8452 15189 8480
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8412 14703 8415
rect 15028 8412 15056 8452
rect 15177 8449 15189 8452
rect 15223 8449 15235 8483
rect 16758 8480 16764 8492
rect 16671 8452 16764 8480
rect 15177 8443 15235 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 14691 8384 15056 8412
rect 14691 8381 14703 8384
rect 14645 8375 14703 8381
rect 13679 8316 14596 8344
rect 13679 8313 13691 8316
rect 13633 8307 13691 8313
rect 13538 8276 13544 8288
rect 13004 8248 13544 8276
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 16301 8279 16359 8285
rect 16301 8276 16313 8279
rect 14516 8248 16313 8276
rect 14516 8236 14522 8248
rect 16301 8245 16313 8248
rect 16347 8276 16359 8279
rect 17494 8276 17500 8288
rect 16347 8248 17500 8276
rect 16347 8245 16359 8248
rect 16301 8239 16359 8245
rect 17494 8236 17500 8248
rect 17552 8236 17558 8288
rect 18138 8276 18144 8288
rect 18099 8248 18144 8276
rect 18138 8236 18144 8248
rect 18196 8236 18202 8288
rect 1104 8186 18860 8208
rect 1104 8134 3915 8186
rect 3967 8134 3979 8186
rect 4031 8134 4043 8186
rect 4095 8134 4107 8186
rect 4159 8134 4171 8186
rect 4223 8134 9846 8186
rect 9898 8134 9910 8186
rect 9962 8134 9974 8186
rect 10026 8134 10038 8186
rect 10090 8134 10102 8186
rect 10154 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 15904 8186
rect 15956 8134 15968 8186
rect 16020 8134 16032 8186
rect 16084 8134 18860 8186
rect 1104 8112 18860 8134
rect 4617 8075 4675 8081
rect 4617 8041 4629 8075
rect 4663 8072 4675 8075
rect 5626 8072 5632 8084
rect 4663 8044 5632 8072
rect 4663 8041 4675 8044
rect 4617 8035 4675 8041
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6457 8075 6515 8081
rect 6457 8072 6469 8075
rect 6144 8044 6469 8072
rect 6144 8032 6150 8044
rect 6457 8041 6469 8044
rect 6503 8041 6515 8075
rect 6457 8035 6515 8041
rect 11793 8075 11851 8081
rect 11793 8041 11805 8075
rect 11839 8072 11851 8075
rect 11839 8044 12204 8072
rect 11839 8041 11851 8044
rect 11793 8035 11851 8041
rect 7377 8007 7435 8013
rect 7377 7973 7389 8007
rect 7423 7973 7435 8007
rect 7377 7967 7435 7973
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7936 3111 7939
rect 3142 7936 3148 7948
rect 3099 7908 3148 7936
rect 3099 7905 3111 7908
rect 3053 7899 3111 7905
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4338 7936 4344 7948
rect 4111 7908 4344 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4338 7896 4344 7908
rect 4396 7936 4402 7948
rect 4706 7936 4712 7948
rect 4396 7908 4712 7936
rect 4396 7896 4402 7908
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 5902 7896 5908 7948
rect 5960 7896 5966 7948
rect 7392 7936 7420 7967
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 7800 7976 12112 8004
rect 7800 7964 7806 7976
rect 7834 7936 7840 7948
rect 6656 7908 7420 7936
rect 7795 7908 7840 7936
rect 2038 7828 2044 7880
rect 2096 7868 2102 7880
rect 2133 7871 2191 7877
rect 2133 7868 2145 7871
rect 2096 7840 2145 7868
rect 2096 7828 2102 7840
rect 2133 7837 2145 7840
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 4157 7871 4215 7877
rect 4157 7868 4169 7871
rect 2832 7840 4169 7868
rect 2832 7828 2838 7840
rect 4157 7837 4169 7840
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 5166 7868 5172 7880
rect 4295 7840 5172 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 5920 7868 5948 7896
rect 6089 7871 6147 7877
rect 5920 7840 6040 7868
rect 5534 7760 5540 7812
rect 5592 7800 5598 7812
rect 5905 7803 5963 7809
rect 5905 7800 5917 7803
rect 5592 7772 5917 7800
rect 5592 7760 5598 7772
rect 5905 7769 5917 7772
rect 5951 7769 5963 7803
rect 6012 7800 6040 7840
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6546 7868 6552 7880
rect 6135 7840 6552 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 6656 7877 6684 7908
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 8021 7939 8079 7945
rect 8021 7905 8033 7939
rect 8067 7936 8079 7939
rect 8478 7936 8484 7948
rect 8067 7908 8484 7936
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 9180 7908 9229 7936
rect 9180 7896 9186 7908
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 11054 7896 11060 7948
rect 11112 7936 11118 7948
rect 11112 7908 11376 7936
rect 11112 7896 11118 7908
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6748 7800 6776 7831
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 7432 7840 8953 7868
rect 7432 7828 7438 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 10410 7868 10416 7880
rect 10371 7840 10416 7868
rect 8941 7831 8999 7837
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 10686 7868 10692 7880
rect 10647 7840 10692 7868
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 7742 7800 7748 7812
rect 6012 7772 6776 7800
rect 7703 7772 7748 7800
rect 5905 7763 5963 7769
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 10502 7760 10508 7812
rect 10560 7800 10566 7812
rect 10597 7803 10655 7809
rect 10597 7800 10609 7803
rect 10560 7772 10609 7800
rect 10560 7760 10566 7772
rect 10597 7769 10609 7772
rect 10643 7769 10655 7803
rect 10597 7763 10655 7769
rect 10796 7800 10824 7831
rect 10870 7828 10876 7880
rect 10928 7868 10934 7880
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 10928 7840 11253 7868
rect 10928 7828 10934 7840
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11348 7868 11376 7908
rect 12084 7877 12112 7976
rect 12176 7936 12204 8044
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 13173 8075 13231 8081
rect 13173 8072 13185 8075
rect 12400 8044 13185 8072
rect 12400 8032 12406 8044
rect 13173 8041 13185 8044
rect 13219 8041 13231 8075
rect 14090 8072 14096 8084
rect 14051 8044 14096 8072
rect 13173 8035 13231 8041
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 14918 8032 14924 8084
rect 14976 8072 14982 8084
rect 15197 8075 15255 8081
rect 15197 8072 15209 8075
rect 14976 8044 15209 8072
rect 14976 8032 14982 8044
rect 15197 8041 15209 8044
rect 15243 8041 15255 8075
rect 15197 8035 15255 8041
rect 16301 8075 16359 8081
rect 16301 8041 16313 8075
rect 16347 8072 16359 8075
rect 16390 8072 16396 8084
rect 16347 8044 16396 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 14550 8004 14556 8016
rect 12912 7976 14556 8004
rect 12176 7908 12664 7936
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 11348 7840 11989 7868
rect 11241 7831 11299 7837
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7837 12219 7871
rect 12342 7868 12348 7880
rect 12303 7840 12348 7868
rect 12161 7831 12219 7837
rect 11514 7800 11520 7812
rect 10796 7772 11520 7800
rect 1946 7732 1952 7744
rect 1907 7704 1952 7732
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 2130 7692 2136 7744
rect 2188 7732 2194 7744
rect 2409 7735 2467 7741
rect 2409 7732 2421 7735
rect 2188 7704 2421 7732
rect 2188 7692 2194 7704
rect 2409 7701 2421 7704
rect 2455 7701 2467 7735
rect 2409 7695 2467 7701
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 3050 7732 3056 7744
rect 2915 7704 3056 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 3050 7692 3056 7704
rect 3108 7692 3114 7744
rect 8938 7692 8944 7744
rect 8996 7732 9002 7744
rect 10796 7732 10824 7772
rect 11514 7760 11520 7772
rect 11572 7760 11578 7812
rect 12176 7800 12204 7831
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 12636 7877 12664 7908
rect 12621 7871 12679 7877
rect 12621 7837 12633 7871
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 12710 7828 12716 7880
rect 12768 7868 12774 7880
rect 12912 7877 12940 7976
rect 14550 7964 14556 7976
rect 14608 7964 14614 8016
rect 16482 7964 16488 8016
rect 16540 8004 16546 8016
rect 16540 7976 17540 8004
rect 16540 7964 16546 7976
rect 13446 7936 13452 7948
rect 13004 7908 13452 7936
rect 13004 7877 13032 7908
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13725 7939 13783 7945
rect 13725 7905 13737 7939
rect 13771 7936 13783 7939
rect 14366 7936 14372 7948
rect 13771 7908 14372 7936
rect 13771 7905 13783 7908
rect 13725 7899 13783 7905
rect 14366 7896 14372 7908
rect 14424 7936 14430 7948
rect 14424 7908 15148 7936
rect 14424 7896 14430 7908
rect 12897 7871 12955 7877
rect 12768 7840 12813 7868
rect 12768 7828 12774 7840
rect 12897 7837 12909 7871
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13262 7828 13268 7880
rect 13320 7868 13326 7880
rect 14274 7877 14280 7880
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13320 7840 13553 7868
rect 13320 7828 13326 7840
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 14272 7868 14280 7877
rect 13541 7831 13599 7837
rect 13648 7840 14280 7868
rect 12250 7800 12256 7812
rect 12163 7772 12256 7800
rect 12250 7760 12256 7772
rect 12308 7800 12314 7812
rect 13648 7800 13676 7840
rect 14272 7831 14280 7840
rect 14274 7828 14280 7831
rect 14332 7828 14338 7880
rect 14458 7868 14464 7880
rect 14419 7840 14464 7868
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 14642 7868 14648 7880
rect 14603 7840 14648 7868
rect 14642 7828 14648 7840
rect 14700 7828 14706 7880
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7868 14795 7871
rect 14918 7868 14924 7880
rect 14783 7840 14924 7868
rect 14783 7837 14795 7840
rect 14737 7831 14795 7837
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 15120 7877 15148 7908
rect 16114 7896 16120 7948
rect 16172 7936 16178 7948
rect 17512 7945 17540 7976
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 16172 7908 16865 7936
rect 16172 7896 16178 7908
rect 16853 7905 16865 7908
rect 16899 7905 16911 7939
rect 16853 7899 16911 7905
rect 17497 7939 17555 7945
rect 17497 7905 17509 7939
rect 17543 7905 17555 7939
rect 17497 7899 17555 7905
rect 15105 7871 15163 7877
rect 15105 7837 15117 7871
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7868 16083 7871
rect 16298 7868 16304 7880
rect 16071 7840 16304 7868
rect 16071 7837 16083 7840
rect 16025 7831 16083 7837
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 16666 7868 16672 7880
rect 16579 7840 16672 7868
rect 16666 7828 16672 7840
rect 16724 7868 16730 7880
rect 17218 7868 17224 7880
rect 16724 7840 17224 7868
rect 16724 7828 16730 7840
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 17770 7868 17776 7880
rect 17731 7840 17776 7868
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 12308 7772 13676 7800
rect 14369 7803 14427 7809
rect 12308 7760 12314 7772
rect 14369 7769 14381 7803
rect 14415 7800 14427 7803
rect 14550 7800 14556 7812
rect 14415 7772 14556 7800
rect 14415 7769 14427 7772
rect 14369 7763 14427 7769
rect 14550 7760 14556 7772
rect 14608 7760 14614 7812
rect 14660 7800 14688 7828
rect 14660 7772 15884 7800
rect 10962 7732 10968 7744
rect 8996 7704 10824 7732
rect 10923 7704 10968 7732
rect 8996 7692 9002 7704
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11422 7732 11428 7744
rect 11383 7704 11428 7732
rect 11422 7692 11428 7704
rect 11480 7692 11486 7744
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 14918 7732 14924 7744
rect 12768 7704 14924 7732
rect 12768 7692 12774 7704
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 15856 7732 15884 7772
rect 16761 7735 16819 7741
rect 16761 7732 16773 7735
rect 15856 7704 16773 7732
rect 16761 7701 16773 7704
rect 16807 7732 16819 7735
rect 18138 7732 18144 7744
rect 16807 7704 18144 7732
rect 16807 7701 16819 7704
rect 16761 7695 16819 7701
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 1104 7642 18860 7664
rect 1104 7590 6880 7642
rect 6932 7590 6944 7642
rect 6996 7590 7008 7642
rect 7060 7590 7072 7642
rect 7124 7590 7136 7642
rect 7188 7590 12811 7642
rect 12863 7590 12875 7642
rect 12927 7590 12939 7642
rect 12991 7590 13003 7642
rect 13055 7590 13067 7642
rect 13119 7590 18860 7642
rect 1104 7568 18860 7590
rect 7466 7528 7472 7540
rect 7427 7500 7472 7528
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 9674 7528 9680 7540
rect 9635 7500 9680 7528
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 11146 7528 11152 7540
rect 9784 7500 11152 7528
rect 1946 7469 1952 7472
rect 1940 7460 1952 7469
rect 1907 7432 1952 7460
rect 1940 7423 1952 7432
rect 1946 7420 1952 7423
rect 2004 7420 2010 7472
rect 6638 7460 6644 7472
rect 4448 7432 6644 7460
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 4448 7401 4476 7432
rect 6638 7420 6644 7432
rect 6696 7460 6702 7472
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 6696 7432 6837 7460
rect 6696 7420 6702 7432
rect 6825 7429 6837 7432
rect 6871 7429 6883 7463
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 6825 7423 6883 7429
rect 7300 7432 7849 7460
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1636 7364 1685 7392
rect 1636 7352 1642 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4890 7392 4896 7404
rect 4851 7364 4896 7392
rect 4433 7355 4491 7361
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 5350 7392 5356 7404
rect 5311 7364 5356 7392
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 7300 7401 7328 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 7837 7423 7895 7429
rect 8053 7463 8111 7469
rect 8053 7429 8065 7463
rect 8099 7460 8111 7463
rect 8938 7460 8944 7472
rect 8099 7432 8944 7460
rect 8099 7429 8111 7432
rect 8053 7423 8111 7429
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 2682 7284 2688 7336
rect 2740 7324 2746 7336
rect 4157 7327 4215 7333
rect 4157 7324 4169 7327
rect 2740 7296 4169 7324
rect 2740 7284 2746 7296
rect 4157 7293 4169 7296
rect 4203 7293 4215 7327
rect 4157 7287 4215 7293
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 4798 7324 4804 7336
rect 4755 7296 4804 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 7300 7324 7328 7355
rect 7374 7352 7380 7404
rect 7432 7392 7438 7404
rect 7561 7395 7619 7401
rect 7432 7364 7512 7392
rect 7432 7352 7438 7364
rect 7300 7296 7420 7324
rect 7392 7268 7420 7296
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5902 7256 5908 7268
rect 5123 7228 5908 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 6638 7256 6644 7268
rect 6599 7228 6644 7256
rect 6638 7216 6644 7228
rect 6696 7216 6702 7268
rect 7374 7216 7380 7268
rect 7432 7216 7438 7268
rect 3050 7188 3056 7200
rect 3011 7160 3056 7188
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 5537 7191 5595 7197
rect 5537 7157 5549 7191
rect 5583 7188 5595 7191
rect 6270 7188 6276 7200
rect 5583 7160 6276 7188
rect 5583 7157 5595 7160
rect 5537 7151 5595 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 7484 7188 7512 7364
rect 7561 7361 7573 7395
rect 7607 7361 7619 7395
rect 7852 7392 7880 7423
rect 8938 7420 8944 7432
rect 8996 7420 9002 7472
rect 9784 7401 9812 7500
rect 11146 7488 11152 7500
rect 11204 7528 11210 7540
rect 14458 7528 14464 7540
rect 11204 7500 13492 7528
rect 11204 7488 11210 7500
rect 10318 7420 10324 7472
rect 10376 7460 10382 7472
rect 12618 7460 12624 7472
rect 10376 7432 10824 7460
rect 10376 7420 10382 7432
rect 10796 7401 10824 7432
rect 11072 7432 12624 7460
rect 8481 7395 8539 7401
rect 8481 7392 8493 7395
rect 7852 7364 8493 7392
rect 7561 7355 7619 7361
rect 8481 7361 8493 7364
rect 8527 7361 8539 7395
rect 9769 7395 9827 7401
rect 8481 7355 8539 7361
rect 8588 7364 9674 7392
rect 7576 7324 7604 7355
rect 8588 7336 8616 7364
rect 8570 7324 8576 7336
rect 7576 7296 8576 7324
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7324 8815 7327
rect 9490 7324 9496 7336
rect 8803 7296 9496 7324
rect 8803 7293 8815 7296
rect 8757 7287 8815 7293
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 9646 7324 9674 7364
rect 9769 7361 9781 7395
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 10689 7395 10747 7401
rect 10689 7361 10701 7395
rect 10735 7361 10747 7395
rect 10689 7355 10747 7361
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7361 10839 7395
rect 10962 7392 10968 7404
rect 10923 7364 10968 7392
rect 10781 7355 10839 7361
rect 10704 7324 10732 7355
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11072 7401 11100 7432
rect 12618 7420 12624 7432
rect 12676 7420 12682 7472
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7361 11115 7395
rect 11514 7392 11520 7404
rect 11475 7364 11520 7392
rect 11057 7355 11115 7361
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 12768 7364 12813 7392
rect 12768 7352 12774 7364
rect 11790 7324 11796 7336
rect 9646 7296 11008 7324
rect 11703 7296 11796 7324
rect 10980 7268 11008 7296
rect 11790 7284 11796 7296
rect 11848 7324 11854 7336
rect 12250 7324 12256 7336
rect 11848 7296 12256 7324
rect 11848 7284 11854 7296
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 12986 7324 12992 7336
rect 12400 7296 12992 7324
rect 12400 7284 12406 7296
rect 12986 7284 12992 7296
rect 13044 7324 13050 7336
rect 13464 7324 13492 7500
rect 13556 7500 14464 7528
rect 13556 7401 13584 7500
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 13633 7463 13691 7469
rect 13633 7429 13645 7463
rect 13679 7460 13691 7463
rect 14829 7463 14887 7469
rect 13679 7432 14044 7460
rect 13679 7429 13691 7432
rect 13633 7423 13691 7429
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7361 13599 7395
rect 13541 7355 13599 7361
rect 13648 7324 13676 7423
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7361 13783 7395
rect 13906 7392 13912 7404
rect 13867 7364 13912 7392
rect 13725 7355 13783 7361
rect 13044 7296 13400 7324
rect 13464 7296 13676 7324
rect 13740 7324 13768 7355
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 13740 7296 13860 7324
rect 13044 7284 13050 7296
rect 8205 7259 8263 7265
rect 8205 7225 8217 7259
rect 8251 7256 8263 7259
rect 9766 7256 9772 7268
rect 8251 7228 9772 7256
rect 8251 7225 8263 7228
rect 8205 7219 8263 7225
rect 9766 7216 9772 7228
rect 9824 7256 9830 7268
rect 10870 7256 10876 7268
rect 9824 7228 10876 7256
rect 9824 7216 9830 7228
rect 10870 7216 10876 7228
rect 10928 7216 10934 7268
rect 10962 7216 10968 7268
rect 11020 7216 11026 7268
rect 11146 7216 11152 7268
rect 11204 7256 11210 7268
rect 12710 7256 12716 7268
rect 11204 7228 12716 7256
rect 11204 7216 11210 7228
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 12894 7256 12900 7268
rect 12855 7228 12900 7256
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 13372 7256 13400 7296
rect 13372 7228 13676 7256
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7484 7160 8033 7188
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 10505 7191 10563 7197
rect 10505 7157 10517 7191
rect 10551 7188 10563 7191
rect 10594 7188 10600 7200
rect 10551 7160 10600 7188
rect 10551 7157 10563 7160
rect 10505 7151 10563 7157
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12912 7188 12940 7216
rect 12676 7160 12940 7188
rect 12676 7148 12682 7160
rect 13262 7148 13268 7200
rect 13320 7188 13326 7200
rect 13357 7191 13415 7197
rect 13357 7188 13369 7191
rect 13320 7160 13369 7188
rect 13320 7148 13326 7160
rect 13357 7157 13369 7160
rect 13403 7157 13415 7191
rect 13648 7188 13676 7228
rect 13832 7188 13860 7296
rect 14016 7256 14044 7432
rect 14384 7432 14780 7460
rect 14182 7392 14188 7404
rect 14143 7364 14188 7392
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 14384 7401 14412 7432
rect 14348 7395 14412 7401
rect 14348 7361 14360 7395
rect 14394 7364 14412 7395
rect 14394 7361 14406 7364
rect 14348 7355 14406 7361
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 14642 7401 14648 7404
rect 14599 7395 14648 7401
rect 14516 7364 14561 7392
rect 14516 7352 14522 7364
rect 14599 7361 14611 7395
rect 14645 7361 14648 7395
rect 14599 7355 14648 7361
rect 14642 7352 14648 7355
rect 14700 7352 14706 7404
rect 14752 7392 14780 7432
rect 14829 7429 14841 7463
rect 14875 7460 14887 7463
rect 15010 7460 15016 7472
rect 14875 7432 15016 7460
rect 14875 7429 14887 7432
rect 14829 7423 14887 7429
rect 15010 7420 15016 7432
rect 15068 7420 15074 7472
rect 15378 7460 15384 7472
rect 15339 7432 15384 7460
rect 15378 7420 15384 7432
rect 15436 7420 15442 7472
rect 16574 7420 16580 7472
rect 16632 7460 16638 7472
rect 17190 7463 17248 7469
rect 17190 7460 17202 7463
rect 16632 7432 17202 7460
rect 16632 7420 16638 7432
rect 17190 7429 17202 7432
rect 17236 7429 17248 7463
rect 17190 7423 17248 7429
rect 14918 7392 14924 7404
rect 14752 7364 14924 7392
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15102 7392 15108 7404
rect 15063 7364 15108 7392
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 15286 7392 15292 7404
rect 15247 7364 15292 7392
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 16206 7392 16212 7404
rect 16163 7364 16212 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 15488 7324 15516 7355
rect 16206 7352 16212 7364
rect 16264 7352 16270 7404
rect 16758 7352 16764 7404
rect 16816 7392 16822 7404
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16816 7364 16957 7392
rect 16816 7352 16822 7364
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 15068 7296 15516 7324
rect 16301 7327 16359 7333
rect 15068 7284 15074 7296
rect 16301 7293 16313 7327
rect 16347 7324 16359 7327
rect 16482 7324 16488 7336
rect 16347 7296 16488 7324
rect 16347 7293 16359 7296
rect 16301 7287 16359 7293
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 14016 7228 14412 7256
rect 13648 7160 13860 7188
rect 14384 7188 14412 7228
rect 14550 7216 14556 7268
rect 14608 7256 14614 7268
rect 14608 7228 16896 7256
rect 14608 7216 14614 7228
rect 16868 7200 16896 7228
rect 15102 7188 15108 7200
rect 14384 7160 15108 7188
rect 13357 7151 13415 7157
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 15657 7191 15715 7197
rect 15657 7188 15669 7191
rect 15436 7160 15669 7188
rect 15436 7148 15442 7160
rect 15657 7157 15669 7160
rect 15703 7157 15715 7191
rect 15657 7151 15715 7157
rect 15933 7191 15991 7197
rect 15933 7157 15945 7191
rect 15979 7188 15991 7191
rect 16114 7188 16120 7200
rect 15979 7160 16120 7188
rect 15979 7157 15991 7160
rect 15933 7151 15991 7157
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 16850 7148 16856 7200
rect 16908 7188 16914 7200
rect 18325 7191 18383 7197
rect 18325 7188 18337 7191
rect 16908 7160 18337 7188
rect 16908 7148 16914 7160
rect 18325 7157 18337 7160
rect 18371 7157 18383 7191
rect 18325 7151 18383 7157
rect 1104 7098 18860 7120
rect 1104 7046 3915 7098
rect 3967 7046 3979 7098
rect 4031 7046 4043 7098
rect 4095 7046 4107 7098
rect 4159 7046 4171 7098
rect 4223 7046 9846 7098
rect 9898 7046 9910 7098
rect 9962 7046 9974 7098
rect 10026 7046 10038 7098
rect 10090 7046 10102 7098
rect 10154 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 15904 7098
rect 15956 7046 15968 7098
rect 16020 7046 16032 7098
rect 16084 7046 18860 7098
rect 1104 7024 18860 7046
rect 1949 6987 2007 6993
rect 1949 6953 1961 6987
rect 1995 6984 2007 6987
rect 2038 6984 2044 6996
rect 1995 6956 2044 6984
rect 1995 6953 2007 6956
rect 1949 6947 2007 6953
rect 2038 6944 2044 6956
rect 2096 6944 2102 6996
rect 4890 6984 4896 6996
rect 4851 6956 4896 6984
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 8113 6987 8171 6993
rect 8113 6953 8125 6987
rect 8159 6953 8171 6987
rect 8938 6984 8944 6996
rect 8899 6956 8944 6984
rect 8113 6947 8171 6953
rect 4798 6916 4804 6928
rect 4172 6888 4804 6916
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 1820 6820 2329 6848
rect 1820 6808 1826 6820
rect 2317 6817 2329 6820
rect 2363 6848 2375 6851
rect 2682 6848 2688 6860
rect 2363 6820 2688 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 3053 6851 3111 6857
rect 3053 6817 3065 6851
rect 3099 6848 3111 6851
rect 3510 6848 3516 6860
rect 3099 6820 3516 6848
rect 3099 6817 3111 6820
rect 3053 6811 3111 6817
rect 3510 6808 3516 6820
rect 3568 6848 3574 6860
rect 4172 6848 4200 6888
rect 4798 6876 4804 6888
rect 4856 6876 4862 6928
rect 8128 6916 8156 6947
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 11422 6944 11428 6996
rect 11480 6984 11486 6996
rect 11480 6956 12434 6984
rect 11480 6944 11486 6956
rect 8202 6916 8208 6928
rect 8115 6888 8208 6916
rect 8202 6876 8208 6888
rect 8260 6916 8266 6928
rect 9398 6916 9404 6928
rect 8260 6888 9404 6916
rect 8260 6876 8266 6888
rect 9398 6876 9404 6888
rect 9456 6876 9462 6928
rect 12253 6919 12311 6925
rect 12253 6916 12265 6919
rect 10336 6888 12265 6916
rect 4338 6848 4344 6860
rect 3568 6820 4200 6848
rect 4299 6820 4344 6848
rect 3568 6808 3574 6820
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7282 6848 7288 6860
rect 6595 6820 7288 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 7282 6808 7288 6820
rect 7340 6808 7346 6860
rect 9217 6851 9275 6857
rect 9217 6817 9229 6851
rect 9263 6848 9275 6851
rect 10336 6848 10364 6888
rect 12253 6885 12265 6888
rect 12299 6885 12311 6919
rect 12406 6916 12434 6956
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 14550 6984 14556 6996
rect 13504 6956 14556 6984
rect 13504 6944 13510 6956
rect 14550 6944 14556 6956
rect 14608 6944 14614 6996
rect 14918 6984 14924 6996
rect 14879 6956 14924 6984
rect 14918 6944 14924 6956
rect 14976 6944 14982 6996
rect 16206 6944 16212 6996
rect 16264 6984 16270 6996
rect 16301 6987 16359 6993
rect 16301 6984 16313 6987
rect 16264 6956 16313 6984
rect 16264 6944 16270 6956
rect 16301 6953 16313 6956
rect 16347 6953 16359 6987
rect 16301 6947 16359 6953
rect 12406 6888 16896 6916
rect 12253 6879 12311 6885
rect 9263 6820 10364 6848
rect 9263 6817 9275 6820
rect 9217 6811 9275 6817
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3237 6783 3295 6789
rect 2832 6752 2877 6780
rect 2832 6740 2838 6752
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 4154 6780 4160 6792
rect 3283 6752 4160 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 6270 6740 6276 6792
rect 6328 6789 6334 6792
rect 6328 6780 6340 6789
rect 6328 6752 6373 6780
rect 6328 6743 6340 6752
rect 6328 6740 6334 6743
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7708 6752 7757 6780
rect 7708 6740 7714 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 9585 6783 9643 6789
rect 9585 6749 9597 6783
rect 9631 6780 9643 6783
rect 9674 6780 9680 6792
rect 9631 6752 9680 6780
rect 9631 6749 9643 6752
rect 9585 6743 9643 6749
rect 9674 6740 9680 6752
rect 9732 6780 9738 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9732 6752 9873 6780
rect 9732 6740 9738 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 10042 6780 10048 6792
rect 10003 6752 10048 6780
rect 9861 6743 9919 6749
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10336 6780 10364 6820
rect 11698 6808 11704 6860
rect 11756 6848 11762 6860
rect 12342 6848 12348 6860
rect 11756 6820 11928 6848
rect 12303 6820 12348 6848
rect 11756 6808 11762 6820
rect 10413 6783 10471 6789
rect 10284 6752 10377 6780
rect 10284 6740 10290 6752
rect 10413 6749 10425 6783
rect 10459 6780 10471 6783
rect 11054 6780 11060 6792
rect 10459 6752 11060 6780
rect 10459 6749 10471 6752
rect 10413 6743 10471 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 11388 6752 11437 6780
rect 11388 6740 11394 6752
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 11790 6780 11796 6792
rect 11751 6752 11796 6780
rect 11425 6743 11483 6749
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 11900 6780 11928 6820
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 12434 6808 12440 6860
rect 12492 6808 12498 6860
rect 12529 6851 12587 6857
rect 12529 6817 12541 6851
rect 12575 6848 12587 6851
rect 12710 6848 12716 6860
rect 12575 6820 12716 6848
rect 12575 6817 12587 6820
rect 12529 6811 12587 6817
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 12805 6851 12863 6857
rect 12805 6817 12817 6851
rect 12851 6848 12863 6851
rect 13814 6848 13820 6860
rect 12851 6820 13820 6848
rect 12851 6817 12863 6820
rect 12805 6811 12863 6817
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 11900 6752 12265 6780
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 12452 6780 12480 6808
rect 12820 6780 12848 6811
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 13906 6808 13912 6860
rect 13964 6808 13970 6860
rect 14274 6808 14280 6860
rect 14332 6848 14338 6860
rect 15010 6848 15016 6860
rect 14332 6820 15016 6848
rect 14332 6808 14338 6820
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 15620 6820 16252 6848
rect 15620 6808 15626 6820
rect 12452 6752 12848 6780
rect 13081 6783 13139 6789
rect 12253 6743 12311 6749
rect 13081 6749 13093 6783
rect 13127 6780 13139 6783
rect 13446 6780 13452 6792
rect 13127 6752 13452 6780
rect 13127 6749 13139 6752
rect 13081 6743 13139 6749
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 13924 6780 13952 6808
rect 14113 6783 14171 6789
rect 14113 6780 14125 6783
rect 13924 6752 14125 6780
rect 14113 6749 14125 6752
rect 14159 6749 14171 6783
rect 14113 6743 14171 6749
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6780 14519 6783
rect 14550 6780 14556 6792
rect 14507 6752 14556 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 14550 6740 14556 6752
rect 14608 6780 14614 6792
rect 14918 6780 14924 6792
rect 14608 6752 14924 6780
rect 14608 6740 14614 6752
rect 14918 6740 14924 6752
rect 14976 6780 14982 6792
rect 15105 6783 15163 6789
rect 15105 6780 15117 6783
rect 14976 6752 15117 6780
rect 14976 6740 14982 6752
rect 15105 6749 15117 6752
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 15197 6783 15255 6789
rect 15197 6749 15209 6783
rect 15243 6749 15255 6783
rect 15378 6780 15384 6792
rect 15339 6752 15384 6780
rect 15197 6743 15255 6749
rect 3421 6715 3479 6721
rect 3421 6681 3433 6715
rect 3467 6712 3479 6715
rect 5350 6712 5356 6724
rect 3467 6684 5356 6712
rect 3467 6681 3479 6684
rect 3421 6675 3479 6681
rect 5350 6672 5356 6684
rect 5408 6672 5414 6724
rect 7558 6672 7564 6724
rect 7616 6712 7622 6724
rect 9100 6715 9158 6721
rect 9100 6712 9112 6715
rect 7616 6684 9112 6712
rect 7616 6672 7622 6684
rect 9100 6681 9112 6684
rect 9146 6681 9158 6715
rect 9100 6675 9158 6681
rect 10318 6672 10324 6724
rect 10376 6712 10382 6724
rect 10502 6712 10508 6724
rect 10376 6684 10508 6712
rect 10376 6672 10382 6684
rect 10502 6672 10508 6684
rect 10560 6712 10566 6724
rect 10781 6715 10839 6721
rect 10781 6712 10793 6715
rect 10560 6684 10793 6712
rect 10560 6672 10566 6684
rect 10781 6681 10793 6684
rect 10827 6712 10839 6715
rect 11609 6715 11667 6721
rect 11609 6712 11621 6715
rect 10827 6684 11621 6712
rect 10827 6681 10839 6684
rect 10781 6675 10839 6681
rect 11609 6681 11621 6684
rect 11655 6681 11667 6715
rect 11609 6675 11667 6681
rect 11701 6715 11759 6721
rect 11701 6681 11713 6715
rect 11747 6681 11759 6715
rect 11701 6675 11759 6681
rect 2590 6644 2596 6656
rect 2551 6616 2596 6644
rect 2590 6604 2596 6616
rect 2648 6604 2654 6656
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 4433 6647 4491 6653
rect 4433 6644 4445 6647
rect 3108 6616 4445 6644
rect 3108 6604 3114 6616
rect 4433 6613 4445 6616
rect 4479 6613 4491 6647
rect 4433 6607 4491 6613
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 5166 6644 5172 6656
rect 4580 6616 4625 6644
rect 5127 6616 5172 6644
rect 4580 6604 4586 6616
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 8110 6644 8116 6656
rect 8071 6616 8116 6644
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 8294 6644 8300 6656
rect 8255 6616 8300 6644
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 9309 6647 9367 6653
rect 9309 6613 9321 6647
rect 9355 6644 9367 6647
rect 10134 6644 10140 6656
rect 9355 6616 10140 6644
rect 9355 6613 9367 6616
rect 9309 6607 9367 6613
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 10870 6644 10876 6656
rect 10831 6616 10876 6644
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 11716 6644 11744 6675
rect 12986 6672 12992 6724
rect 13044 6712 13050 6724
rect 13814 6712 13820 6724
rect 13044 6684 13820 6712
rect 13044 6672 13050 6684
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 13906 6672 13912 6724
rect 13964 6712 13970 6724
rect 14277 6715 14335 6721
rect 14277 6712 14289 6715
rect 13964 6684 14289 6712
rect 13964 6672 13970 6684
rect 14277 6681 14289 6684
rect 14323 6681 14335 6715
rect 14277 6675 14335 6681
rect 14369 6715 14427 6721
rect 14369 6681 14381 6715
rect 14415 6712 14427 6715
rect 15010 6712 15016 6724
rect 14415 6684 15016 6712
rect 14415 6681 14427 6684
rect 14369 6675 14427 6681
rect 15010 6672 15016 6684
rect 15068 6672 15074 6724
rect 11790 6644 11796 6656
rect 11716 6616 11796 6644
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 11974 6644 11980 6656
rect 11935 6616 11980 6644
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 12618 6644 12624 6656
rect 12308 6616 12624 6644
rect 12308 6604 12314 6616
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 14608 6616 14657 6644
rect 14608 6604 14614 6616
rect 14645 6613 14657 6616
rect 14691 6613 14703 6647
rect 15212 6644 15240 6743
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 15473 6783 15531 6789
rect 15473 6749 15485 6783
rect 15519 6749 15531 6783
rect 15473 6743 15531 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6780 15899 6783
rect 16114 6780 16120 6792
rect 15887 6752 16120 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 15488 6712 15516 6743
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16224 6780 16252 6820
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 16868 6857 16896 6888
rect 16761 6851 16819 6857
rect 16761 6848 16773 6851
rect 16724 6820 16773 6848
rect 16724 6808 16730 6820
rect 16761 6817 16773 6820
rect 16807 6817 16819 6851
rect 16761 6811 16819 6817
rect 16853 6851 16911 6857
rect 16853 6817 16865 6851
rect 16899 6848 16911 6851
rect 16942 6848 16948 6860
rect 16899 6820 16948 6848
rect 16899 6817 16911 6820
rect 16853 6811 16911 6817
rect 16942 6808 16948 6820
rect 17000 6848 17006 6860
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 17000 6820 17877 6848
rect 17000 6808 17006 6820
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 16224 6752 17693 6780
rect 17681 6749 17693 6752
rect 17727 6780 17739 6783
rect 18230 6780 18236 6792
rect 17727 6752 18236 6780
rect 17727 6749 17739 6752
rect 17681 6743 17739 6749
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 15562 6712 15568 6724
rect 15488 6684 15568 6712
rect 15562 6672 15568 6684
rect 15620 6672 15626 6724
rect 16206 6672 16212 6724
rect 16264 6712 16270 6724
rect 17773 6715 17831 6721
rect 16264 6684 17356 6712
rect 16264 6672 16270 6684
rect 15654 6644 15660 6656
rect 15212 6616 15660 6644
rect 14645 6607 14703 6613
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 16025 6647 16083 6653
rect 16025 6613 16037 6647
rect 16071 6644 16083 6647
rect 16574 6644 16580 6656
rect 16071 6616 16580 6644
rect 16071 6613 16083 6616
rect 16025 6607 16083 6613
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 16669 6647 16727 6653
rect 16669 6613 16681 6647
rect 16715 6644 16727 6647
rect 16850 6644 16856 6656
rect 16715 6616 16856 6644
rect 16715 6613 16727 6616
rect 16669 6607 16727 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 17328 6653 17356 6684
rect 17773 6681 17785 6715
rect 17819 6712 17831 6715
rect 17862 6712 17868 6724
rect 17819 6684 17868 6712
rect 17819 6681 17831 6684
rect 17773 6675 17831 6681
rect 17862 6672 17868 6684
rect 17920 6672 17926 6724
rect 17313 6647 17371 6653
rect 17313 6613 17325 6647
rect 17359 6613 17371 6647
rect 17313 6607 17371 6613
rect 1104 6554 18860 6576
rect 1104 6502 6880 6554
rect 6932 6502 6944 6554
rect 6996 6502 7008 6554
rect 7060 6502 7072 6554
rect 7124 6502 7136 6554
rect 7188 6502 12811 6554
rect 12863 6502 12875 6554
rect 12927 6502 12939 6554
rect 12991 6502 13003 6554
rect 13055 6502 13067 6554
rect 13119 6502 18860 6554
rect 1104 6480 18860 6502
rect 2869 6443 2927 6449
rect 2869 6409 2881 6443
rect 2915 6440 2927 6443
rect 3050 6440 3056 6452
rect 2915 6412 3056 6440
rect 2915 6409 2927 6412
rect 2869 6403 2927 6409
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 4154 6440 4160 6452
rect 4115 6412 4160 6440
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 4525 6443 4583 6449
rect 4525 6409 4537 6443
rect 4571 6440 4583 6443
rect 5166 6440 5172 6452
rect 4571 6412 5172 6440
rect 4571 6409 4583 6412
rect 4525 6403 4583 6409
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6440 6883 6443
rect 7282 6440 7288 6452
rect 6871 6412 7288 6440
rect 6871 6409 6883 6412
rect 6825 6403 6883 6409
rect 6932 6384 6960 6412
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 7558 6440 7564 6452
rect 7519 6412 7564 6440
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 8352 6412 9413 6440
rect 8352 6400 8358 6412
rect 9401 6409 9413 6412
rect 9447 6440 9459 6443
rect 10042 6440 10048 6452
rect 9447 6412 10048 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 10284 6412 10333 6440
rect 10284 6400 10290 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 11146 6440 11152 6452
rect 11107 6412 11152 6440
rect 10321 6403 10379 6409
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 12342 6440 12348 6452
rect 11532 6412 12348 6440
rect 2958 6372 2964 6384
rect 1688 6344 2774 6372
rect 2871 6344 2964 6372
rect 1688 6313 1716 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 2746 6304 2774 6344
rect 2958 6332 2964 6344
rect 3016 6372 3022 6384
rect 4617 6375 4675 6381
rect 4617 6372 4629 6375
rect 3016 6344 4629 6372
rect 3016 6332 3022 6344
rect 4617 6341 4629 6344
rect 4663 6341 4675 6375
rect 4617 6335 4675 6341
rect 5353 6375 5411 6381
rect 5353 6341 5365 6375
rect 5399 6372 5411 6375
rect 5534 6372 5540 6384
rect 5399 6344 5540 6372
rect 5399 6341 5411 6344
rect 5353 6335 5411 6341
rect 5534 6332 5540 6344
rect 5592 6372 5598 6384
rect 6733 6375 6791 6381
rect 6733 6372 6745 6375
rect 5592 6344 6745 6372
rect 5592 6332 5598 6344
rect 6733 6341 6745 6344
rect 6779 6341 6791 6375
rect 6733 6335 6791 6341
rect 6914 6332 6920 6384
rect 6972 6332 6978 6384
rect 7193 6375 7251 6381
rect 7193 6341 7205 6375
rect 7239 6341 7251 6375
rect 7193 6335 7251 6341
rect 7409 6375 7467 6381
rect 7409 6341 7421 6375
rect 7455 6372 7467 6375
rect 8386 6372 8392 6384
rect 7455 6344 8248 6372
rect 8347 6344 8392 6372
rect 7455 6341 7467 6344
rect 7409 6335 7467 6341
rect 3697 6307 3755 6313
rect 2746 6276 3648 6304
rect 1673 6267 1731 6273
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 3142 6236 3148 6248
rect 3103 6208 3148 6236
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 3510 6236 3516 6248
rect 3471 6208 3516 6236
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 3620 6236 3648 6276
rect 3697 6273 3709 6307
rect 3743 6304 3755 6307
rect 3786 6304 3792 6316
rect 3743 6276 3792 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 3786 6264 3792 6276
rect 3844 6264 3850 6316
rect 5902 6304 5908 6316
rect 4264 6276 5764 6304
rect 5863 6276 5908 6304
rect 4264 6236 4292 6276
rect 3620 6208 4292 6236
rect 4338 6196 4344 6248
rect 4396 6236 4402 6248
rect 4709 6239 4767 6245
rect 4709 6236 4721 6239
rect 4396 6208 4721 6236
rect 4396 6196 4402 6208
rect 4709 6205 4721 6208
rect 4755 6205 4767 6239
rect 5736 6236 5764 6276
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 7208 6304 7236 6335
rect 8220 6316 8248 6344
rect 8386 6332 8392 6344
rect 8444 6332 8450 6384
rect 8570 6332 8576 6384
rect 8628 6372 8634 6384
rect 8941 6375 8999 6381
rect 8941 6372 8953 6375
rect 8628 6344 8953 6372
rect 8628 6332 8634 6344
rect 8941 6341 8953 6344
rect 8987 6341 8999 6375
rect 8941 6335 8999 6341
rect 9217 6375 9275 6381
rect 9217 6341 9229 6375
rect 9263 6372 9275 6375
rect 10244 6372 10272 6400
rect 9263 6344 10272 6372
rect 9263 6341 9275 6344
rect 9217 6335 9275 6341
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7208 6276 7941 6304
rect 7929 6273 7941 6276
rect 7975 6304 7987 6307
rect 8018 6304 8024 6316
rect 7975 6276 8024 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 7374 6236 7380 6248
rect 5736 6208 7380 6236
rect 4709 6199 4767 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 8128 6236 8156 6267
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8260 6276 8677 6304
rect 8260 6264 8266 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 10502 6304 10508 6316
rect 8812 6276 10508 6304
rect 8812 6264 8818 6276
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 10965 6264 10971 6316
rect 11023 6304 11029 6316
rect 11023 6276 11068 6304
rect 11023 6264 11029 6276
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11532 6304 11560 6412
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 15470 6440 15476 6452
rect 13004 6412 15476 6440
rect 11606 6332 11612 6384
rect 11664 6372 11670 6384
rect 11664 6344 11836 6372
rect 11664 6332 11670 6344
rect 11808 6313 11836 6344
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11204 6276 11713 6304
rect 11204 6264 11210 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11974 6304 11980 6316
rect 11935 6276 11980 6304
rect 11793 6267 11851 6273
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6304 12127 6307
rect 12250 6304 12256 6316
rect 12115 6276 12256 6304
rect 12115 6273 12127 6276
rect 12069 6267 12127 6273
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 12400 6276 12449 6304
rect 12400 6264 12406 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 12526 6264 12532 6316
rect 12584 6304 12590 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12584 6276 12909 6304
rect 12584 6264 12590 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 13004 6304 13032 6412
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 15657 6443 15715 6449
rect 15657 6409 15669 6443
rect 15703 6409 15715 6443
rect 18230 6440 18236 6452
rect 18191 6412 18236 6440
rect 15657 6403 15715 6409
rect 13170 6372 13176 6384
rect 13131 6344 13176 6372
rect 13170 6332 13176 6344
rect 13228 6332 13234 6384
rect 13906 6372 13912 6384
rect 13867 6344 13912 6372
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 14001 6375 14059 6381
rect 14001 6341 14013 6375
rect 14047 6341 14059 6375
rect 15102 6372 15108 6384
rect 14001 6335 14059 6341
rect 14568 6344 15108 6372
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 13004 6276 13093 6304
rect 12897 6267 12955 6273
rect 13081 6273 13093 6276
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6273 13323 6307
rect 13722 6304 13728 6316
rect 13683 6276 13728 6304
rect 13265 6267 13323 6273
rect 7668 6208 8156 6236
rect 9309 6239 9367 6245
rect 1578 6128 1584 6180
rect 1636 6168 1642 6180
rect 5169 6171 5227 6177
rect 5169 6168 5181 6171
rect 1636 6140 5181 6168
rect 1636 6128 1642 6140
rect 5169 6137 5181 6140
rect 5215 6168 5227 6171
rect 5258 6168 5264 6180
rect 5215 6140 5264 6168
rect 5215 6137 5227 6140
rect 5169 6131 5227 6137
rect 5258 6128 5264 6140
rect 5316 6128 5322 6180
rect 7668 6112 7696 6208
rect 9309 6205 9321 6239
rect 9355 6205 9367 6239
rect 9309 6199 9367 6205
rect 9324 6168 9352 6199
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9732 6208 9965 6236
rect 9732 6196 9738 6208
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 10781 6239 10839 6245
rect 10781 6205 10793 6239
rect 10827 6205 10839 6239
rect 13280 6236 13308 6267
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 14016 6248 14044 6335
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6304 14151 6307
rect 14274 6304 14280 6316
rect 14139 6276 14280 6304
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 14568 6313 14596 6344
rect 15102 6332 15108 6344
rect 15160 6372 15166 6384
rect 15562 6372 15568 6384
rect 15160 6344 15568 6372
rect 15160 6332 15166 6344
rect 15562 6332 15568 6344
rect 15620 6332 15626 6384
rect 15672 6372 15700 6403
rect 18230 6400 18236 6412
rect 18288 6400 18294 6452
rect 17098 6375 17156 6381
rect 17098 6372 17110 6375
rect 15672 6344 17110 6372
rect 17098 6341 17110 6344
rect 17144 6341 17156 6375
rect 17098 6335 17156 6341
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 13998 6236 14004 6248
rect 13280 6208 14004 6236
rect 10781 6199 10839 6205
rect 10134 6168 10140 6180
rect 9324 6140 10140 6168
rect 10134 6128 10140 6140
rect 10192 6168 10198 6180
rect 10686 6168 10692 6180
rect 10192 6140 10692 6168
rect 10192 6128 10198 6140
rect 1946 6060 1952 6112
rect 2004 6100 2010 6112
rect 2501 6103 2559 6109
rect 2501 6100 2513 6103
rect 2004 6072 2513 6100
rect 2004 6060 2010 6072
rect 2501 6069 2513 6072
rect 2547 6069 2559 6103
rect 2501 6063 2559 6069
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 3881 6103 3939 6109
rect 3881 6100 3893 6103
rect 3844 6072 3893 6100
rect 3844 6060 3850 6072
rect 3881 6069 3893 6072
rect 3927 6069 3939 6103
rect 3881 6063 3939 6069
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 5721 6103 5779 6109
rect 5721 6100 5733 6103
rect 5592 6072 5733 6100
rect 5592 6060 5598 6072
rect 5721 6069 5733 6072
rect 5767 6069 5779 6103
rect 5721 6063 5779 6069
rect 7377 6103 7435 6109
rect 7377 6069 7389 6103
rect 7423 6100 7435 6103
rect 7650 6100 7656 6112
rect 7423 6072 7656 6100
rect 7423 6069 7435 6072
rect 7377 6063 7435 6069
rect 7650 6060 7656 6072
rect 7708 6060 7714 6112
rect 10336 6109 10364 6140
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 10321 6103 10379 6109
rect 10321 6069 10333 6103
rect 10367 6069 10379 6103
rect 10502 6100 10508 6112
rect 10463 6072 10508 6100
rect 10321 6063 10379 6069
rect 10502 6060 10508 6072
rect 10560 6100 10566 6112
rect 10796 6100 10824 6199
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14660 6236 14688 6267
rect 14734 6264 14740 6316
rect 14792 6304 14798 6316
rect 14829 6307 14887 6313
rect 14829 6304 14841 6307
rect 14792 6276 14841 6304
rect 14792 6264 14798 6276
rect 14829 6273 14841 6276
rect 14875 6273 14887 6307
rect 14829 6267 14887 6273
rect 14918 6264 14924 6316
rect 14976 6304 14982 6316
rect 15473 6307 15531 6313
rect 14976 6276 15021 6304
rect 14976 6264 14982 6276
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 15933 6307 15991 6313
rect 15933 6304 15945 6307
rect 15519 6276 15945 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 15933 6273 15945 6276
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 16206 6304 16212 6316
rect 16163 6276 16212 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 16758 6264 16764 6316
rect 16816 6304 16822 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16816 6276 16865 6304
rect 16816 6264 16822 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 14292 6208 14688 6236
rect 12621 6171 12679 6177
rect 12621 6137 12633 6171
rect 12667 6168 12679 6171
rect 13354 6168 13360 6180
rect 12667 6140 13360 6168
rect 12667 6137 12679 6140
rect 12621 6131 12679 6137
rect 13354 6128 13360 6140
rect 13412 6168 13418 6180
rect 14292 6177 14320 6208
rect 15654 6196 15660 6248
rect 15712 6236 15718 6248
rect 16301 6239 16359 6245
rect 16301 6236 16313 6239
rect 15712 6208 16313 6236
rect 15712 6196 15718 6208
rect 16301 6205 16313 6208
rect 16347 6236 16359 6239
rect 16482 6236 16488 6248
rect 16347 6208 16488 6236
rect 16347 6205 16359 6208
rect 16301 6199 16359 6205
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 14277 6171 14335 6177
rect 13412 6140 14044 6168
rect 13412 6128 13418 6140
rect 11514 6100 11520 6112
rect 10560 6072 10824 6100
rect 11475 6072 11520 6100
rect 10560 6060 10566 6072
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 13449 6103 13507 6109
rect 13449 6069 13461 6103
rect 13495 6100 13507 6103
rect 13722 6100 13728 6112
rect 13495 6072 13728 6100
rect 13495 6069 13507 6072
rect 13449 6063 13507 6069
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 14016 6100 14044 6140
rect 14277 6137 14289 6171
rect 14323 6137 14335 6171
rect 14277 6131 14335 6137
rect 14458 6100 14464 6112
rect 14016 6072 14464 6100
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 15105 6103 15163 6109
rect 15105 6069 15117 6103
rect 15151 6100 15163 6103
rect 15562 6100 15568 6112
rect 15151 6072 15568 6100
rect 15151 6069 15163 6072
rect 15105 6063 15163 6069
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 1104 6010 18860 6032
rect 1104 5958 3915 6010
rect 3967 5958 3979 6010
rect 4031 5958 4043 6010
rect 4095 5958 4107 6010
rect 4159 5958 4171 6010
rect 4223 5958 9846 6010
rect 9898 5958 9910 6010
rect 9962 5958 9974 6010
rect 10026 5958 10038 6010
rect 10090 5958 10102 6010
rect 10154 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 15904 6010
rect 15956 5958 15968 6010
rect 16020 5958 16032 6010
rect 16084 5958 18860 6010
rect 1104 5936 18860 5958
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 2958 5896 2964 5908
rect 2915 5868 2964 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3752 5868 3893 5896
rect 3752 5856 3758 5868
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 3881 5859 3939 5865
rect 4522 5856 4528 5908
rect 4580 5896 4586 5908
rect 6641 5899 6699 5905
rect 6641 5896 6653 5899
rect 4580 5868 6653 5896
rect 4580 5856 4586 5868
rect 6641 5865 6653 5868
rect 6687 5896 6699 5899
rect 10318 5896 10324 5908
rect 6687 5868 10180 5896
rect 10279 5868 10324 5896
rect 6687 5865 6699 5868
rect 6641 5859 6699 5865
rect 8846 5788 8852 5840
rect 8904 5828 8910 5840
rect 9674 5828 9680 5840
rect 8904 5800 9680 5828
rect 8904 5788 8910 5800
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 10152 5828 10180 5868
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 10870 5896 10876 5908
rect 10744 5868 10876 5896
rect 10744 5856 10750 5868
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 11977 5899 12035 5905
rect 11977 5896 11989 5899
rect 11940 5868 11989 5896
rect 11940 5856 11946 5868
rect 11977 5865 11989 5868
rect 12023 5865 12035 5899
rect 11977 5859 12035 5865
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 12897 5899 12955 5905
rect 12897 5896 12909 5899
rect 12676 5868 12909 5896
rect 12676 5856 12682 5868
rect 12897 5865 12909 5868
rect 12943 5865 12955 5899
rect 12897 5859 12955 5865
rect 11149 5831 11207 5837
rect 9784 5800 10088 5828
rect 10152 5800 10824 5828
rect 4338 5720 4344 5772
rect 4396 5760 4402 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4396 5732 4445 5760
rect 4396 5720 4402 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 5258 5760 5264 5772
rect 5219 5732 5264 5760
rect 4433 5723 4491 5729
rect 5258 5720 5264 5732
rect 5316 5720 5322 5772
rect 6914 5760 6920 5772
rect 6875 5732 6920 5760
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 9784 5760 9812 5800
rect 9508 5732 9812 5760
rect 10060 5760 10088 5800
rect 10502 5760 10508 5772
rect 10060 5732 10508 5760
rect 1489 5695 1547 5701
rect 1489 5661 1501 5695
rect 1535 5692 1547 5695
rect 1578 5692 1584 5704
rect 1535 5664 1584 5692
rect 1535 5661 1547 5664
rect 1489 5655 1547 5661
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 1756 5695 1814 5701
rect 1756 5661 1768 5695
rect 1802 5692 1814 5695
rect 2590 5692 2596 5704
rect 1802 5664 2596 5692
rect 1802 5661 1814 5664
rect 1756 5655 1814 5661
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4982 5692 4988 5704
rect 4295 5664 4988 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5534 5701 5540 5704
rect 5528 5692 5540 5701
rect 5495 5664 5540 5692
rect 5528 5655 5540 5664
rect 5534 5652 5540 5655
rect 5592 5652 5598 5704
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 9508 5701 9536 5732
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 10796 5769 10824 5800
rect 11149 5797 11161 5831
rect 11195 5828 11207 5831
rect 14642 5828 14648 5840
rect 11195 5800 14648 5828
rect 11195 5797 11207 5800
rect 11149 5791 11207 5797
rect 14642 5788 14648 5800
rect 14700 5788 14706 5840
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5729 10839 5763
rect 11701 5763 11759 5769
rect 11701 5760 11713 5763
rect 10781 5723 10839 5729
rect 10888 5732 11713 5760
rect 9309 5695 9367 5701
rect 9309 5692 9321 5695
rect 8444 5664 9321 5692
rect 8444 5652 8450 5664
rect 9309 5661 9321 5664
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5661 9551 5695
rect 10137 5695 10195 5701
rect 9493 5655 9551 5661
rect 9600 5692 9720 5694
rect 10137 5692 10149 5695
rect 9600 5666 10149 5692
rect 7184 5627 7242 5633
rect 7184 5593 7196 5627
rect 7230 5624 7242 5627
rect 7466 5624 7472 5636
rect 7230 5596 7472 5624
rect 7230 5593 7242 5596
rect 7184 5587 7242 5593
rect 7466 5584 7472 5596
rect 7524 5584 7530 5636
rect 9324 5624 9352 5655
rect 9600 5624 9628 5666
rect 9692 5664 10149 5666
rect 10137 5661 10149 5664
rect 10183 5692 10195 5695
rect 10183 5664 10364 5692
rect 10183 5661 10195 5664
rect 10137 5655 10195 5661
rect 9324 5596 9628 5624
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 9769 5627 9827 5633
rect 9769 5624 9781 5627
rect 9732 5596 9781 5624
rect 9732 5584 9738 5596
rect 9769 5593 9781 5596
rect 9815 5593 9827 5627
rect 9950 5624 9956 5636
rect 9911 5596 9956 5624
rect 9769 5587 9827 5593
rect 9950 5584 9956 5596
rect 10008 5584 10014 5636
rect 10226 5624 10232 5636
rect 10152 5596 10232 5624
rect 4338 5516 4344 5568
rect 4396 5556 4402 5568
rect 8294 5556 8300 5568
rect 4396 5528 4441 5556
rect 8255 5528 8300 5556
rect 4396 5516 4402 5528
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 9493 5559 9551 5565
rect 9493 5525 9505 5559
rect 9539 5556 9551 5559
rect 9858 5556 9864 5568
rect 9539 5528 9864 5556
rect 9539 5525 9551 5528
rect 9493 5519 9551 5525
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 10045 5559 10103 5565
rect 10045 5525 10057 5559
rect 10091 5556 10103 5559
rect 10152 5556 10180 5596
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 10091 5528 10180 5556
rect 10336 5556 10364 5664
rect 10520 5624 10548 5720
rect 10686 5692 10692 5704
rect 10647 5664 10692 5692
rect 10686 5652 10692 5664
rect 10744 5652 10750 5704
rect 10888 5701 10916 5732
rect 11701 5729 11713 5732
rect 11747 5729 11759 5763
rect 11701 5723 11759 5729
rect 12066 5720 12072 5772
rect 12124 5760 12130 5772
rect 12253 5763 12311 5769
rect 12253 5760 12265 5763
rect 12124 5732 12265 5760
rect 12124 5720 12130 5732
rect 12253 5729 12265 5732
rect 12299 5729 12311 5763
rect 16942 5760 16948 5772
rect 16903 5732 16948 5760
rect 12253 5723 12311 5729
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 17773 5763 17831 5769
rect 17773 5760 17785 5763
rect 17144 5732 17785 5760
rect 17144 5704 17172 5732
rect 17773 5729 17785 5732
rect 17819 5729 17831 5763
rect 17773 5723 17831 5729
rect 10873 5695 10931 5701
rect 10873 5661 10885 5695
rect 10919 5661 10931 5695
rect 10873 5655 10931 5661
rect 10888 5624 10916 5655
rect 10962 5652 10968 5704
rect 11020 5701 11026 5704
rect 11020 5692 11031 5701
rect 11020 5664 11113 5692
rect 11020 5655 11031 5664
rect 11020 5652 11026 5655
rect 11146 5652 11152 5704
rect 11204 5692 11210 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11204 5664 11529 5692
rect 11204 5652 11210 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5661 11667 5695
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11609 5655 11667 5661
rect 11716 5664 11805 5692
rect 10520 5596 10916 5624
rect 10980 5556 11008 5652
rect 11054 5584 11060 5636
rect 11112 5624 11118 5636
rect 11624 5624 11652 5655
rect 11112 5596 11652 5624
rect 11112 5584 11118 5596
rect 11716 5556 11744 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 13262 5692 13268 5704
rect 12492 5664 12537 5692
rect 13223 5664 13268 5692
rect 12492 5652 12498 5664
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 13722 5692 13728 5704
rect 13587 5664 13728 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 14277 5695 14335 5701
rect 13872 5664 14228 5692
rect 13872 5652 13878 5664
rect 12158 5584 12164 5636
rect 12216 5624 12222 5636
rect 14093 5627 14151 5633
rect 14093 5624 14105 5627
rect 12216 5596 14105 5624
rect 12216 5584 12222 5596
rect 14093 5593 14105 5596
rect 14139 5593 14151 5627
rect 14200 5624 14228 5664
rect 14277 5661 14289 5695
rect 14323 5692 14335 5695
rect 14366 5692 14372 5704
rect 14323 5664 14372 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 14826 5692 14832 5704
rect 14783 5664 14832 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 16666 5692 16672 5704
rect 14936 5664 16672 5692
rect 14936 5624 14964 5664
rect 16666 5652 16672 5664
rect 16724 5692 16730 5704
rect 16761 5695 16819 5701
rect 16761 5692 16773 5695
rect 16724 5664 16773 5692
rect 16724 5652 16730 5664
rect 16761 5661 16773 5664
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 16853 5695 16911 5701
rect 16853 5661 16865 5695
rect 16899 5692 16911 5695
rect 17126 5692 17132 5704
rect 16899 5664 17132 5692
rect 16899 5661 16911 5664
rect 16853 5655 16911 5661
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 14200 5596 14964 5624
rect 15004 5627 15062 5633
rect 14093 5587 14151 5593
rect 15004 5593 15016 5627
rect 15050 5624 15062 5627
rect 15102 5624 15108 5636
rect 15050 5596 15108 5624
rect 15050 5593 15062 5596
rect 15004 5587 15062 5593
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 12618 5556 12624 5568
rect 10336 5528 11744 5556
rect 12579 5528 12624 5556
rect 10091 5525 10103 5528
rect 10045 5519 10103 5525
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 13354 5556 13360 5568
rect 13315 5528 13360 5556
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 13722 5556 13728 5568
rect 13683 5528 13728 5556
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 16117 5559 16175 5565
rect 16117 5556 16129 5559
rect 15252 5528 16129 5556
rect 15252 5516 15258 5528
rect 16117 5525 16129 5528
rect 16163 5556 16175 5559
rect 16206 5556 16212 5568
rect 16163 5528 16212 5556
rect 16163 5525 16175 5528
rect 16117 5519 16175 5525
rect 16206 5516 16212 5528
rect 16264 5516 16270 5568
rect 16390 5556 16396 5568
rect 16351 5528 16396 5556
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 1104 5466 18860 5488
rect 1104 5414 6880 5466
rect 6932 5414 6944 5466
rect 6996 5414 7008 5466
rect 7060 5414 7072 5466
rect 7124 5414 7136 5466
rect 7188 5414 12811 5466
rect 12863 5414 12875 5466
rect 12927 5414 12939 5466
rect 12991 5414 13003 5466
rect 13055 5414 13067 5466
rect 13119 5414 18860 5466
rect 1104 5392 18860 5414
rect 1394 5352 1400 5364
rect 1355 5324 1400 5352
rect 1394 5312 1400 5324
rect 1452 5312 1458 5364
rect 2133 5355 2191 5361
rect 2133 5321 2145 5355
rect 2179 5352 2191 5355
rect 2774 5352 2780 5364
rect 2179 5324 2780 5352
rect 2179 5321 2191 5324
rect 2133 5315 2191 5321
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 2869 5355 2927 5361
rect 2869 5321 2881 5355
rect 2915 5352 2927 5355
rect 3050 5352 3056 5364
rect 2915 5324 3056 5352
rect 2915 5321 2927 5324
rect 2869 5315 2927 5321
rect 3050 5312 3056 5324
rect 3108 5352 3114 5364
rect 4338 5352 4344 5364
rect 3108 5324 4344 5352
rect 3108 5312 3114 5324
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 5353 5355 5411 5361
rect 5353 5321 5365 5355
rect 5399 5352 5411 5355
rect 5442 5352 5448 5364
rect 5399 5324 5448 5352
rect 5399 5321 5411 5324
rect 5353 5315 5411 5321
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 6365 5355 6423 5361
rect 6365 5321 6377 5355
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 6733 5355 6791 5361
rect 6733 5321 6745 5355
rect 6779 5352 6791 5355
rect 8294 5352 8300 5364
rect 6779 5324 8300 5352
rect 6779 5321 6791 5324
rect 6733 5315 6791 5321
rect 2958 5284 2964 5296
rect 2792 5256 2964 5284
rect 1762 5216 1768 5228
rect 1723 5188 1768 5216
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 1946 5216 1952 5228
rect 1907 5188 1952 5216
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 2792 5225 2820 5256
rect 2958 5244 2964 5256
rect 3016 5244 3022 5296
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5185 2835 5219
rect 2777 5179 2835 5185
rect 3694 5176 3700 5228
rect 3752 5216 3758 5228
rect 3861 5219 3919 5225
rect 3861 5216 3873 5219
rect 3752 5188 3873 5216
rect 3752 5176 3758 5188
rect 3861 5185 3873 5188
rect 3907 5185 3919 5219
rect 3861 5179 3919 5185
rect 5350 5176 5356 5228
rect 5408 5216 5414 5228
rect 5813 5219 5871 5225
rect 5408 5188 5764 5216
rect 5408 5176 5414 5188
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3142 5148 3148 5160
rect 3099 5120 3148 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5117 3663 5151
rect 3605 5111 3663 5117
rect 1578 5040 1584 5092
rect 1636 5080 1642 5092
rect 3620 5080 3648 5111
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 5629 5151 5687 5157
rect 5629 5148 5641 5151
rect 5500 5120 5641 5148
rect 5500 5108 5506 5120
rect 5629 5117 5641 5120
rect 5675 5117 5687 5151
rect 5736 5148 5764 5188
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 6380 5216 6408 5315
rect 8294 5312 8300 5324
rect 8352 5352 8358 5364
rect 11054 5352 11060 5364
rect 8352 5324 11060 5352
rect 8352 5312 8358 5324
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 13354 5352 13360 5364
rect 12032 5324 13360 5352
rect 12032 5312 12038 5324
rect 13354 5312 13360 5324
rect 13412 5352 13418 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 13412 5324 13553 5352
rect 13412 5312 13418 5324
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 15102 5352 15108 5364
rect 15063 5324 15108 5352
rect 13541 5315 13599 5321
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 16666 5312 16672 5364
rect 16724 5352 16730 5364
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 16724 5324 18061 5352
rect 16724 5312 16730 5324
rect 18049 5321 18061 5324
rect 18095 5321 18107 5355
rect 18049 5315 18107 5321
rect 9858 5244 9864 5296
rect 9916 5284 9922 5296
rect 10502 5284 10508 5296
rect 9916 5256 10508 5284
rect 9916 5244 9922 5256
rect 10502 5244 10508 5256
rect 10560 5284 10566 5296
rect 11514 5284 11520 5296
rect 10560 5256 10824 5284
rect 10560 5244 10566 5256
rect 7558 5216 7564 5228
rect 5859 5188 6408 5216
rect 6656 5188 6960 5216
rect 7519 5188 7564 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 6656 5148 6684 5188
rect 5736 5120 6684 5148
rect 5629 5111 5687 5117
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6932 5157 6960 5188
rect 7558 5176 7564 5188
rect 7616 5176 7622 5228
rect 8656 5219 8714 5225
rect 8656 5185 8668 5219
rect 8702 5216 8714 5219
rect 9766 5216 9772 5228
rect 8702 5188 9772 5216
rect 8702 5185 8714 5188
rect 8656 5179 8714 5185
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 10226 5176 10232 5228
rect 10284 5216 10290 5228
rect 10796 5225 10824 5256
rect 10888 5256 11520 5284
rect 10888 5225 10916 5256
rect 11514 5244 11520 5256
rect 11572 5244 11578 5296
rect 11790 5244 11796 5296
rect 11848 5284 11854 5296
rect 11848 5256 15792 5284
rect 11848 5244 11854 5256
rect 10689 5219 10747 5225
rect 10689 5216 10701 5219
rect 10284 5188 10701 5216
rect 10284 5176 10290 5188
rect 10689 5185 10701 5188
rect 10735 5185 10747 5219
rect 10689 5179 10747 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 11057 5219 11115 5225
rect 11057 5185 11069 5219
rect 11103 5216 11115 5219
rect 11330 5216 11336 5228
rect 11103 5188 11336 5216
rect 11103 5185 11115 5188
rect 11057 5179 11115 5185
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 12158 5216 12164 5228
rect 12119 5188 12164 5216
rect 11701 5179 11759 5185
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6788 5120 6837 5148
rect 6788 5108 6794 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 8389 5151 8447 5157
rect 8389 5148 8401 5151
rect 7340 5120 8401 5148
rect 7340 5108 7346 5120
rect 8389 5117 8401 5120
rect 8435 5117 8447 5151
rect 8389 5111 8447 5117
rect 11146 5108 11152 5160
rect 11204 5148 11210 5160
rect 11716 5148 11744 5179
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12417 5219 12475 5225
rect 12417 5216 12429 5219
rect 12308 5188 12429 5216
rect 12308 5176 12314 5188
rect 12417 5185 12429 5188
rect 12463 5185 12475 5219
rect 12417 5179 12475 5185
rect 13909 5219 13967 5225
rect 13909 5185 13921 5219
rect 13955 5216 13967 5219
rect 14182 5216 14188 5228
rect 13955 5188 14188 5216
rect 13955 5185 13967 5188
rect 13909 5179 13967 5185
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 14366 5216 14372 5228
rect 14327 5188 14372 5216
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 14550 5216 14556 5228
rect 14511 5188 14556 5216
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 14642 5176 14648 5228
rect 14700 5216 14706 5228
rect 14921 5219 14979 5225
rect 14700 5188 14745 5216
rect 14700 5176 14706 5188
rect 14921 5185 14933 5219
rect 14967 5185 14979 5219
rect 14921 5179 14979 5185
rect 15381 5219 15439 5225
rect 15381 5185 15393 5219
rect 15427 5185 15439 5219
rect 15562 5216 15568 5228
rect 15523 5188 15568 5216
rect 15381 5179 15439 5185
rect 11204 5120 11744 5148
rect 11885 5151 11943 5157
rect 11204 5108 11210 5120
rect 11885 5117 11897 5151
rect 11931 5117 11943 5151
rect 11885 5111 11943 5117
rect 4982 5080 4988 5092
rect 1636 5052 3648 5080
rect 4895 5052 4988 5080
rect 1636 5040 1642 5052
rect 4982 5040 4988 5052
rect 5040 5080 5046 5092
rect 7742 5080 7748 5092
rect 5040 5052 7748 5080
rect 5040 5040 5046 5052
rect 7742 5040 7748 5052
rect 7800 5040 7806 5092
rect 11900 5080 11928 5111
rect 14090 5108 14096 5160
rect 14148 5148 14154 5160
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 14148 5120 14749 5148
rect 14148 5108 14154 5120
rect 14737 5117 14749 5120
rect 14783 5117 14795 5151
rect 14936 5148 14964 5179
rect 15194 5148 15200 5160
rect 14936 5120 15200 5148
rect 14737 5111 14795 5117
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 10244 5052 10916 5080
rect 2406 5012 2412 5024
rect 2367 4984 2412 5012
rect 2406 4972 2412 4984
rect 2464 4972 2470 5024
rect 5997 5015 6055 5021
rect 5997 4981 6009 5015
rect 6043 5012 6055 5015
rect 6270 5012 6276 5024
rect 6043 4984 6276 5012
rect 6043 4981 6055 4984
rect 5997 4975 6055 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 7374 5012 7380 5024
rect 7335 4984 7380 5012
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9732 4984 9781 5012
rect 9732 4972 9738 4984
rect 9769 4981 9781 4984
rect 9815 5012 9827 5015
rect 10244 5012 10272 5052
rect 10410 5012 10416 5024
rect 9815 4984 10272 5012
rect 10371 4984 10416 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 10888 5012 10916 5052
rect 11348 5052 11928 5080
rect 11348 5012 11376 5052
rect 14182 5040 14188 5092
rect 14240 5080 14246 5092
rect 15396 5080 15424 5179
rect 15562 5176 15568 5188
rect 15620 5176 15626 5228
rect 15764 5225 15792 5256
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 16758 5216 16764 5228
rect 16715 5188 16764 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 14240 5052 15424 5080
rect 14240 5040 14246 5052
rect 11514 5012 11520 5024
rect 10888 4984 11376 5012
rect 11475 4984 11520 5012
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 14001 5015 14059 5021
rect 14001 4981 14013 5015
rect 14047 5012 14059 5015
rect 14090 5012 14096 5024
rect 14047 4984 14096 5012
rect 14047 4981 14059 4984
rect 14001 4975 14059 4981
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14458 4972 14464 5024
rect 14516 5012 14522 5024
rect 15672 5012 15700 5179
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 16942 5225 16948 5228
rect 16936 5179 16948 5225
rect 17000 5216 17006 5228
rect 17000 5188 17036 5216
rect 16942 5176 16948 5179
rect 17000 5176 17006 5188
rect 14516 4984 15700 5012
rect 16025 5015 16083 5021
rect 14516 4972 14522 4984
rect 16025 4981 16037 5015
rect 16071 5012 16083 5015
rect 16114 5012 16120 5024
rect 16071 4984 16120 5012
rect 16071 4981 16083 4984
rect 16025 4975 16083 4981
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 1104 4922 18860 4944
rect 1104 4870 3915 4922
rect 3967 4870 3979 4922
rect 4031 4870 4043 4922
rect 4095 4870 4107 4922
rect 4159 4870 4171 4922
rect 4223 4870 9846 4922
rect 9898 4870 9910 4922
rect 9962 4870 9974 4922
rect 10026 4870 10038 4922
rect 10090 4870 10102 4922
rect 10154 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 15904 4922
rect 15956 4870 15968 4922
rect 16020 4870 16032 4922
rect 16084 4870 18860 4922
rect 1104 4848 18860 4870
rect 3050 4808 3056 4820
rect 3011 4780 3056 4808
rect 3050 4768 3056 4780
rect 3108 4768 3114 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 3881 4811 3939 4817
rect 3881 4808 3893 4811
rect 3752 4780 3893 4808
rect 3752 4768 3758 4780
rect 3881 4777 3893 4780
rect 3927 4777 3939 4811
rect 3881 4771 3939 4777
rect 6457 4811 6515 4817
rect 6457 4777 6469 4811
rect 6503 4808 6515 4811
rect 7466 4808 7472 4820
rect 6503 4780 7472 4808
rect 6503 4777 6515 4780
rect 6457 4771 6515 4777
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 11790 4808 11796 4820
rect 7800 4780 11796 4808
rect 7800 4768 7806 4780
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 12529 4811 12587 4817
rect 12529 4808 12541 4811
rect 12492 4780 12541 4808
rect 12492 4768 12498 4780
rect 12529 4777 12541 4780
rect 12575 4777 12587 4811
rect 12529 4771 12587 4777
rect 15933 4811 15991 4817
rect 15933 4777 15945 4811
rect 15979 4808 15991 4811
rect 16206 4808 16212 4820
rect 15979 4780 16212 4808
rect 15979 4777 15991 4780
rect 15933 4771 15991 4777
rect 16206 4768 16212 4780
rect 16264 4768 16270 4820
rect 9490 4740 9496 4752
rect 9451 4712 9496 4740
rect 9490 4700 9496 4712
rect 9548 4700 9554 4752
rect 1578 4632 1584 4684
rect 1636 4672 1642 4684
rect 1673 4675 1731 4681
rect 1673 4672 1685 4675
rect 1636 4644 1685 4672
rect 1636 4632 1642 4644
rect 1673 4641 1685 4644
rect 1719 4641 1731 4675
rect 1673 4635 1731 4641
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 4893 4675 4951 4681
rect 4893 4672 4905 4675
rect 4663 4644 4905 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 4893 4641 4905 4644
rect 4939 4672 4951 4675
rect 5442 4672 5448 4684
rect 4939 4644 5448 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 5442 4632 5448 4644
rect 5500 4672 5506 4684
rect 6546 4672 6552 4684
rect 5500 4644 6552 4672
rect 5500 4632 5506 4644
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 9122 4672 9128 4684
rect 9083 4644 9128 4672
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4672 9643 4675
rect 11330 4672 11336 4684
rect 9631 4644 11336 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 3786 4564 3792 4616
rect 3844 4604 3850 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3844 4576 4077 4604
rect 3844 4564 3850 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 5074 4604 5080 4616
rect 5035 4576 5080 4604
rect 4065 4567 4123 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4604 5319 4607
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5307 4576 5733 4604
rect 5307 4573 5319 4576
rect 5261 4567 5319 4573
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 6270 4604 6276 4616
rect 6231 4576 6276 4604
rect 5721 4567 5779 4573
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4604 7159 4607
rect 7190 4604 7196 4616
rect 7147 4576 7196 4604
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 7374 4613 7380 4616
rect 7368 4604 7380 4613
rect 7335 4576 7380 4604
rect 7368 4567 7380 4576
rect 7374 4564 7380 4567
rect 7432 4564 7438 4616
rect 10428 4613 10456 4644
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 11422 4632 11428 4684
rect 11480 4672 11486 4684
rect 11885 4675 11943 4681
rect 11885 4672 11897 4675
rect 11480 4644 11897 4672
rect 11480 4632 11486 4644
rect 11885 4641 11897 4644
rect 11931 4672 11943 4675
rect 13081 4675 13139 4681
rect 13081 4672 13093 4675
rect 11931 4644 13093 4672
rect 11931 4641 11943 4644
rect 11885 4635 11943 4641
rect 13081 4641 13093 4644
rect 13127 4641 13139 4675
rect 13081 4635 13139 4641
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4573 10471 4607
rect 10594 4604 10600 4616
rect 10555 4576 10600 4604
rect 10413 4567 10471 4573
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4573 10747 4607
rect 10689 4567 10747 4573
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 1670 4496 1676 4548
rect 1728 4536 1734 4548
rect 1918 4539 1976 4545
rect 1918 4536 1930 4539
rect 1728 4508 1930 4536
rect 1728 4496 1734 4508
rect 1918 4505 1930 4508
rect 1964 4505 1976 4539
rect 3329 4539 3387 4545
rect 3329 4536 3341 4539
rect 1918 4499 1976 4505
rect 2746 4508 3341 4536
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 2746 4468 2774 4508
rect 3329 4505 3341 4508
rect 3375 4505 3387 4539
rect 3329 4499 3387 4505
rect 10502 4496 10508 4548
rect 10560 4536 10566 4548
rect 10704 4536 10732 4567
rect 10560 4508 10732 4536
rect 10560 4496 10566 4508
rect 2372 4440 2774 4468
rect 2372 4428 2378 4440
rect 4890 4428 4896 4480
rect 4948 4468 4954 4480
rect 5537 4471 5595 4477
rect 5537 4468 5549 4471
rect 4948 4440 5549 4468
rect 4948 4428 4954 4440
rect 5537 4437 5549 4440
rect 5583 4437 5595 4471
rect 8478 4468 8484 4480
rect 8391 4440 8484 4468
rect 5537 4431 5595 4437
rect 8478 4428 8484 4440
rect 8536 4468 8542 4480
rect 10796 4468 10824 4567
rect 11974 4564 11980 4616
rect 12032 4604 12038 4616
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 12032 4576 12173 4604
rect 12032 4564 12038 4576
rect 12161 4573 12173 4576
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 13265 4607 13323 4613
rect 13265 4573 13277 4607
rect 13311 4604 13323 4607
rect 14458 4604 14464 4616
rect 13311 4576 14464 4604
rect 13311 4573 13323 4576
rect 13265 4567 13323 4573
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 15565 4607 15623 4613
rect 15565 4573 15577 4607
rect 15611 4573 15623 4607
rect 15565 4567 15623 4573
rect 13357 4539 13415 4545
rect 13357 4505 13369 4539
rect 13403 4536 13415 4539
rect 13998 4536 14004 4548
rect 13403 4508 14004 4536
rect 13403 4505 13415 4508
rect 13357 4499 13415 4505
rect 13998 4496 14004 4508
rect 14056 4536 14062 4548
rect 14056 4508 14228 4536
rect 14056 4496 14062 4508
rect 8536 4440 10824 4468
rect 11057 4471 11115 4477
rect 8536 4428 8542 4440
rect 11057 4437 11069 4471
rect 11103 4468 11115 4471
rect 11882 4468 11888 4480
rect 11103 4440 11888 4468
rect 11103 4437 11115 4440
rect 11057 4431 11115 4437
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 12066 4468 12072 4480
rect 12027 4440 12072 4468
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 13725 4471 13783 4477
rect 13725 4437 13737 4471
rect 13771 4468 13783 4471
rect 13814 4468 13820 4480
rect 13771 4440 13820 4468
rect 13771 4437 13783 4440
rect 13725 4431 13783 4437
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 14200 4477 14228 4508
rect 14918 4496 14924 4548
rect 14976 4536 14982 4548
rect 15298 4539 15356 4545
rect 15298 4536 15310 4539
rect 14976 4508 15310 4536
rect 14976 4496 14982 4508
rect 15298 4505 15310 4508
rect 15344 4505 15356 4539
rect 15580 4536 15608 4567
rect 15654 4564 15660 4616
rect 15712 4604 15718 4616
rect 16022 4604 16028 4616
rect 15712 4576 16028 4604
rect 15712 4564 15718 4576
rect 16022 4564 16028 4576
rect 16080 4604 16086 4616
rect 16209 4607 16267 4613
rect 16209 4604 16221 4607
rect 16080 4576 16221 4604
rect 16080 4564 16086 4576
rect 16209 4573 16221 4576
rect 16255 4573 16267 4607
rect 16390 4604 16396 4616
rect 16351 4576 16396 4604
rect 16209 4567 16267 4573
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 16945 4607 17003 4613
rect 16945 4604 16957 4607
rect 16632 4576 16957 4604
rect 16632 4564 16638 4576
rect 16945 4573 16957 4576
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 16758 4536 16764 4548
rect 15580 4508 16764 4536
rect 15298 4499 15356 4505
rect 16758 4496 16764 4508
rect 16816 4496 16822 4548
rect 17212 4539 17270 4545
rect 17212 4505 17224 4539
rect 17258 4536 17270 4539
rect 17310 4536 17316 4548
rect 17258 4508 17316 4536
rect 17258 4505 17270 4508
rect 17212 4499 17270 4505
rect 17310 4496 17316 4508
rect 17368 4496 17374 4548
rect 14185 4471 14243 4477
rect 14185 4437 14197 4471
rect 14231 4437 14243 4471
rect 14185 4431 14243 4437
rect 16577 4471 16635 4477
rect 16577 4437 16589 4471
rect 16623 4468 16635 4471
rect 16666 4468 16672 4480
rect 16623 4440 16672 4468
rect 16623 4437 16635 4440
rect 16577 4431 16635 4437
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 18322 4468 18328 4480
rect 18283 4440 18328 4468
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 1104 4378 18860 4400
rect 1104 4326 6880 4378
rect 6932 4326 6944 4378
rect 6996 4326 7008 4378
rect 7060 4326 7072 4378
rect 7124 4326 7136 4378
rect 7188 4326 12811 4378
rect 12863 4326 12875 4378
rect 12927 4326 12939 4378
rect 12991 4326 13003 4378
rect 13055 4326 13067 4378
rect 13119 4326 18860 4378
rect 1104 4304 18860 4326
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1670 4224 1676 4236
rect 1728 4224 1734 4276
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3329 4267 3387 4273
rect 3329 4264 3341 4267
rect 3108 4236 3341 4264
rect 3108 4224 3114 4236
rect 3329 4233 3341 4236
rect 3375 4233 3387 4267
rect 3329 4227 3387 4233
rect 7101 4267 7159 4273
rect 7101 4233 7113 4267
rect 7147 4264 7159 4267
rect 8478 4264 8484 4276
rect 7147 4236 8484 4264
rect 7147 4233 7159 4236
rect 7101 4227 7159 4233
rect 8478 4224 8484 4236
rect 8536 4224 8542 4276
rect 9861 4267 9919 4273
rect 9861 4233 9873 4267
rect 9907 4264 9919 4267
rect 10962 4264 10968 4276
rect 9907 4236 10968 4264
rect 9907 4233 9919 4236
rect 9861 4227 9919 4233
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 12250 4264 12256 4276
rect 12211 4236 12256 4264
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 16853 4267 16911 4273
rect 14108 4236 14964 4264
rect 7282 4156 7288 4208
rect 7340 4196 7346 4208
rect 13998 4196 14004 4208
rect 7340 4168 7788 4196
rect 7340 4156 7346 4168
rect 7760 4140 7788 4168
rect 13648 4168 14004 4196
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4128 1547 4131
rect 1949 4131 2007 4137
rect 1949 4128 1961 4131
rect 1535 4100 1961 4128
rect 1535 4097 1547 4100
rect 1489 4091 1547 4097
rect 1949 4097 1961 4100
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2406 4128 2412 4140
rect 2179 4100 2412 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 4157 4131 4215 4137
rect 3528 4100 4108 4128
rect 1762 4020 1768 4072
rect 1820 4060 1826 4072
rect 2317 4063 2375 4069
rect 2317 4060 2329 4063
rect 1820 4032 2329 4060
rect 1820 4020 1826 4032
rect 2317 4029 2329 4032
rect 2363 4060 2375 4063
rect 2498 4060 2504 4072
rect 2363 4032 2504 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 2774 4060 2780 4072
rect 2731 4032 2780 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 3418 4060 3424 4072
rect 3379 4032 3424 4060
rect 3418 4020 3424 4032
rect 3476 4020 3482 4072
rect 3528 4069 3556 4100
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4029 3571 4063
rect 3513 4023 3571 4029
rect 3602 4020 3608 4072
rect 3660 4060 3666 4072
rect 3973 4063 4031 4069
rect 3973 4060 3985 4063
rect 3660 4032 3985 4060
rect 3660 4020 3666 4032
rect 3973 4029 3985 4032
rect 4019 4029 4031 4063
rect 4080 4060 4108 4100
rect 4157 4097 4169 4131
rect 4203 4128 4215 4131
rect 4246 4128 4252 4140
rect 4203 4100 4252 4128
rect 4203 4097 4215 4100
rect 4157 4091 4215 4097
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4890 4137 4896 4140
rect 4884 4128 4896 4137
rect 4851 4100 4896 4128
rect 4884 4091 4896 4100
rect 4890 4088 4896 4091
rect 4948 4088 4954 4140
rect 5350 4088 5356 4140
rect 5408 4128 5414 4140
rect 7742 4128 7748 4140
rect 5408 4100 7328 4128
rect 7655 4100 7748 4128
rect 5408 4088 5414 4100
rect 4522 4060 4528 4072
rect 4080 4032 4528 4060
rect 3973 4023 4031 4029
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4029 4675 4063
rect 7190 4060 7196 4072
rect 7151 4032 7196 4060
rect 4617 4023 4675 4029
rect 2038 3952 2044 4004
rect 2096 3992 2102 4004
rect 4632 3992 4660 4023
rect 7190 4020 7196 4032
rect 7248 4020 7254 4072
rect 7300 4069 7328 4100
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 8012 4131 8070 4137
rect 8012 4097 8024 4131
rect 8058 4128 8070 4131
rect 8938 4128 8944 4140
rect 8058 4100 8944 4128
rect 8058 4097 8070 4100
rect 8012 4091 8070 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 9582 4128 9588 4140
rect 9447 4100 9588 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 9824 4100 10149 4128
rect 9824 4088 9830 4100
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 2096 3964 4660 3992
rect 2096 3952 2102 3964
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 5997 3995 6055 4001
rect 5997 3992 6009 3995
rect 5684 3964 6009 3992
rect 5684 3952 5690 3964
rect 5997 3961 6009 3964
rect 6043 3992 6055 3995
rect 10226 3992 10232 4004
rect 6043 3964 7328 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 2682 3884 2688 3936
rect 2740 3924 2746 3936
rect 2961 3927 3019 3933
rect 2961 3924 2973 3927
rect 2740 3896 2973 3924
rect 2740 3884 2746 3896
rect 2961 3893 2973 3896
rect 3007 3893 3019 3927
rect 4338 3924 4344 3936
rect 4299 3896 4344 3924
rect 2961 3887 3019 3893
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 6914 3924 6920 3936
rect 6779 3896 6920 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 7300 3924 7328 3964
rect 8680 3964 10232 3992
rect 8680 3924 8708 3964
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 10336 3992 10364 4091
rect 10410 4088 10416 4140
rect 10468 4128 10474 4140
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10468 4100 10517 4128
rect 10468 4088 10474 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10962 4128 10968 4140
rect 10923 4100 10968 4128
rect 10505 4091 10563 4097
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11238 4128 11244 4140
rect 11195 4100 11244 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11624 4100 11713 4128
rect 10597 4063 10655 4069
rect 10597 4029 10609 4063
rect 10643 4060 10655 4063
rect 11514 4060 11520 4072
rect 10643 4032 11520 4060
rect 10643 4029 10655 4032
rect 10597 4023 10655 4029
rect 11514 4020 11520 4032
rect 11572 4020 11578 4072
rect 10778 3992 10784 4004
rect 10336 3964 10784 3992
rect 10778 3952 10784 3964
rect 10836 3992 10842 4004
rect 11624 3992 11652 4100
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11882 4128 11888 4140
rect 11843 4100 11888 4128
rect 11701 4091 11759 4097
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 12437 4131 12495 4137
rect 12437 4097 12449 4131
rect 12483 4128 12495 4131
rect 12618 4128 12624 4140
rect 12483 4100 12624 4128
rect 12483 4097 12495 4100
rect 12437 4091 12495 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13648 4128 13676 4168
rect 13998 4156 14004 4168
rect 14056 4156 14062 4208
rect 13814 4128 13820 4140
rect 13219 4100 13676 4128
rect 13775 4100 13820 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 14108 4128 14136 4236
rect 14936 4196 14964 4236
rect 16853 4233 16865 4267
rect 16899 4264 16911 4267
rect 16942 4264 16948 4276
rect 16899 4236 16948 4264
rect 16899 4233 16911 4236
rect 16853 4227 16911 4233
rect 16942 4224 16948 4236
rect 17000 4224 17006 4276
rect 17310 4264 17316 4276
rect 17271 4236 17316 4264
rect 17310 4224 17316 4236
rect 17368 4224 17374 4276
rect 16022 4196 16028 4208
rect 14936 4168 16028 4196
rect 16022 4156 16028 4168
rect 16080 4156 16086 4208
rect 16298 4196 16304 4208
rect 16259 4168 16304 4196
rect 16298 4156 16304 4168
rect 16356 4156 16362 4208
rect 16500 4168 16804 4196
rect 14274 4128 14280 4140
rect 13924 4100 14136 4128
rect 14235 4100 14280 4128
rect 11974 4060 11980 4072
rect 11935 4032 11980 4060
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 13633 4063 13691 4069
rect 13633 4060 13645 4063
rect 12406 4032 13645 4060
rect 10836 3964 11652 3992
rect 10836 3952 10842 3964
rect 11790 3952 11796 4004
rect 11848 3992 11854 4004
rect 12406 3992 12434 4032
rect 13633 4029 13645 4032
rect 13679 4060 13691 4063
rect 13924 4060 13952 4100
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4097 14795 4131
rect 14737 4091 14795 4097
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4128 16175 4131
rect 16500 4128 16528 4168
rect 16666 4128 16672 4140
rect 16163 4100 16528 4128
rect 16627 4100 16672 4128
rect 16163 4097 16175 4100
rect 16117 4091 16175 4097
rect 13679 4032 13952 4060
rect 14001 4063 14059 4069
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 14001 4029 14013 4063
rect 14047 4060 14059 4063
rect 14752 4060 14780 4091
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 16776 4128 16804 4168
rect 17402 4128 17408 4140
rect 16776 4100 17408 4128
rect 17402 4088 17408 4100
rect 17460 4128 17466 4140
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 17460 4100 17509 4128
rect 17460 4088 17466 4100
rect 17497 4097 17509 4100
rect 17543 4097 17555 4131
rect 17678 4128 17684 4140
rect 17639 4100 17684 4128
rect 17497 4091 17555 4097
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 18049 4131 18107 4137
rect 18049 4097 18061 4131
rect 18095 4128 18107 4131
rect 18322 4128 18328 4140
rect 18095 4100 18328 4128
rect 18095 4097 18107 4100
rect 18049 4091 18107 4097
rect 18322 4088 18328 4100
rect 18380 4088 18386 4140
rect 14047 4032 14780 4060
rect 15841 4063 15899 4069
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 15841 4029 15853 4063
rect 15887 4060 15899 4063
rect 16850 4060 16856 4072
rect 15887 4032 16856 4060
rect 15887 4029 15899 4032
rect 15841 4023 15899 4029
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 17770 4060 17776 4072
rect 17731 4032 17776 4060
rect 17770 4020 17776 4032
rect 17828 4020 17834 4072
rect 12894 3992 12900 4004
rect 11848 3964 12434 3992
rect 12807 3964 12900 3992
rect 11848 3952 11854 3964
rect 12894 3952 12900 3964
rect 12952 3992 12958 4004
rect 15654 3992 15660 4004
rect 12952 3964 15660 3992
rect 12952 3952 12958 3964
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 15933 3995 15991 4001
rect 15933 3961 15945 3995
rect 15979 3992 15991 3995
rect 16114 3992 16120 4004
rect 15979 3964 16120 3992
rect 15979 3961 15991 3964
rect 15933 3955 15991 3961
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 18230 3992 18236 4004
rect 16224 3964 18092 3992
rect 18191 3964 18236 3992
rect 7300 3896 8708 3924
rect 9030 3884 9036 3936
rect 9088 3924 9094 3936
rect 9125 3927 9183 3933
rect 9125 3924 9137 3927
rect 9088 3896 9137 3924
rect 9088 3884 9094 3896
rect 9125 3893 9137 3896
rect 9171 3893 9183 3927
rect 9125 3887 9183 3893
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 9272 3896 9505 3924
rect 9272 3884 9278 3896
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11480 3896 11529 3924
rect 11480 3884 11486 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 13170 3924 13176 3936
rect 12768 3896 13176 3924
rect 12768 3884 12774 3896
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 13357 3927 13415 3933
rect 13357 3893 13369 3927
rect 13403 3924 13415 3927
rect 14366 3924 14372 3936
rect 13403 3896 14372 3924
rect 13403 3893 13415 3896
rect 13357 3887 13415 3893
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 14550 3924 14556 3936
rect 14507 3896 14556 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14918 3924 14924 3936
rect 14879 3896 14924 3924
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 15565 3927 15623 3933
rect 15565 3893 15577 3927
rect 15611 3924 15623 3927
rect 16224 3924 16252 3964
rect 15611 3896 16252 3924
rect 18064 3924 18092 3964
rect 18230 3952 18236 3964
rect 18288 3952 18294 4004
rect 18690 3924 18696 3936
rect 18064 3896 18696 3924
rect 15611 3893 15623 3896
rect 15565 3887 15623 3893
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 1104 3834 18860 3856
rect 1104 3782 3915 3834
rect 3967 3782 3979 3834
rect 4031 3782 4043 3834
rect 4095 3782 4107 3834
rect 4159 3782 4171 3834
rect 4223 3782 9846 3834
rect 9898 3782 9910 3834
rect 9962 3782 9974 3834
rect 10026 3782 10038 3834
rect 10090 3782 10102 3834
rect 10154 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 15904 3834
rect 15956 3782 15968 3834
rect 16020 3782 16032 3834
rect 16084 3782 18860 3834
rect 1104 3760 18860 3782
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 3602 3720 3608 3732
rect 2464 3692 3608 3720
rect 2464 3680 2470 3692
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 4246 3720 4252 3732
rect 3927 3692 4252 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 4893 3723 4951 3729
rect 4893 3689 4905 3723
rect 4939 3720 4951 3723
rect 5074 3720 5080 3732
rect 4939 3692 5080 3720
rect 4939 3689 4951 3692
rect 4893 3683 4951 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 7558 3720 7564 3732
rect 7147 3692 7564 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8938 3720 8944 3732
rect 8899 3692 8944 3720
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 11790 3720 11796 3732
rect 9048 3692 11796 3720
rect 1578 3612 1584 3664
rect 1636 3612 1642 3664
rect 3418 3652 3424 3664
rect 3331 3624 3424 3652
rect 3418 3612 3424 3624
rect 3476 3652 3482 3664
rect 5534 3652 5540 3664
rect 3476 3624 4292 3652
rect 3476 3612 3482 3624
rect 1596 3584 1624 3612
rect 2038 3584 2044 3596
rect 1596 3556 2044 3584
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 2774 3516 2780 3528
rect 1627 3488 2780 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 2774 3476 2780 3488
rect 2832 3516 2838 3528
rect 3234 3516 3240 3528
rect 2832 3488 3240 3516
rect 2832 3476 2838 3488
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 4264 3525 4292 3624
rect 4356 3624 5540 3652
rect 4356 3593 4384 3624
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 5718 3612 5724 3664
rect 5776 3652 5782 3664
rect 6638 3652 6644 3664
rect 5776 3624 6644 3652
rect 5776 3612 5782 3624
rect 6638 3612 6644 3624
rect 6696 3652 6702 3664
rect 9048 3652 9076 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 11974 3720 11980 3732
rect 11935 3692 11980 3720
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 13357 3723 13415 3729
rect 13357 3689 13369 3723
rect 13403 3720 13415 3723
rect 14274 3720 14280 3732
rect 13403 3692 14280 3720
rect 13403 3689 13415 3692
rect 13357 3683 13415 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 16850 3720 16856 3732
rect 14424 3692 16436 3720
rect 16811 3692 16856 3720
rect 14424 3680 14430 3692
rect 6696 3624 9076 3652
rect 6696 3612 6702 3624
rect 12158 3612 12164 3664
rect 12216 3612 12222 3664
rect 13081 3655 13139 3661
rect 13081 3621 13093 3655
rect 13127 3652 13139 3655
rect 13127 3624 16252 3652
rect 13127 3621 13139 3624
rect 13081 3615 13139 3621
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3553 4399 3587
rect 4341 3547 4399 3553
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 4614 3584 4620 3596
rect 4571 3556 4620 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 5442 3584 5448 3596
rect 5403 3556 5448 3584
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 6733 3587 6791 3593
rect 6733 3584 6745 3587
rect 6604 3556 6745 3584
rect 6604 3544 6610 3556
rect 6733 3553 6745 3556
rect 6779 3584 6791 3587
rect 7377 3587 7435 3593
rect 7377 3584 7389 3587
rect 6779 3556 7389 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 7377 3553 7389 3556
rect 7423 3553 7435 3587
rect 7377 3547 7435 3553
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 11701 3587 11759 3593
rect 9180 3556 9352 3584
rect 9180 3544 9186 3556
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 4295 3488 5365 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 6914 3516 6920 3528
rect 6875 3488 6920 3516
rect 5353 3479 5411 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 9214 3516 9220 3528
rect 9175 3488 9220 3516
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9324 3525 9352 3556
rect 11701 3553 11713 3587
rect 11747 3584 11759 3587
rect 12176 3584 12204 3612
rect 11747 3556 12204 3584
rect 11747 3553 11759 3556
rect 11701 3547 11759 3553
rect 13170 3544 13176 3596
rect 13228 3584 13234 3596
rect 14645 3587 14703 3593
rect 14645 3584 14657 3587
rect 13228 3556 14657 3584
rect 13228 3544 13234 3556
rect 14645 3553 14657 3556
rect 14691 3553 14703 3587
rect 14645 3547 14703 3553
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9456 3488 9501 3516
rect 9456 3476 9462 3488
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 9640 3488 9685 3516
rect 9640 3476 9646 3488
rect 11422 3476 11428 3528
rect 11480 3525 11486 3528
rect 11480 3516 11492 3525
rect 12161 3519 12219 3525
rect 11480 3488 11525 3516
rect 11480 3479 11492 3488
rect 12161 3485 12173 3519
rect 12207 3485 12219 3519
rect 12161 3479 12219 3485
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3485 12311 3519
rect 12894 3516 12900 3528
rect 12855 3488 12900 3516
rect 12253 3479 12311 3485
rect 11480 3476 11486 3479
rect 2308 3451 2366 3457
rect 2308 3417 2320 3451
rect 2354 3448 2366 3451
rect 3142 3448 3148 3460
rect 2354 3420 3148 3448
rect 2354 3417 2366 3420
rect 2308 3411 2366 3417
rect 3142 3408 3148 3420
rect 3200 3408 3206 3460
rect 10134 3448 10140 3460
rect 4264 3420 10140 3448
rect 1765 3383 1823 3389
rect 1765 3349 1777 3383
rect 1811 3380 1823 3383
rect 4264 3380 4292 3420
rect 10134 3408 10140 3420
rect 10192 3408 10198 3460
rect 10962 3408 10968 3460
rect 11020 3448 11026 3460
rect 12176 3448 12204 3479
rect 11020 3420 12204 3448
rect 11020 3408 11026 3420
rect 1811 3352 4292 3380
rect 5261 3383 5319 3389
rect 1811 3349 1823 3352
rect 1765 3343 1823 3349
rect 5261 3349 5273 3383
rect 5307 3380 5319 3383
rect 5626 3380 5632 3392
rect 5307 3352 5632 3380
rect 5307 3349 5319 3352
rect 5261 3343 5319 3349
rect 5626 3340 5632 3352
rect 5684 3340 5690 3392
rect 6086 3380 6092 3392
rect 6047 3352 6092 3380
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 10045 3383 10103 3389
rect 10045 3349 10057 3383
rect 10091 3380 10103 3383
rect 10226 3380 10232 3392
rect 10091 3352 10232 3380
rect 10091 3349 10103 3352
rect 10045 3343 10103 3349
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 10321 3383 10379 3389
rect 10321 3349 10333 3383
rect 10367 3380 10379 3383
rect 11054 3380 11060 3392
rect 10367 3352 11060 3380
rect 10367 3349 10379 3352
rect 10321 3343 10379 3349
rect 11054 3340 11060 3352
rect 11112 3380 11118 3392
rect 12268 3380 12296 3479
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13630 3516 13636 3528
rect 13587 3488 13636 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 13446 3448 13452 3460
rect 12492 3420 13452 3448
rect 12492 3408 12498 3420
rect 13446 3408 13452 3420
rect 13504 3448 13510 3460
rect 13556 3448 13584 3479
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 15289 3519 15347 3525
rect 15289 3516 15301 3519
rect 13872 3488 15301 3516
rect 13872 3476 13878 3488
rect 15289 3485 15301 3488
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 16114 3516 16120 3528
rect 15979 3488 16120 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 16224 3525 16252 3624
rect 16408 3525 16436 3692
rect 16850 3680 16856 3692
rect 16908 3680 16914 3732
rect 17770 3720 17776 3732
rect 17731 3692 17776 3720
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 16482 3612 16488 3664
rect 16540 3652 16546 3664
rect 16540 3624 16585 3652
rect 16540 3612 16546 3624
rect 18141 3587 18199 3593
rect 18141 3553 18153 3587
rect 18187 3584 18199 3587
rect 18322 3584 18328 3596
rect 18187 3556 18328 3584
rect 18187 3553 18199 3556
rect 18141 3547 18199 3553
rect 18322 3544 18328 3556
rect 18380 3544 18386 3596
rect 16209 3519 16267 3525
rect 16209 3485 16221 3519
rect 16255 3485 16267 3519
rect 16209 3479 16267 3485
rect 16393 3519 16451 3525
rect 16393 3485 16405 3519
rect 16439 3485 16451 3519
rect 17034 3516 17040 3528
rect 16995 3488 17040 3516
rect 16393 3479 16451 3485
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 17126 3476 17132 3528
rect 17184 3516 17190 3528
rect 17957 3519 18015 3525
rect 17184 3488 17229 3516
rect 17184 3476 17190 3488
rect 17957 3485 17969 3519
rect 18003 3485 18015 3519
rect 17957 3479 18015 3485
rect 13504 3420 13584 3448
rect 13725 3451 13783 3457
rect 13504 3408 13510 3420
rect 13725 3417 13737 3451
rect 13771 3417 13783 3451
rect 13725 3411 13783 3417
rect 11112 3352 12296 3380
rect 13740 3380 13768 3411
rect 13906 3408 13912 3460
rect 13964 3448 13970 3460
rect 14458 3448 14464 3460
rect 13964 3420 14464 3448
rect 13964 3408 13970 3420
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 14553 3451 14611 3457
rect 14553 3417 14565 3451
rect 14599 3448 14611 3451
rect 14642 3448 14648 3460
rect 14599 3420 14648 3448
rect 14599 3417 14611 3420
rect 14553 3411 14611 3417
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 17052 3448 17080 3476
rect 17972 3448 18000 3479
rect 17052 3420 18000 3448
rect 14093 3383 14151 3389
rect 14093 3380 14105 3383
rect 13740 3352 14105 3380
rect 11112 3340 11118 3352
rect 14093 3349 14105 3352
rect 14139 3349 14151 3383
rect 15102 3380 15108 3392
rect 15063 3352 15108 3380
rect 14093 3343 14151 3349
rect 15102 3340 15108 3352
rect 15160 3340 15166 3392
rect 1104 3290 18860 3312
rect 1104 3238 6880 3290
rect 6932 3238 6944 3290
rect 6996 3238 7008 3290
rect 7060 3238 7072 3290
rect 7124 3238 7136 3290
rect 7188 3238 12811 3290
rect 12863 3238 12875 3290
rect 12927 3238 12939 3290
rect 12991 3238 13003 3290
rect 13055 3238 13067 3290
rect 13119 3238 18860 3290
rect 1104 3216 18860 3238
rect 3142 3176 3148 3188
rect 3103 3148 3148 3176
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 5997 3179 6055 3185
rect 5997 3145 6009 3179
rect 6043 3176 6055 3179
rect 6043 3148 8248 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 2038 3068 2044 3120
rect 2096 3108 2102 3120
rect 2096 3080 4016 3108
rect 2096 3068 2102 3080
rect 2498 3040 2504 3052
rect 2459 3012 2504 3040
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 2682 3040 2688 3052
rect 2643 3012 2688 3040
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 3988 3049 4016 3080
rect 4614 3068 4620 3120
rect 4672 3108 4678 3120
rect 7098 3108 7104 3120
rect 4672 3080 7104 3108
rect 4672 3068 4678 3080
rect 7098 3068 7104 3080
rect 7156 3068 7162 3120
rect 7500 3111 7558 3117
rect 7500 3077 7512 3111
rect 7546 3108 7558 3111
rect 7834 3108 7840 3120
rect 7546 3080 7840 3108
rect 7546 3077 7558 3080
rect 7500 3071 7558 3077
rect 7834 3068 7840 3080
rect 7892 3068 7898 3120
rect 4246 3049 4252 3052
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 2915 3012 3341 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3329 3009 3341 3012
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4240 3003 4252 3049
rect 4304 3040 4310 3052
rect 5718 3040 5724 3052
rect 4304 3012 4340 3040
rect 5679 3012 5724 3040
rect 4246 3000 4252 3003
rect 4304 3000 4310 3012
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 6546 3040 6552 3052
rect 5859 3012 6552 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 7742 3040 7748 3052
rect 7703 3012 7748 3040
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 8220 3049 8248 3148
rect 9214 3136 9220 3188
rect 9272 3176 9278 3188
rect 9582 3176 9588 3188
rect 9272 3148 9588 3176
rect 9272 3136 9278 3148
rect 9582 3136 9588 3148
rect 9640 3176 9646 3188
rect 9953 3179 10011 3185
rect 9953 3176 9965 3179
rect 9640 3148 9965 3176
rect 9640 3136 9646 3148
rect 9953 3145 9965 3148
rect 9999 3145 10011 3179
rect 9953 3139 10011 3145
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 13725 3179 13783 3185
rect 13725 3176 13737 3179
rect 10192 3148 13737 3176
rect 10192 3136 10198 3148
rect 13725 3145 13737 3148
rect 13771 3145 13783 3179
rect 13725 3139 13783 3145
rect 13998 3136 14004 3188
rect 14056 3176 14062 3188
rect 14461 3179 14519 3185
rect 14461 3176 14473 3179
rect 14056 3148 14473 3176
rect 14056 3136 14062 3148
rect 14461 3145 14473 3148
rect 14507 3176 14519 3179
rect 15194 3176 15200 3188
rect 14507 3148 15200 3176
rect 14507 3145 14519 3148
rect 14461 3139 14519 3145
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 15436 3148 16129 3176
rect 15436 3136 15442 3148
rect 16117 3145 16129 3148
rect 16163 3145 16175 3179
rect 16117 3139 16175 3145
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 17184 3148 18061 3176
rect 17184 3136 17190 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 9030 3068 9036 3120
rect 9088 3108 9094 3120
rect 9088 3080 9352 3108
rect 9088 3068 9094 3080
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8840 3043 8898 3049
rect 8840 3009 8852 3043
rect 8886 3040 8898 3043
rect 9122 3040 9128 3052
rect 8886 3012 9128 3040
rect 8886 3009 8898 3012
rect 8840 3003 8898 3009
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 9324 3040 9352 3080
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 10321 3111 10379 3117
rect 10321 3108 10333 3111
rect 9456 3080 10333 3108
rect 9456 3068 9462 3080
rect 10321 3077 10333 3080
rect 10367 3077 10379 3111
rect 10965 3111 11023 3117
rect 10965 3108 10977 3111
rect 10321 3071 10379 3077
rect 10428 3080 10977 3108
rect 10428 3049 10456 3080
rect 10965 3077 10977 3080
rect 11011 3108 11023 3111
rect 11011 3080 11284 3108
rect 11011 3077 11023 3080
rect 10965 3071 11023 3077
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 9324 3012 10241 3040
rect 10229 3009 10241 3012
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 10413 3043 10471 3049
rect 10413 3009 10425 3043
rect 10459 3009 10471 3043
rect 11146 3040 11152 3052
rect 11107 3012 11152 3040
rect 10413 3003 10471 3009
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 11256 3040 11284 3080
rect 12158 3068 12164 3120
rect 12216 3108 12222 3120
rect 14274 3108 14280 3120
rect 12216 3080 14280 3108
rect 12216 3068 12222 3080
rect 12434 3040 12440 3052
rect 11256 3012 12440 3040
rect 12434 3000 12440 3012
rect 12492 3000 12498 3052
rect 12710 3040 12716 3052
rect 12768 3049 12774 3052
rect 13004 3049 13032 3080
rect 14274 3068 14280 3080
rect 14332 3108 14338 3120
rect 15004 3111 15062 3117
rect 14332 3080 14780 3108
rect 14332 3068 14338 3080
rect 12680 3012 12716 3040
rect 12710 3000 12716 3012
rect 12768 3003 12780 3049
rect 12989 3043 13047 3049
rect 12989 3009 13001 3043
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 12768 3000 12774 3003
rect 13630 3000 13636 3052
rect 13688 3040 13694 3052
rect 14752 3049 14780 3080
rect 15004 3077 15016 3111
rect 15050 3108 15062 3111
rect 15102 3108 15108 3120
rect 15050 3080 15108 3108
rect 15050 3077 15062 3080
rect 15004 3071 15062 3077
rect 15102 3068 15108 3080
rect 15160 3068 15166 3120
rect 16298 3068 16304 3120
rect 16356 3108 16362 3120
rect 16914 3111 16972 3117
rect 16914 3108 16926 3111
rect 16356 3080 16926 3108
rect 16356 3068 16362 3080
rect 16914 3077 16926 3080
rect 16960 3077 16972 3111
rect 16914 3071 16972 3077
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13688 3012 13829 3040
rect 13688 3000 13694 3012
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3040 14795 3043
rect 16574 3040 16580 3052
rect 14783 3012 16580 3040
rect 14783 3009 14795 3012
rect 14737 3003 14795 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3040 16727 3043
rect 16758 3040 16764 3052
rect 16715 3012 16764 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 16758 3000 16764 3012
rect 16816 3000 16822 3052
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 2038 2972 2044 2984
rect 1995 2944 2044 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2222 2972 2228 2984
rect 2183 2944 2228 2972
rect 2222 2932 2228 2944
rect 2280 2932 2286 2984
rect 7760 2972 7788 3000
rect 8573 2975 8631 2981
rect 8573 2972 8585 2975
rect 7760 2944 8585 2972
rect 8573 2941 8585 2944
rect 8619 2941 8631 2975
rect 8573 2935 8631 2941
rect 13170 2932 13176 2984
rect 13228 2972 13234 2984
rect 13909 2975 13967 2981
rect 13909 2972 13921 2975
rect 13228 2944 13921 2972
rect 13228 2932 13234 2944
rect 13909 2941 13921 2944
rect 13955 2941 13967 2975
rect 13909 2935 13967 2941
rect 2240 2904 2268 2932
rect 3605 2907 3663 2913
rect 3605 2904 3617 2907
rect 2240 2876 3617 2904
rect 3605 2873 3617 2876
rect 3651 2873 3663 2907
rect 3605 2867 3663 2873
rect 5353 2907 5411 2913
rect 5353 2873 5365 2907
rect 5399 2904 5411 2907
rect 5534 2904 5540 2916
rect 5399 2876 5540 2904
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 5534 2864 5540 2876
rect 5592 2904 5598 2916
rect 6730 2904 6736 2916
rect 5592 2876 6736 2904
rect 5592 2864 5598 2876
rect 6730 2864 6736 2876
rect 6788 2864 6794 2916
rect 7834 2864 7840 2916
rect 7892 2904 7898 2916
rect 8021 2907 8079 2913
rect 8021 2904 8033 2907
rect 7892 2876 8033 2904
rect 7892 2864 7898 2876
rect 8021 2873 8033 2876
rect 8067 2873 8079 2907
rect 8021 2867 8079 2873
rect 10781 2907 10839 2913
rect 10781 2873 10793 2907
rect 10827 2904 10839 2907
rect 10827 2876 11744 2904
rect 10827 2873 10839 2876
rect 10781 2867 10839 2873
rect 6365 2839 6423 2845
rect 6365 2805 6377 2839
rect 6411 2836 6423 2839
rect 7374 2836 7380 2848
rect 6411 2808 7380 2836
rect 6411 2805 6423 2808
rect 6365 2799 6423 2805
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 11606 2836 11612 2848
rect 11567 2808 11612 2836
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 11716 2836 11744 2876
rect 12618 2836 12624 2848
rect 11716 2808 12624 2836
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 13354 2836 13360 2848
rect 13315 2808 13360 2836
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 1104 2746 18860 2768
rect 1104 2694 3915 2746
rect 3967 2694 3979 2746
rect 4031 2694 4043 2746
rect 4095 2694 4107 2746
rect 4159 2694 4171 2746
rect 4223 2694 9846 2746
rect 9898 2694 9910 2746
rect 9962 2694 9974 2746
rect 10026 2694 10038 2746
rect 10090 2694 10102 2746
rect 10154 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 15904 2746
rect 15956 2694 15968 2746
rect 16020 2694 16032 2746
rect 16084 2694 18860 2746
rect 1104 2672 18860 2694
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 9306 2632 9312 2644
rect 3476 2604 9312 2632
rect 3476 2592 3482 2604
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 11204 2604 11621 2632
rect 11204 2592 11210 2604
rect 11609 2601 11621 2604
rect 11655 2601 11667 2635
rect 11609 2595 11667 2601
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 12805 2635 12863 2641
rect 12805 2632 12817 2635
rect 12768 2604 12817 2632
rect 12768 2592 12774 2604
rect 12805 2601 12817 2604
rect 12851 2601 12863 2635
rect 12805 2595 12863 2601
rect 13725 2635 13783 2641
rect 13725 2601 13737 2635
rect 13771 2632 13783 2635
rect 13814 2632 13820 2644
rect 13771 2604 13820 2632
rect 13771 2601 13783 2604
rect 13725 2595 13783 2601
rect 13814 2592 13820 2604
rect 13872 2592 13878 2644
rect 14642 2592 14648 2644
rect 14700 2632 14706 2644
rect 15657 2635 15715 2641
rect 15657 2632 15669 2635
rect 14700 2604 15669 2632
rect 14700 2592 14706 2604
rect 15657 2601 15669 2604
rect 15703 2601 15715 2635
rect 15657 2595 15715 2601
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2564 4215 2567
rect 4246 2564 4252 2576
rect 4203 2536 4252 2564
rect 4203 2533 4215 2536
rect 4157 2527 4215 2533
rect 4246 2524 4252 2536
rect 4304 2524 4310 2576
rect 6546 2564 6552 2576
rect 6507 2536 6552 2564
rect 6546 2524 6552 2536
rect 6604 2524 6610 2576
rect 8846 2564 8852 2576
rect 6886 2536 8852 2564
rect 1302 2456 1308 2508
rect 1360 2496 1366 2508
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 1360 2468 2237 2496
rect 1360 2456 1366 2468
rect 2225 2465 2237 2468
rect 2271 2496 2283 2499
rect 2314 2496 2320 2508
rect 2271 2468 2320 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 2314 2456 2320 2468
rect 2372 2456 2378 2508
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6886 2496 6914 2536
rect 8846 2524 8852 2536
rect 8904 2524 8910 2576
rect 9122 2564 9128 2576
rect 9083 2536 9128 2564
rect 9122 2524 9128 2536
rect 9180 2524 9186 2576
rect 10137 2567 10195 2573
rect 10137 2533 10149 2567
rect 10183 2533 10195 2567
rect 10137 2527 10195 2533
rect 10597 2567 10655 2573
rect 10597 2533 10609 2567
rect 10643 2564 10655 2567
rect 11698 2564 11704 2576
rect 10643 2536 11704 2564
rect 10643 2533 10655 2536
rect 10597 2527 10655 2533
rect 7098 2496 7104 2508
rect 5767 2468 6914 2496
rect 7059 2468 7104 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 9582 2496 9588 2508
rect 9543 2468 9588 2496
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 10152 2496 10180 2527
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 13170 2564 13176 2576
rect 12268 2536 13176 2564
rect 10152 2468 11560 2496
rect 1946 2428 1952 2440
rect 1907 2400 1952 2428
rect 1946 2388 1952 2400
rect 2004 2388 2010 2440
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 2774 2428 2780 2440
rect 2547 2400 2780 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 3878 2428 3884 2440
rect 3467 2400 3884 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4338 2428 4344 2440
rect 4019 2400 4344 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 4908 2360 4936 2391
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 5592 2400 6009 2428
rect 5592 2388 5598 2400
rect 5997 2397 6009 2400
rect 6043 2428 6055 2431
rect 6086 2428 6092 2440
rect 6043 2400 6092 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6086 2388 6092 2400
rect 6144 2388 6150 2440
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6788 2400 6929 2428
rect 6788 2388 6794 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 7282 2428 7288 2440
rect 7055 2400 7288 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2428 8171 2431
rect 9030 2428 9036 2440
rect 8159 2400 9036 2428
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 9030 2388 9036 2400
rect 9088 2388 9094 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9398 2428 9404 2440
rect 9355 2400 9404 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 9490 2388 9496 2440
rect 9548 2428 9554 2440
rect 9953 2431 10011 2437
rect 9548 2400 9593 2428
rect 9548 2388 9554 2400
rect 9953 2397 9965 2431
rect 9999 2428 10011 2431
rect 10318 2428 10324 2440
rect 9999 2400 10324 2428
rect 9999 2397 10011 2400
rect 9953 2391 10011 2397
rect 6454 2360 6460 2372
rect 4908 2332 6460 2360
rect 6454 2320 6460 2332
rect 6512 2320 6518 2372
rect 8573 2363 8631 2369
rect 8573 2329 8585 2363
rect 8619 2360 8631 2363
rect 9968 2360 9996 2391
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 8619 2332 9996 2360
rect 8619 2329 8631 2332
rect 8573 2323 8631 2329
rect 10226 2320 10232 2372
rect 10284 2360 10290 2372
rect 10428 2360 10456 2391
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11532 2428 11560 2468
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 12268 2505 12296 2536
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 15470 2524 15476 2576
rect 15528 2564 15534 2576
rect 16025 2567 16083 2573
rect 16025 2564 16037 2567
rect 15528 2536 16037 2564
rect 15528 2524 15534 2536
rect 16025 2533 16037 2536
rect 16071 2533 16083 2567
rect 16025 2527 16083 2533
rect 12069 2499 12127 2505
rect 12069 2496 12081 2499
rect 11664 2468 12081 2496
rect 11664 2456 11670 2468
rect 12069 2465 12081 2468
rect 12115 2465 12127 2499
rect 12069 2459 12127 2465
rect 12253 2499 12311 2505
rect 12253 2465 12265 2499
rect 12299 2465 12311 2499
rect 13906 2496 13912 2508
rect 12253 2459 12311 2465
rect 12452 2468 13912 2496
rect 12452 2428 12480 2468
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 14274 2496 14280 2508
rect 14235 2468 14280 2496
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 12618 2428 12624 2440
rect 11204 2400 11249 2428
rect 11532 2400 12480 2428
rect 12579 2400 12624 2428
rect 11204 2388 11210 2400
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 13354 2428 13360 2440
rect 13315 2400 13360 2428
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13446 2388 13452 2440
rect 13504 2428 13510 2440
rect 14550 2437 14556 2440
rect 13541 2431 13599 2437
rect 13541 2428 13553 2431
rect 13504 2400 13553 2428
rect 13504 2388 13510 2400
rect 13541 2397 13553 2400
rect 13587 2397 13599 2431
rect 14544 2428 14556 2437
rect 14511 2400 14556 2428
rect 13541 2391 13599 2397
rect 14544 2391 14556 2400
rect 14550 2388 14556 2391
rect 14608 2388 14614 2440
rect 16206 2428 16212 2440
rect 16167 2400 16212 2428
rect 16206 2388 16212 2400
rect 16264 2388 16270 2440
rect 17126 2428 17132 2440
rect 17087 2400 17132 2428
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 17678 2388 17684 2440
rect 17736 2428 17742 2440
rect 17773 2431 17831 2437
rect 17773 2428 17785 2431
rect 17736 2400 17785 2428
rect 17736 2388 17742 2400
rect 17773 2397 17785 2400
rect 17819 2397 17831 2431
rect 17773 2391 17831 2397
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 12710 2360 12716 2372
rect 10284 2332 12716 2360
rect 10284 2320 10290 2332
rect 12710 2320 12716 2332
rect 12768 2320 12774 2372
rect 13722 2320 13728 2372
rect 13780 2360 13786 2372
rect 18064 2360 18092 2391
rect 13780 2332 18092 2360
rect 13780 2320 13786 2332
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 7650 2292 7656 2304
rect 2096 2264 7656 2292
rect 2096 2252 2102 2264
rect 7650 2252 7656 2264
rect 7708 2252 7714 2304
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 7800 2264 7941 2292
rect 7800 2252 7806 2264
rect 7929 2261 7941 2264
rect 7975 2261 7987 2295
rect 7929 2255 7987 2261
rect 10965 2295 11023 2301
rect 10965 2261 10977 2295
rect 11011 2292 11023 2295
rect 11514 2292 11520 2304
rect 11011 2264 11520 2292
rect 11011 2261 11023 2264
rect 10965 2255 11023 2261
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 11974 2292 11980 2304
rect 11935 2264 11980 2292
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 16945 2295 17003 2301
rect 16945 2292 16957 2295
rect 16816 2264 16957 2292
rect 16816 2252 16822 2264
rect 16945 2261 16957 2264
rect 16991 2261 17003 2295
rect 16945 2255 17003 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18233 2295 18291 2301
rect 18233 2292 18245 2295
rect 18104 2264 18245 2292
rect 18104 2252 18110 2264
rect 18233 2261 18245 2264
rect 18279 2261 18291 2295
rect 18233 2255 18291 2261
rect 1104 2202 18860 2224
rect 1104 2150 6880 2202
rect 6932 2150 6944 2202
rect 6996 2150 7008 2202
rect 7060 2150 7072 2202
rect 7124 2150 7136 2202
rect 7188 2150 12811 2202
rect 12863 2150 12875 2202
rect 12927 2150 12939 2202
rect 12991 2150 13003 2202
rect 13055 2150 13067 2202
rect 13119 2150 18860 2202
rect 1104 2128 18860 2150
rect 1946 2048 1952 2100
rect 2004 2088 2010 2100
rect 7466 2088 7472 2100
rect 2004 2060 7472 2088
rect 2004 2048 2010 2060
rect 7466 2048 7472 2060
rect 7524 2048 7530 2100
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 11974 2088 11980 2100
rect 7708 2060 11980 2088
rect 7708 2048 7714 2060
rect 11974 2048 11980 2060
rect 12032 2048 12038 2100
rect 9490 1980 9496 2032
rect 9548 2020 9554 2032
rect 14182 2020 14188 2032
rect 9548 1992 14188 2020
rect 9548 1980 9554 1992
rect 14182 1980 14188 1992
rect 14240 1980 14246 2032
<< via1 >>
rect 6880 17382 6932 17434
rect 6944 17382 6996 17434
rect 7008 17382 7060 17434
rect 7072 17382 7124 17434
rect 7136 17382 7188 17434
rect 12811 17382 12863 17434
rect 12875 17382 12927 17434
rect 12939 17382 12991 17434
rect 13003 17382 13055 17434
rect 13067 17382 13119 17434
rect 4344 17280 4396 17332
rect 7748 17280 7800 17332
rect 9680 17280 9732 17332
rect 14188 17280 14240 17332
rect 18052 17280 18104 17332
rect 1308 17144 1360 17196
rect 2872 17144 2924 17196
rect 6552 17144 6604 17196
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 6736 17144 6788 17153
rect 6644 17076 6696 17128
rect 7288 17144 7340 17196
rect 12440 17212 12492 17264
rect 7932 17008 7984 17060
rect 2964 16983 3016 16992
rect 2964 16949 2973 16983
rect 2973 16949 3007 16983
rect 3007 16949 3016 16983
rect 2964 16940 3016 16949
rect 7196 16983 7248 16992
rect 7196 16949 7205 16983
rect 7205 16949 7239 16983
rect 7239 16949 7248 16983
rect 7196 16940 7248 16949
rect 9036 17144 9088 17196
rect 10416 17144 10468 17196
rect 11612 17144 11664 17196
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 15016 17187 15068 17196
rect 9496 17076 9548 17128
rect 10324 17076 10376 17128
rect 12624 17076 12676 17128
rect 11060 17008 11112 17060
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 16764 17144 16816 17196
rect 17040 17144 17092 17196
rect 17592 17144 17644 17196
rect 18052 17187 18104 17196
rect 18052 17153 18061 17187
rect 18061 17153 18095 17187
rect 18095 17153 18104 17187
rect 18052 17144 18104 17153
rect 16304 17119 16356 17128
rect 16304 17085 16313 17119
rect 16313 17085 16347 17119
rect 16347 17085 16356 17119
rect 16304 17076 16356 17085
rect 15384 17008 15436 17060
rect 17224 17008 17276 17060
rect 17684 17051 17736 17060
rect 17684 17017 17693 17051
rect 17693 17017 17727 17051
rect 17727 17017 17736 17051
rect 17684 17008 17736 17017
rect 10600 16940 10652 16992
rect 11888 16940 11940 16992
rect 14832 16983 14884 16992
rect 14832 16949 14841 16983
rect 14841 16949 14875 16983
rect 14875 16949 14884 16983
rect 14832 16940 14884 16949
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 3915 16838 3967 16890
rect 3979 16838 4031 16890
rect 4043 16838 4095 16890
rect 4107 16838 4159 16890
rect 4171 16838 4223 16890
rect 9846 16838 9898 16890
rect 9910 16838 9962 16890
rect 9974 16838 10026 16890
rect 10038 16838 10090 16890
rect 10102 16838 10154 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 15904 16838 15956 16890
rect 15968 16838 16020 16890
rect 16032 16838 16084 16890
rect 2872 16736 2924 16788
rect 6736 16736 6788 16788
rect 2504 16668 2556 16720
rect 3148 16711 3200 16720
rect 3148 16677 3157 16711
rect 3157 16677 3191 16711
rect 3191 16677 3200 16711
rect 3148 16668 3200 16677
rect 2412 16643 2464 16652
rect 2412 16609 2421 16643
rect 2421 16609 2455 16643
rect 2455 16609 2464 16643
rect 2412 16600 2464 16609
rect 9036 16736 9088 16788
rect 7748 16668 7800 16720
rect 11612 16711 11664 16720
rect 11612 16677 11621 16711
rect 11621 16677 11655 16711
rect 11655 16677 11664 16711
rect 11612 16668 11664 16677
rect 9128 16643 9180 16652
rect 9128 16609 9137 16643
rect 9137 16609 9171 16643
rect 9171 16609 9180 16643
rect 9128 16600 9180 16609
rect 10324 16600 10376 16652
rect 10968 16600 11020 16652
rect 12256 16600 12308 16652
rect 16580 16643 16632 16652
rect 16580 16609 16589 16643
rect 16589 16609 16623 16643
rect 16623 16609 16632 16643
rect 16580 16600 16632 16609
rect 20 16532 72 16584
rect 2964 16532 3016 16584
rect 4344 16532 4396 16584
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 5172 16532 5224 16541
rect 6368 16532 6420 16584
rect 7564 16532 7616 16584
rect 2228 16507 2280 16516
rect 2228 16473 2237 16507
rect 2237 16473 2271 16507
rect 2271 16473 2280 16507
rect 2228 16464 2280 16473
rect 3332 16464 3384 16516
rect 7472 16464 7524 16516
rect 1952 16396 2004 16448
rect 2780 16396 2832 16448
rect 3792 16439 3844 16448
rect 3792 16405 3801 16439
rect 3801 16405 3835 16439
rect 3835 16405 3844 16439
rect 3792 16396 3844 16405
rect 5540 16396 5592 16448
rect 6644 16396 6696 16448
rect 7932 16575 7984 16584
rect 7932 16541 7941 16575
rect 7941 16541 7975 16575
rect 7975 16541 7984 16575
rect 7932 16532 7984 16541
rect 10232 16532 10284 16584
rect 11704 16532 11756 16584
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 12440 16532 12492 16584
rect 14832 16532 14884 16584
rect 16672 16532 16724 16584
rect 9404 16507 9456 16516
rect 9404 16473 9438 16507
rect 9438 16473 9456 16507
rect 9404 16464 9456 16473
rect 11244 16396 11296 16448
rect 15936 16507 15988 16516
rect 15936 16473 15945 16507
rect 15945 16473 15979 16507
rect 15979 16473 15988 16507
rect 15936 16464 15988 16473
rect 16120 16507 16172 16516
rect 16120 16473 16129 16507
rect 16129 16473 16163 16507
rect 16163 16473 16172 16507
rect 16120 16464 16172 16473
rect 12164 16396 12216 16448
rect 13452 16396 13504 16448
rect 13728 16439 13780 16448
rect 13728 16405 13737 16439
rect 13737 16405 13771 16439
rect 13771 16405 13780 16439
rect 13728 16396 13780 16405
rect 15476 16396 15528 16448
rect 16856 16396 16908 16448
rect 17500 16396 17552 16448
rect 6880 16294 6932 16346
rect 6944 16294 6996 16346
rect 7008 16294 7060 16346
rect 7072 16294 7124 16346
rect 7136 16294 7188 16346
rect 12811 16294 12863 16346
rect 12875 16294 12927 16346
rect 12939 16294 12991 16346
rect 13003 16294 13055 16346
rect 13067 16294 13119 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 2228 16235 2280 16244
rect 2228 16201 2237 16235
rect 2237 16201 2271 16235
rect 2271 16201 2280 16235
rect 2228 16192 2280 16201
rect 3516 16235 3568 16244
rect 3516 16201 3525 16235
rect 3525 16201 3559 16235
rect 3559 16201 3568 16235
rect 3516 16192 3568 16201
rect 3700 16235 3752 16244
rect 3700 16201 3709 16235
rect 3709 16201 3743 16235
rect 3743 16201 3752 16235
rect 3700 16192 3752 16201
rect 5632 16192 5684 16244
rect 6368 16235 6420 16244
rect 6368 16201 6377 16235
rect 6377 16201 6411 16235
rect 6411 16201 6420 16235
rect 6368 16192 6420 16201
rect 9404 16235 9456 16244
rect 9404 16201 9413 16235
rect 9413 16201 9447 16235
rect 9447 16201 9456 16235
rect 9404 16192 9456 16201
rect 10232 16235 10284 16244
rect 10232 16201 10241 16235
rect 10241 16201 10275 16235
rect 10275 16201 10284 16235
rect 10232 16192 10284 16201
rect 3608 16167 3660 16176
rect 3608 16133 3617 16167
rect 3617 16133 3651 16167
rect 3651 16133 3660 16167
rect 3608 16124 3660 16133
rect 6552 16167 6604 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 2780 16099 2832 16108
rect 2780 16065 2789 16099
rect 2789 16065 2823 16099
rect 2823 16065 2832 16099
rect 2780 16056 2832 16065
rect 1768 15920 1820 15972
rect 3332 16056 3384 16108
rect 4252 16056 4304 16108
rect 5632 16099 5684 16108
rect 5632 16065 5641 16099
rect 5641 16065 5675 16099
rect 5675 16065 5684 16099
rect 6552 16133 6561 16167
rect 6561 16133 6595 16167
rect 6595 16133 6604 16167
rect 6552 16124 6604 16133
rect 6736 16124 6788 16176
rect 12532 16192 12584 16244
rect 5632 16056 5684 16065
rect 6644 16056 6696 16108
rect 7196 16099 7248 16108
rect 7196 16065 7205 16099
rect 7205 16065 7239 16099
rect 7239 16065 7248 16099
rect 7196 16056 7248 16065
rect 7564 16056 7616 16108
rect 8024 16099 8076 16108
rect 8024 16065 8058 16099
rect 8058 16065 8076 16099
rect 8024 16056 8076 16065
rect 3516 15988 3568 16040
rect 3792 15988 3844 16040
rect 3424 15920 3476 15972
rect 5264 15852 5316 15904
rect 5448 16031 5500 16040
rect 5448 15997 5457 16031
rect 5457 15997 5491 16031
rect 5491 15997 5500 16031
rect 5448 15988 5500 15997
rect 9220 15920 9272 15972
rect 10324 16099 10376 16108
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 12716 16124 12768 16176
rect 13452 16192 13504 16244
rect 15016 16192 15068 16244
rect 15292 16192 15344 16244
rect 15200 16124 15252 16176
rect 15476 16167 15528 16176
rect 15476 16133 15485 16167
rect 15485 16133 15519 16167
rect 15519 16133 15528 16167
rect 15476 16124 15528 16133
rect 15936 16192 15988 16244
rect 17040 16235 17092 16244
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 16672 16167 16724 16176
rect 10876 16056 10928 16108
rect 13268 16056 13320 16108
rect 13728 16056 13780 16108
rect 16212 16056 16264 16108
rect 16672 16133 16681 16167
rect 16681 16133 16715 16167
rect 16715 16133 16724 16167
rect 16672 16124 16724 16133
rect 17500 16099 17552 16108
rect 17500 16065 17509 16099
rect 17509 16065 17543 16099
rect 17543 16065 17552 16099
rect 17500 16056 17552 16065
rect 11704 15988 11756 16040
rect 12072 15988 12124 16040
rect 7288 15852 7340 15904
rect 7932 15852 7984 15904
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 12624 15963 12676 15972
rect 12624 15929 12633 15963
rect 12633 15929 12667 15963
rect 12667 15929 12676 15963
rect 12624 15920 12676 15929
rect 11980 15852 12032 15904
rect 12348 15852 12400 15904
rect 12992 15895 13044 15904
rect 12992 15861 13001 15895
rect 13001 15861 13035 15895
rect 13035 15861 13044 15895
rect 12992 15852 13044 15861
rect 13544 15852 13596 15904
rect 17408 15988 17460 16040
rect 14004 15852 14056 15904
rect 15660 15895 15712 15904
rect 15660 15861 15669 15895
rect 15669 15861 15703 15895
rect 15703 15861 15712 15895
rect 15660 15852 15712 15861
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 3915 15750 3967 15802
rect 3979 15750 4031 15802
rect 4043 15750 4095 15802
rect 4107 15750 4159 15802
rect 4171 15750 4223 15802
rect 9846 15750 9898 15802
rect 9910 15750 9962 15802
rect 9974 15750 10026 15802
rect 10038 15750 10090 15802
rect 10102 15750 10154 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 15904 15750 15956 15802
rect 15968 15750 16020 15802
rect 16032 15750 16084 15802
rect 2780 15648 2832 15700
rect 3332 15691 3384 15700
rect 3332 15657 3341 15691
rect 3341 15657 3375 15691
rect 3375 15657 3384 15691
rect 3332 15648 3384 15657
rect 3608 15648 3660 15700
rect 5264 15648 5316 15700
rect 7196 15648 7248 15700
rect 10876 15691 10928 15700
rect 10876 15657 10885 15691
rect 10885 15657 10919 15691
rect 10919 15657 10928 15691
rect 10876 15648 10928 15657
rect 12624 15648 12676 15700
rect 15200 15691 15252 15700
rect 15200 15657 15209 15691
rect 15209 15657 15243 15691
rect 15243 15657 15252 15691
rect 15200 15648 15252 15657
rect 16212 15648 16264 15700
rect 7840 15580 7892 15632
rect 3148 15555 3200 15564
rect 3148 15521 3157 15555
rect 3157 15521 3191 15555
rect 3191 15521 3200 15555
rect 3148 15512 3200 15521
rect 3792 15555 3844 15564
rect 3792 15521 3801 15555
rect 3801 15521 3835 15555
rect 3835 15521 3844 15555
rect 3792 15512 3844 15521
rect 1768 15419 1820 15428
rect 1768 15385 1802 15419
rect 1802 15385 1820 15419
rect 1768 15376 1820 15385
rect 1860 15376 1912 15428
rect 3424 15487 3476 15496
rect 3424 15453 3433 15487
rect 3433 15453 3467 15487
rect 3467 15453 3476 15487
rect 5172 15512 5224 15564
rect 8300 15580 8352 15632
rect 11244 15623 11296 15632
rect 11244 15589 11253 15623
rect 11253 15589 11287 15623
rect 11287 15589 11296 15623
rect 11244 15580 11296 15589
rect 3424 15444 3476 15453
rect 4344 15444 4396 15496
rect 5356 15444 5408 15496
rect 5540 15487 5592 15496
rect 5540 15453 5574 15487
rect 5574 15453 5592 15487
rect 5540 15444 5592 15453
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 8484 15512 8536 15564
rect 8300 15444 8352 15496
rect 9588 15444 9640 15496
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 11336 15512 11388 15564
rect 12992 15580 13044 15632
rect 16672 15580 16724 15632
rect 15292 15512 15344 15564
rect 9772 15444 9824 15453
rect 4068 15376 4120 15428
rect 7932 15419 7984 15428
rect 7932 15385 7941 15419
rect 7941 15385 7975 15419
rect 7975 15385 7984 15419
rect 7932 15376 7984 15385
rect 8668 15376 8720 15428
rect 11152 15444 11204 15496
rect 12072 15487 12124 15496
rect 12072 15453 12081 15487
rect 12081 15453 12115 15487
rect 12115 15453 12124 15487
rect 12072 15444 12124 15453
rect 12532 15444 12584 15496
rect 7472 15308 7524 15360
rect 8208 15351 8260 15360
rect 8208 15317 8217 15351
rect 8217 15317 8251 15351
rect 8251 15317 8260 15351
rect 8208 15308 8260 15317
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 11704 15308 11756 15360
rect 11980 15351 12032 15360
rect 11980 15317 11989 15351
rect 11989 15317 12023 15351
rect 12023 15317 12032 15351
rect 13176 15419 13228 15428
rect 13176 15385 13185 15419
rect 13185 15385 13219 15419
rect 13219 15385 13228 15419
rect 13176 15376 13228 15385
rect 13544 15444 13596 15496
rect 14004 15444 14056 15496
rect 15476 15444 15528 15496
rect 16580 15512 16632 15564
rect 16028 15444 16080 15496
rect 15200 15376 15252 15428
rect 16304 15419 16356 15428
rect 16304 15385 16313 15419
rect 16313 15385 16347 15419
rect 16347 15385 16356 15419
rect 16304 15376 16356 15385
rect 17316 15376 17368 15428
rect 11980 15308 12032 15317
rect 12624 15351 12676 15360
rect 12624 15317 12633 15351
rect 12633 15317 12667 15351
rect 12667 15317 12676 15351
rect 12624 15308 12676 15317
rect 13268 15308 13320 15360
rect 13452 15351 13504 15360
rect 13452 15317 13461 15351
rect 13461 15317 13495 15351
rect 13495 15317 13504 15351
rect 13452 15308 13504 15317
rect 15660 15308 15712 15360
rect 16856 15308 16908 15360
rect 6880 15206 6932 15258
rect 6944 15206 6996 15258
rect 7008 15206 7060 15258
rect 7072 15206 7124 15258
rect 7136 15206 7188 15258
rect 12811 15206 12863 15258
rect 12875 15206 12927 15258
rect 12939 15206 12991 15258
rect 13003 15206 13055 15258
rect 13067 15206 13119 15258
rect 3792 15104 3844 15156
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 8024 15104 8076 15156
rect 11980 15104 12032 15156
rect 12716 15147 12768 15156
rect 12716 15113 12725 15147
rect 12725 15113 12759 15147
rect 12759 15113 12768 15147
rect 12716 15104 12768 15113
rect 13176 15104 13228 15156
rect 5632 15036 5684 15088
rect 1860 14943 1912 14952
rect 1860 14909 1869 14943
rect 1869 14909 1903 14943
rect 1903 14909 1912 14943
rect 1860 14900 1912 14909
rect 3700 14943 3752 14952
rect 3700 14909 3709 14943
rect 3709 14909 3743 14943
rect 3743 14909 3752 14943
rect 3700 14900 3752 14909
rect 4068 14900 4120 14952
rect 3884 14832 3936 14884
rect 4896 14807 4948 14816
rect 4896 14773 4905 14807
rect 4905 14773 4939 14807
rect 4939 14773 4948 14807
rect 4896 14764 4948 14773
rect 5264 14900 5316 14952
rect 5540 14943 5592 14952
rect 5540 14909 5549 14943
rect 5549 14909 5583 14943
rect 5583 14909 5592 14943
rect 5540 14900 5592 14909
rect 6276 14900 6328 14952
rect 7288 14968 7340 15020
rect 7012 14900 7064 14952
rect 7472 14968 7524 15020
rect 7840 15011 7892 15020
rect 7840 14977 7849 15011
rect 7849 14977 7883 15011
rect 7883 14977 7892 15011
rect 7840 14968 7892 14977
rect 8208 14968 8260 15020
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 8668 15011 8720 15020
rect 8668 14977 8677 15011
rect 8677 14977 8711 15011
rect 8711 14977 8720 15011
rect 8668 14968 8720 14977
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 9312 14900 9364 14952
rect 12348 15079 12400 15088
rect 12348 15045 12357 15079
rect 12357 15045 12391 15079
rect 12391 15045 12400 15079
rect 12348 15036 12400 15045
rect 12532 15079 12584 15088
rect 12532 15045 12541 15079
rect 12541 15045 12575 15079
rect 12575 15045 12584 15079
rect 13452 15079 13504 15088
rect 12532 15036 12584 15045
rect 13452 15045 13486 15079
rect 13486 15045 13504 15079
rect 13452 15036 13504 15045
rect 15200 15104 15252 15156
rect 17316 15147 17368 15156
rect 16120 15036 16172 15088
rect 16672 15079 16724 15088
rect 16672 15045 16681 15079
rect 16681 15045 16715 15079
rect 16715 15045 16724 15079
rect 16672 15036 16724 15045
rect 16764 15036 16816 15088
rect 9588 14968 9640 15020
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 10232 14968 10284 15020
rect 10876 15011 10928 15020
rect 10876 14977 10885 15011
rect 10885 14977 10919 15011
rect 10919 14977 10928 15011
rect 12072 15011 12124 15020
rect 10876 14968 10928 14977
rect 12072 14977 12081 15011
rect 12081 14977 12115 15011
rect 12115 14977 12124 15011
rect 12072 14968 12124 14977
rect 15476 14968 15528 15020
rect 16304 14968 16356 15020
rect 17316 15113 17325 15147
rect 17325 15113 17359 15147
rect 17359 15113 17368 15147
rect 17316 15104 17368 15113
rect 18328 15011 18380 15020
rect 18328 14977 18337 15011
rect 18337 14977 18371 15011
rect 18371 14977 18380 15011
rect 18328 14968 18380 14977
rect 12440 14900 12492 14952
rect 12716 14900 12768 14952
rect 11336 14832 11388 14884
rect 6552 14764 6604 14816
rect 6644 14764 6696 14816
rect 7012 14764 7064 14816
rect 8208 14764 8260 14816
rect 9404 14764 9456 14816
rect 10508 14807 10560 14816
rect 10508 14773 10517 14807
rect 10517 14773 10551 14807
rect 10551 14773 10560 14807
rect 10508 14764 10560 14773
rect 10876 14764 10928 14816
rect 11704 14807 11756 14816
rect 11704 14773 11713 14807
rect 11713 14773 11747 14807
rect 11747 14773 11756 14807
rect 16212 14832 16264 14884
rect 16856 14807 16908 14816
rect 11704 14764 11756 14773
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 3915 14662 3967 14714
rect 3979 14662 4031 14714
rect 4043 14662 4095 14714
rect 4107 14662 4159 14714
rect 4171 14662 4223 14714
rect 9846 14662 9898 14714
rect 9910 14662 9962 14714
rect 9974 14662 10026 14714
rect 10038 14662 10090 14714
rect 10102 14662 10154 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 15904 14662 15956 14714
rect 15968 14662 16020 14714
rect 16032 14662 16084 14714
rect 4896 14560 4948 14612
rect 5724 14560 5776 14612
rect 6276 14603 6328 14612
rect 6276 14569 6285 14603
rect 6285 14569 6319 14603
rect 6319 14569 6328 14603
rect 6276 14560 6328 14569
rect 9312 14560 9364 14612
rect 9680 14560 9732 14612
rect 10784 14560 10836 14612
rect 10968 14603 11020 14612
rect 10968 14569 10977 14603
rect 10977 14569 11011 14603
rect 11011 14569 11020 14603
rect 10968 14560 11020 14569
rect 11980 14560 12032 14612
rect 16764 14560 16816 14612
rect 17868 14603 17920 14612
rect 17868 14569 17877 14603
rect 17877 14569 17911 14603
rect 17911 14569 17920 14603
rect 17868 14560 17920 14569
rect 3700 14424 3752 14476
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 4252 14399 4304 14408
rect 4252 14365 4261 14399
rect 4261 14365 4295 14399
rect 4295 14365 4304 14399
rect 4252 14356 4304 14365
rect 6920 14492 6972 14544
rect 7380 14492 7432 14544
rect 7288 14424 7340 14476
rect 8300 14492 8352 14544
rect 8944 14535 8996 14544
rect 8944 14501 8953 14535
rect 8953 14501 8987 14535
rect 8987 14501 8996 14535
rect 8944 14492 8996 14501
rect 10140 14492 10192 14544
rect 12624 14492 12676 14544
rect 10876 14424 10928 14476
rect 14004 14492 14056 14544
rect 4344 14288 4396 14340
rect 4988 14331 5040 14340
rect 4988 14297 4997 14331
rect 4997 14297 5031 14331
rect 5031 14297 5040 14331
rect 4988 14288 5040 14297
rect 5540 14288 5592 14340
rect 5724 14356 5776 14408
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 7012 14399 7064 14408
rect 7012 14365 7021 14399
rect 7021 14365 7055 14399
rect 7055 14365 7064 14399
rect 7012 14356 7064 14365
rect 5816 14288 5868 14340
rect 6000 14288 6052 14340
rect 7104 14288 7156 14340
rect 5264 14220 5316 14272
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 7288 14220 7340 14229
rect 7472 14220 7524 14272
rect 7748 14399 7800 14408
rect 7748 14365 7758 14399
rect 7758 14365 7792 14399
rect 7792 14365 7800 14399
rect 7748 14356 7800 14365
rect 8300 14331 8352 14340
rect 8300 14297 8309 14331
rect 8309 14297 8343 14331
rect 8343 14297 8352 14331
rect 8300 14288 8352 14297
rect 8484 14331 8536 14340
rect 8484 14297 8493 14331
rect 8493 14297 8527 14331
rect 8527 14297 8536 14331
rect 8484 14288 8536 14297
rect 9036 14288 9088 14340
rect 7932 14220 7984 14272
rect 8116 14263 8168 14272
rect 8116 14229 8125 14263
rect 8125 14229 8159 14263
rect 8159 14229 8168 14263
rect 8116 14220 8168 14229
rect 9588 14356 9640 14408
rect 11244 14356 11296 14408
rect 12532 14356 12584 14408
rect 9772 14288 9824 14340
rect 10692 14288 10744 14340
rect 11152 14331 11204 14340
rect 11152 14297 11161 14331
rect 11161 14297 11195 14331
rect 11195 14297 11204 14331
rect 11152 14288 11204 14297
rect 11336 14331 11388 14340
rect 11336 14297 11345 14331
rect 11345 14297 11379 14331
rect 11379 14297 11388 14331
rect 11336 14288 11388 14297
rect 12440 14288 12492 14340
rect 13268 14356 13320 14408
rect 14096 14356 14148 14408
rect 9312 14220 9364 14272
rect 9680 14220 9732 14272
rect 10232 14263 10284 14272
rect 10232 14229 10241 14263
rect 10241 14229 10275 14263
rect 10275 14229 10284 14263
rect 10232 14220 10284 14229
rect 13360 14263 13412 14272
rect 13360 14229 13369 14263
rect 13369 14229 13403 14263
rect 13403 14229 13412 14263
rect 13360 14220 13412 14229
rect 14464 14263 14516 14272
rect 14464 14229 14473 14263
rect 14473 14229 14507 14263
rect 14507 14229 14516 14263
rect 14464 14220 14516 14229
rect 15568 14356 15620 14408
rect 16120 14399 16172 14408
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 18328 14399 18380 14408
rect 18328 14365 18337 14399
rect 18337 14365 18371 14399
rect 18371 14365 18380 14399
rect 18328 14356 18380 14365
rect 18236 14288 18288 14340
rect 15384 14220 15436 14272
rect 15568 14263 15620 14272
rect 15568 14229 15577 14263
rect 15577 14229 15611 14263
rect 15611 14229 15620 14263
rect 15568 14220 15620 14229
rect 6880 14118 6932 14170
rect 6944 14118 6996 14170
rect 7008 14118 7060 14170
rect 7072 14118 7124 14170
rect 7136 14118 7188 14170
rect 12811 14118 12863 14170
rect 12875 14118 12927 14170
rect 12939 14118 12991 14170
rect 13003 14118 13055 14170
rect 13067 14118 13119 14170
rect 6000 14016 6052 14068
rect 7380 14016 7432 14068
rect 5172 13948 5224 14000
rect 6092 13948 6144 14000
rect 3608 13923 3660 13932
rect 3608 13889 3642 13923
rect 3642 13889 3660 13923
rect 3608 13880 3660 13889
rect 4528 13880 4580 13932
rect 4988 13880 5040 13932
rect 5724 13880 5776 13932
rect 4344 13812 4396 13864
rect 7472 13880 7524 13932
rect 7748 13923 7800 13932
rect 7748 13889 7757 13923
rect 7757 13889 7791 13923
rect 7791 13889 7800 13923
rect 7748 13880 7800 13889
rect 7932 13880 7984 13932
rect 8852 13948 8904 14000
rect 9404 13948 9456 14000
rect 11152 14016 11204 14068
rect 8852 13812 8904 13864
rect 5264 13744 5316 13796
rect 9680 13880 9732 13932
rect 10784 13948 10836 14000
rect 13268 14016 13320 14068
rect 14464 14016 14516 14068
rect 15200 14016 15252 14068
rect 16672 14016 16724 14068
rect 10140 13923 10192 13932
rect 10140 13889 10149 13923
rect 10149 13889 10183 13923
rect 10183 13889 10192 13923
rect 10140 13880 10192 13889
rect 12348 13948 12400 14000
rect 12256 13923 12308 13932
rect 12256 13889 12265 13923
rect 12265 13889 12299 13923
rect 12299 13889 12308 13923
rect 12256 13880 12308 13889
rect 12716 13923 12768 13932
rect 12716 13889 12725 13923
rect 12725 13889 12759 13923
rect 12759 13889 12768 13923
rect 12716 13880 12768 13889
rect 13360 13948 13412 14000
rect 14648 13880 14700 13932
rect 15292 13880 15344 13932
rect 16580 13880 16632 13932
rect 16764 13880 16816 13932
rect 12624 13812 12676 13864
rect 4712 13719 4764 13728
rect 4712 13685 4721 13719
rect 4721 13685 4755 13719
rect 4755 13685 4764 13719
rect 5540 13719 5592 13728
rect 4712 13676 4764 13685
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 6552 13676 6604 13728
rect 6644 13719 6696 13728
rect 6644 13685 6653 13719
rect 6653 13685 6687 13719
rect 6687 13685 6696 13719
rect 6644 13676 6696 13685
rect 7932 13676 7984 13728
rect 8208 13676 8260 13728
rect 10508 13744 10560 13796
rect 10692 13787 10744 13796
rect 10692 13753 10701 13787
rect 10701 13753 10735 13787
rect 10735 13753 10744 13787
rect 10692 13744 10744 13753
rect 9588 13676 9640 13728
rect 11796 13719 11848 13728
rect 11796 13685 11805 13719
rect 11805 13685 11839 13719
rect 11839 13685 11848 13719
rect 11796 13676 11848 13685
rect 14096 13719 14148 13728
rect 14096 13685 14105 13719
rect 14105 13685 14139 13719
rect 14139 13685 14148 13719
rect 14096 13676 14148 13685
rect 3915 13574 3967 13626
rect 3979 13574 4031 13626
rect 4043 13574 4095 13626
rect 4107 13574 4159 13626
rect 4171 13574 4223 13626
rect 9846 13574 9898 13626
rect 9910 13574 9962 13626
rect 9974 13574 10026 13626
rect 10038 13574 10090 13626
rect 10102 13574 10154 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 15904 13574 15956 13626
rect 15968 13574 16020 13626
rect 16032 13574 16084 13626
rect 3608 13472 3660 13524
rect 5264 13515 5316 13524
rect 1860 13268 1912 13320
rect 3792 13268 3844 13320
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 5356 13472 5408 13524
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 7380 13472 7432 13524
rect 8208 13515 8260 13524
rect 8208 13481 8217 13515
rect 8217 13481 8251 13515
rect 8251 13481 8260 13515
rect 8208 13472 8260 13481
rect 11888 13472 11940 13524
rect 18236 13472 18288 13524
rect 11060 13404 11112 13456
rect 11244 13447 11296 13456
rect 11244 13413 11253 13447
rect 11253 13413 11287 13447
rect 11287 13413 11296 13447
rect 11244 13404 11296 13413
rect 12716 13404 12768 13456
rect 2596 13200 2648 13252
rect 4528 13268 4580 13320
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 5448 13311 5500 13320
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 5448 13268 5500 13277
rect 7840 13311 7892 13320
rect 5264 13200 5316 13252
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 7932 13268 7984 13320
rect 9036 13268 9088 13320
rect 11428 13268 11480 13320
rect 15384 13404 15436 13456
rect 15200 13336 15252 13388
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 16580 13336 16632 13388
rect 16948 13379 17000 13388
rect 16948 13345 16957 13379
rect 16957 13345 16991 13379
rect 16991 13345 17000 13379
rect 16948 13336 17000 13345
rect 6736 13200 6788 13252
rect 4252 13132 4304 13184
rect 5540 13132 5592 13184
rect 7288 13132 7340 13184
rect 8116 13200 8168 13252
rect 10416 13200 10468 13252
rect 11796 13243 11848 13252
rect 11796 13209 11830 13243
rect 11830 13209 11848 13243
rect 11796 13200 11848 13209
rect 13452 13200 13504 13252
rect 14372 13243 14424 13252
rect 14372 13209 14381 13243
rect 14381 13209 14415 13243
rect 14415 13209 14424 13243
rect 14372 13200 14424 13209
rect 16672 13268 16724 13320
rect 9220 13132 9272 13184
rect 13176 13132 13228 13184
rect 13728 13132 13780 13184
rect 15016 13132 15068 13184
rect 16488 13200 16540 13252
rect 16856 13200 16908 13252
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 17040 13132 17092 13184
rect 6880 13030 6932 13082
rect 6944 13030 6996 13082
rect 7008 13030 7060 13082
rect 7072 13030 7124 13082
rect 7136 13030 7188 13082
rect 12811 13030 12863 13082
rect 12875 13030 12927 13082
rect 12939 13030 12991 13082
rect 13003 13030 13055 13082
rect 13067 13030 13119 13082
rect 2596 12971 2648 12980
rect 2596 12937 2605 12971
rect 2605 12937 2639 12971
rect 2639 12937 2648 12971
rect 2596 12928 2648 12937
rect 3792 12928 3844 12980
rect 5172 12928 5224 12980
rect 10416 12971 10468 12980
rect 5632 12860 5684 12912
rect 7564 12860 7616 12912
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 5540 12792 5592 12844
rect 5724 12792 5776 12844
rect 3700 12656 3752 12708
rect 5264 12724 5316 12776
rect 5356 12656 5408 12708
rect 5724 12656 5776 12708
rect 7196 12792 7248 12844
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 13176 12971 13228 12980
rect 13176 12937 13185 12971
rect 13185 12937 13219 12971
rect 13219 12937 13228 12971
rect 13176 12928 13228 12937
rect 12348 12860 12400 12912
rect 14096 12860 14148 12912
rect 9312 12835 9364 12844
rect 9312 12801 9321 12835
rect 9321 12801 9355 12835
rect 9355 12801 9364 12835
rect 9312 12792 9364 12801
rect 10692 12835 10744 12844
rect 9036 12767 9088 12776
rect 9036 12733 9045 12767
rect 9045 12733 9079 12767
rect 9079 12733 9088 12767
rect 9036 12724 9088 12733
rect 9220 12724 9272 12776
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 11060 12835 11112 12844
rect 10876 12792 10928 12801
rect 11060 12801 11069 12835
rect 11069 12801 11103 12835
rect 11103 12801 11112 12835
rect 11060 12792 11112 12801
rect 11244 12792 11296 12844
rect 12532 12792 12584 12844
rect 15016 12860 15068 12912
rect 12624 12656 12676 12708
rect 14372 12724 14424 12776
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 15292 12928 15344 12980
rect 16764 12928 16816 12980
rect 17040 12928 17092 12980
rect 18236 12971 18288 12980
rect 18236 12937 18245 12971
rect 18245 12937 18279 12971
rect 18279 12937 18288 12971
rect 18236 12928 18288 12937
rect 15660 12835 15712 12844
rect 14924 12792 14976 12801
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 15384 12724 15436 12776
rect 16396 12792 16448 12844
rect 17776 12792 17828 12844
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 16488 12724 16540 12776
rect 13728 12656 13780 12708
rect 14740 12656 14792 12708
rect 15936 12656 15988 12708
rect 1952 12588 2004 12640
rect 3056 12631 3108 12640
rect 3056 12597 3065 12631
rect 3065 12597 3099 12631
rect 3099 12597 3108 12631
rect 3056 12588 3108 12597
rect 4252 12588 4304 12640
rect 5264 12588 5316 12640
rect 5448 12631 5500 12640
rect 5448 12597 5457 12631
rect 5457 12597 5491 12631
rect 5491 12597 5500 12631
rect 5448 12588 5500 12597
rect 5540 12588 5592 12640
rect 5816 12588 5868 12640
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 3915 12486 3967 12538
rect 3979 12486 4031 12538
rect 4043 12486 4095 12538
rect 4107 12486 4159 12538
rect 4171 12486 4223 12538
rect 9846 12486 9898 12538
rect 9910 12486 9962 12538
rect 9974 12486 10026 12538
rect 10038 12486 10090 12538
rect 10102 12486 10154 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 15904 12486 15956 12538
rect 15968 12486 16020 12538
rect 16032 12486 16084 12538
rect 3700 12384 3752 12436
rect 5356 12384 5408 12436
rect 5540 12384 5592 12436
rect 5724 12427 5776 12436
rect 5724 12393 5733 12427
rect 5733 12393 5767 12427
rect 5767 12393 5776 12427
rect 5724 12384 5776 12393
rect 6276 12427 6328 12436
rect 6276 12393 6285 12427
rect 6285 12393 6319 12427
rect 6319 12393 6328 12427
rect 6276 12384 6328 12393
rect 7196 12427 7248 12436
rect 7196 12393 7205 12427
rect 7205 12393 7239 12427
rect 7239 12393 7248 12427
rect 7196 12384 7248 12393
rect 7564 12384 7616 12436
rect 10876 12384 10928 12436
rect 12440 12384 12492 12436
rect 14740 12427 14792 12436
rect 14740 12393 14749 12427
rect 14749 12393 14783 12427
rect 14783 12393 14792 12427
rect 14740 12384 14792 12393
rect 15384 12427 15436 12436
rect 15384 12393 15393 12427
rect 15393 12393 15427 12427
rect 15427 12393 15436 12427
rect 15384 12384 15436 12393
rect 17132 12384 17184 12436
rect 1768 12180 1820 12232
rect 1952 12223 2004 12232
rect 1952 12189 1986 12223
rect 1986 12189 2004 12223
rect 1952 12180 2004 12189
rect 4252 12223 4304 12232
rect 4252 12189 4261 12223
rect 4261 12189 4295 12223
rect 4295 12189 4304 12223
rect 4252 12180 4304 12189
rect 4528 12316 4580 12368
rect 6736 12316 6788 12368
rect 5264 12248 5316 12300
rect 9036 12316 9088 12368
rect 12256 12316 12308 12368
rect 5080 12180 5132 12232
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 7288 12248 7340 12300
rect 8852 12248 8904 12300
rect 9220 12291 9272 12300
rect 9220 12257 9229 12291
rect 9229 12257 9263 12291
rect 9263 12257 9272 12291
rect 9220 12248 9272 12257
rect 7656 12180 7708 12232
rect 5632 12112 5684 12164
rect 5816 12112 5868 12164
rect 9036 12112 9088 12164
rect 10324 12112 10376 12164
rect 3700 12044 3752 12096
rect 5540 12044 5592 12096
rect 9312 12044 9364 12096
rect 11612 12112 11664 12164
rect 12072 12180 12124 12232
rect 12532 12248 12584 12300
rect 12624 12180 12676 12232
rect 13268 12180 13320 12232
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 15660 12180 15712 12232
rect 16212 12223 16264 12232
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 16672 12248 16724 12300
rect 16396 12223 16448 12232
rect 16396 12189 16405 12223
rect 16405 12189 16439 12223
rect 16439 12189 16448 12223
rect 16396 12180 16448 12189
rect 16764 12180 16816 12232
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 14740 12112 14792 12164
rect 15292 12112 15344 12164
rect 12716 12044 12768 12096
rect 13176 12044 13228 12096
rect 14464 12044 14516 12096
rect 6880 11942 6932 11994
rect 6944 11942 6996 11994
rect 7008 11942 7060 11994
rect 7072 11942 7124 11994
rect 7136 11942 7188 11994
rect 12811 11942 12863 11994
rect 12875 11942 12927 11994
rect 12939 11942 12991 11994
rect 13003 11942 13055 11994
rect 13067 11942 13119 11994
rect 5816 11840 5868 11892
rect 5908 11840 5960 11892
rect 3056 11772 3108 11824
rect 6276 11772 6328 11824
rect 7840 11772 7892 11824
rect 13728 11840 13780 11892
rect 13544 11772 13596 11824
rect 14924 11772 14976 11824
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 6552 11704 6604 11756
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 7472 11704 7524 11756
rect 9128 11704 9180 11756
rect 9312 11747 9364 11756
rect 9312 11713 9346 11747
rect 9346 11713 9364 11747
rect 9312 11704 9364 11713
rect 9588 11704 9640 11756
rect 3792 11679 3844 11688
rect 3792 11645 3801 11679
rect 3801 11645 3835 11679
rect 3835 11645 3844 11679
rect 3792 11636 3844 11645
rect 6092 11636 6144 11688
rect 10968 11704 11020 11756
rect 12624 11704 12676 11756
rect 15016 11747 15068 11756
rect 15016 11713 15025 11747
rect 15025 11713 15059 11747
rect 15059 11713 15068 11747
rect 15016 11704 15068 11713
rect 15660 11747 15712 11756
rect 1400 11611 1452 11620
rect 1400 11577 1409 11611
rect 1409 11577 1443 11611
rect 1443 11577 1452 11611
rect 1400 11568 1452 11577
rect 4988 11568 5040 11620
rect 3240 11543 3292 11552
rect 3240 11509 3249 11543
rect 3249 11509 3283 11543
rect 3283 11509 3292 11543
rect 3240 11500 3292 11509
rect 5172 11543 5224 11552
rect 5172 11509 5181 11543
rect 5181 11509 5215 11543
rect 5215 11509 5224 11543
rect 5172 11500 5224 11509
rect 6644 11568 6696 11620
rect 11336 11636 11388 11688
rect 11428 11636 11480 11688
rect 7564 11500 7616 11552
rect 10324 11500 10376 11552
rect 10784 11500 10836 11552
rect 12716 11500 12768 11552
rect 14648 11636 14700 11688
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 16396 11704 16448 11756
rect 16120 11636 16172 11688
rect 16764 11679 16816 11688
rect 16764 11645 16773 11679
rect 16773 11645 16807 11679
rect 16807 11645 16816 11679
rect 16764 11636 16816 11645
rect 14280 11500 14332 11552
rect 14464 11500 14516 11552
rect 16304 11500 16356 11552
rect 16580 11500 16632 11552
rect 17776 11500 17828 11552
rect 3915 11398 3967 11450
rect 3979 11398 4031 11450
rect 4043 11398 4095 11450
rect 4107 11398 4159 11450
rect 4171 11398 4223 11450
rect 9846 11398 9898 11450
rect 9910 11398 9962 11450
rect 9974 11398 10026 11450
rect 10038 11398 10090 11450
rect 10102 11398 10154 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 15904 11398 15956 11450
rect 15968 11398 16020 11450
rect 16032 11398 16084 11450
rect 3240 11296 3292 11348
rect 4160 11228 4212 11280
rect 5908 11296 5960 11348
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 6736 11296 6788 11348
rect 9312 11296 9364 11348
rect 10968 11339 11020 11348
rect 10968 11305 10977 11339
rect 10977 11305 11011 11339
rect 11011 11305 11020 11339
rect 10968 11296 11020 11305
rect 11336 11296 11388 11348
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 5172 11271 5224 11280
rect 2136 11160 2188 11212
rect 5172 11237 5181 11271
rect 5181 11237 5215 11271
rect 5215 11237 5224 11271
rect 5172 11228 5224 11237
rect 7472 11228 7524 11280
rect 8852 11228 8904 11280
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 3700 11024 3752 11076
rect 2320 10956 2372 11008
rect 5356 11160 5408 11212
rect 4988 11067 5040 11076
rect 4988 11033 4997 11067
rect 4997 11033 5031 11067
rect 5031 11033 5040 11067
rect 4988 11024 5040 11033
rect 5540 11135 5592 11144
rect 5540 11101 5549 11135
rect 5549 11101 5583 11135
rect 5583 11101 5592 11135
rect 5540 11092 5592 11101
rect 6000 11092 6052 11144
rect 7564 11160 7616 11212
rect 16212 11228 16264 11280
rect 6736 11092 6788 11144
rect 7656 11092 7708 11144
rect 8116 11092 8168 11144
rect 12164 11160 12216 11212
rect 16488 11160 16540 11212
rect 9588 11092 9640 11144
rect 9772 11092 9824 11144
rect 10600 11092 10652 11144
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 15568 11092 15620 11144
rect 16580 11135 16632 11144
rect 16580 11101 16589 11135
rect 16589 11101 16623 11135
rect 16623 11101 16632 11135
rect 16580 11092 16632 11101
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 5540 10956 5592 11008
rect 7564 11024 7616 11076
rect 10324 11024 10376 11076
rect 11152 11024 11204 11076
rect 12072 11024 12124 11076
rect 12716 11024 12768 11076
rect 13268 11067 13320 11076
rect 13268 11033 13277 11067
rect 13277 11033 13311 11067
rect 13311 11033 13320 11067
rect 13268 11024 13320 11033
rect 13452 11067 13504 11076
rect 13452 11033 13461 11067
rect 13461 11033 13495 11067
rect 13495 11033 13504 11067
rect 13452 11024 13504 11033
rect 14004 11024 14056 11076
rect 14556 11024 14608 11076
rect 14924 11067 14976 11076
rect 14924 11033 14933 11067
rect 14933 11033 14967 11067
rect 14967 11033 14976 11067
rect 14924 11024 14976 11033
rect 15016 11024 15068 11076
rect 15660 11067 15712 11076
rect 15660 11033 15669 11067
rect 15669 11033 15703 11067
rect 15703 11033 15712 11067
rect 15660 11024 15712 11033
rect 16304 11024 16356 11076
rect 17592 11024 17644 11076
rect 7288 10956 7340 11008
rect 10968 10956 11020 11008
rect 12256 10956 12308 11008
rect 17868 10956 17920 11008
rect 6880 10854 6932 10906
rect 6944 10854 6996 10906
rect 7008 10854 7060 10906
rect 7072 10854 7124 10906
rect 7136 10854 7188 10906
rect 12811 10854 12863 10906
rect 12875 10854 12927 10906
rect 12939 10854 12991 10906
rect 13003 10854 13055 10906
rect 13067 10854 13119 10906
rect 5080 10752 5132 10804
rect 9772 10795 9824 10804
rect 3792 10684 3844 10736
rect 1860 10616 1912 10668
rect 2044 10659 2096 10668
rect 2044 10625 2078 10659
rect 2078 10625 2096 10659
rect 6000 10684 6052 10736
rect 7472 10684 7524 10736
rect 7748 10684 7800 10736
rect 9772 10761 9781 10795
rect 9781 10761 9815 10795
rect 9815 10761 9824 10795
rect 9772 10752 9824 10761
rect 11152 10752 11204 10804
rect 13176 10752 13228 10804
rect 14280 10752 14332 10804
rect 2044 10616 2096 10625
rect 4160 10659 4212 10668
rect 4160 10625 4194 10659
rect 4194 10625 4212 10659
rect 4160 10616 4212 10625
rect 5540 10616 5592 10668
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 10692 10684 10744 10736
rect 11336 10684 11388 10736
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 10232 10616 10284 10668
rect 11520 10616 11572 10668
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 7472 10548 7524 10600
rect 9772 10548 9824 10600
rect 11980 10548 12032 10600
rect 12256 10616 12308 10668
rect 13452 10684 13504 10736
rect 12624 10548 12676 10600
rect 14096 10616 14148 10668
rect 14280 10659 14332 10668
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 14556 10659 14608 10668
rect 14556 10625 14590 10659
rect 14590 10625 14608 10659
rect 14556 10616 14608 10625
rect 16764 10616 16816 10668
rect 16948 10659 17000 10668
rect 16948 10625 16982 10659
rect 16982 10625 17000 10659
rect 16948 10616 17000 10625
rect 13544 10548 13596 10600
rect 6644 10480 6696 10532
rect 7564 10523 7616 10532
rect 7564 10489 7573 10523
rect 7573 10489 7607 10523
rect 7607 10489 7616 10523
rect 7564 10480 7616 10489
rect 13268 10480 13320 10532
rect 15476 10480 15528 10532
rect 15660 10523 15712 10532
rect 15660 10489 15669 10523
rect 15669 10489 15703 10523
rect 15703 10489 15712 10523
rect 15660 10480 15712 10489
rect 2872 10412 2924 10464
rect 5264 10455 5316 10464
rect 5264 10421 5273 10455
rect 5273 10421 5307 10455
rect 5307 10421 5316 10455
rect 5264 10412 5316 10421
rect 7932 10412 7984 10464
rect 9588 10412 9640 10464
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 12256 10412 12308 10464
rect 15384 10412 15436 10464
rect 16212 10412 16264 10464
rect 3915 10310 3967 10362
rect 3979 10310 4031 10362
rect 4043 10310 4095 10362
rect 4107 10310 4159 10362
rect 4171 10310 4223 10362
rect 9846 10310 9898 10362
rect 9910 10310 9962 10362
rect 9974 10310 10026 10362
rect 10038 10310 10090 10362
rect 10102 10310 10154 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 15904 10310 15956 10362
rect 15968 10310 16020 10362
rect 16032 10310 16084 10362
rect 2044 10208 2096 10260
rect 2412 10208 2464 10260
rect 5356 10251 5408 10260
rect 5356 10217 5365 10251
rect 5365 10217 5399 10251
rect 5399 10217 5408 10251
rect 5356 10208 5408 10217
rect 14188 10208 14240 10260
rect 18052 10208 18104 10260
rect 7748 10140 7800 10192
rect 3148 10072 3200 10124
rect 11428 10072 11480 10124
rect 16120 10115 16172 10124
rect 16120 10081 16129 10115
rect 16129 10081 16163 10115
rect 16163 10081 16172 10115
rect 16120 10072 16172 10081
rect 16764 10072 16816 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 4344 10004 4396 10056
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 5540 10004 5592 10056
rect 7656 10004 7708 10056
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 10416 10004 10468 10056
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 11704 10004 11756 10056
rect 11980 10004 12032 10056
rect 2872 9936 2924 9988
rect 4620 9936 4672 9988
rect 6736 9936 6788 9988
rect 9312 9936 9364 9988
rect 10784 9936 10836 9988
rect 12348 9936 12400 9988
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 5724 9868 5776 9920
rect 7564 9868 7616 9920
rect 9680 9868 9732 9920
rect 10692 9868 10744 9920
rect 10876 9911 10928 9920
rect 10876 9877 10885 9911
rect 10885 9877 10919 9911
rect 10919 9877 10928 9911
rect 10876 9868 10928 9877
rect 12624 9868 12676 9920
rect 14280 10004 14332 10056
rect 17776 10004 17828 10056
rect 13820 9936 13872 9988
rect 17316 9936 17368 9988
rect 13912 9868 13964 9920
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 14464 9868 14516 9920
rect 15292 9868 15344 9920
rect 15660 9868 15712 9920
rect 16212 9911 16264 9920
rect 16212 9877 16221 9911
rect 16221 9877 16255 9911
rect 16255 9877 16264 9911
rect 16212 9868 16264 9877
rect 16856 9868 16908 9920
rect 6880 9766 6932 9818
rect 6944 9766 6996 9818
rect 7008 9766 7060 9818
rect 7072 9766 7124 9818
rect 7136 9766 7188 9818
rect 12811 9766 12863 9818
rect 12875 9766 12927 9818
rect 12939 9766 12991 9818
rect 13003 9766 13055 9818
rect 13067 9766 13119 9818
rect 6736 9664 6788 9716
rect 5540 9596 5592 9648
rect 7564 9664 7616 9716
rect 8116 9664 8168 9716
rect 9680 9664 9732 9716
rect 10784 9664 10836 9716
rect 10876 9664 10928 9716
rect 13636 9664 13688 9716
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 4252 9528 4304 9580
rect 5724 9571 5776 9580
rect 5724 9537 5742 9571
rect 5742 9537 5776 9571
rect 6000 9571 6052 9580
rect 5724 9528 5776 9537
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 7288 9571 7340 9580
rect 4712 9460 4764 9512
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 7748 9596 7800 9648
rect 12532 9596 12584 9648
rect 12624 9639 12676 9648
rect 12624 9605 12642 9639
rect 12642 9605 12676 9639
rect 12624 9596 12676 9605
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 7932 9571 7984 9580
rect 7932 9537 7966 9571
rect 7966 9537 7984 9571
rect 7932 9528 7984 9537
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 14556 9664 14608 9716
rect 14924 9664 14976 9716
rect 17316 9707 17368 9716
rect 17316 9673 17325 9707
rect 17325 9673 17359 9707
rect 17359 9673 17368 9707
rect 17316 9664 17368 9673
rect 14096 9528 14148 9580
rect 14188 9528 14240 9580
rect 16764 9596 16816 9648
rect 17592 9596 17644 9648
rect 18236 9639 18288 9648
rect 18236 9605 18245 9639
rect 18245 9605 18279 9639
rect 18279 9605 18288 9639
rect 18236 9596 18288 9605
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 17408 9528 17460 9580
rect 17960 9528 18012 9580
rect 7472 9460 7524 9512
rect 14924 9460 14976 9512
rect 17040 9503 17092 9512
rect 17040 9469 17049 9503
rect 17049 9469 17083 9503
rect 17083 9469 17092 9503
rect 17040 9460 17092 9469
rect 17776 9503 17828 9512
rect 17776 9469 17785 9503
rect 17785 9469 17819 9503
rect 17819 9469 17828 9503
rect 17776 9460 17828 9469
rect 13820 9392 13872 9444
rect 16948 9392 17000 9444
rect 2780 9367 2832 9376
rect 2780 9333 2789 9367
rect 2789 9333 2823 9367
rect 2823 9333 2832 9367
rect 2780 9324 2832 9333
rect 4436 9324 4488 9376
rect 10416 9324 10468 9376
rect 10600 9367 10652 9376
rect 10600 9333 10609 9367
rect 10609 9333 10643 9367
rect 10643 9333 10652 9367
rect 10600 9324 10652 9333
rect 11336 9324 11388 9376
rect 13084 9324 13136 9376
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 17684 9367 17736 9376
rect 17684 9333 17693 9367
rect 17693 9333 17727 9367
rect 17727 9333 17736 9367
rect 17684 9324 17736 9333
rect 3915 9222 3967 9274
rect 3979 9222 4031 9274
rect 4043 9222 4095 9274
rect 4107 9222 4159 9274
rect 4171 9222 4223 9274
rect 9846 9222 9898 9274
rect 9910 9222 9962 9274
rect 9974 9222 10026 9274
rect 10038 9222 10090 9274
rect 10102 9222 10154 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 15904 9222 15956 9274
rect 15968 9222 16020 9274
rect 16032 9222 16084 9274
rect 4252 9120 4304 9172
rect 7840 9120 7892 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 10232 9120 10284 9172
rect 10416 9120 10468 9172
rect 11152 9120 11204 9172
rect 11520 9163 11572 9172
rect 11520 9129 11529 9163
rect 11529 9129 11563 9163
rect 11563 9129 11572 9163
rect 11520 9120 11572 9129
rect 11796 9120 11848 9172
rect 12348 9120 12400 9172
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 14188 9120 14240 9172
rect 17776 9163 17828 9172
rect 6552 9095 6604 9104
rect 6552 9061 6561 9095
rect 6561 9061 6595 9095
rect 6595 9061 6604 9095
rect 6552 9052 6604 9061
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 2780 8916 2832 8968
rect 5448 8916 5500 8968
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 10600 8984 10652 9036
rect 11980 9052 12032 9104
rect 12164 9052 12216 9104
rect 11244 8984 11296 9036
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 8208 8916 8260 8968
rect 2872 8848 2924 8900
rect 5264 8891 5316 8900
rect 5264 8857 5273 8891
rect 5273 8857 5307 8891
rect 5307 8857 5316 8891
rect 5264 8848 5316 8857
rect 8760 8916 8812 8968
rect 9588 8959 9640 8968
rect 9588 8925 9597 8959
rect 9597 8925 9631 8959
rect 9631 8925 9640 8959
rect 9588 8916 9640 8925
rect 9680 8916 9732 8968
rect 10968 8916 11020 8968
rect 12532 8984 12584 9036
rect 9496 8848 9548 8900
rect 2780 8780 2832 8832
rect 3424 8823 3476 8832
rect 3424 8789 3433 8823
rect 3433 8789 3467 8823
rect 3467 8789 3476 8823
rect 3424 8780 3476 8789
rect 4436 8823 4488 8832
rect 4436 8789 4445 8823
rect 4445 8789 4479 8823
rect 4479 8789 4488 8823
rect 4436 8780 4488 8789
rect 6460 8780 6512 8832
rect 8392 8780 8444 8832
rect 8484 8780 8536 8832
rect 11060 8848 11112 8900
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 11888 8916 11940 8968
rect 12256 8959 12308 8968
rect 11704 8848 11756 8900
rect 12256 8925 12265 8959
rect 12265 8925 12299 8959
rect 12299 8925 12308 8959
rect 12256 8916 12308 8925
rect 13084 8984 13136 9036
rect 17776 9129 17785 9163
rect 17785 9129 17819 9163
rect 17819 9129 17828 9163
rect 17776 9120 17828 9129
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 13452 8916 13504 8968
rect 15568 8959 15620 8968
rect 15568 8925 15577 8959
rect 15577 8925 15611 8959
rect 15611 8925 15620 8959
rect 15568 8916 15620 8925
rect 17040 8984 17092 9036
rect 16120 8916 16172 8968
rect 16396 8959 16448 8968
rect 16396 8925 16405 8959
rect 16405 8925 16439 8959
rect 16439 8925 16448 8959
rect 16396 8916 16448 8925
rect 17500 8959 17552 8968
rect 17500 8925 17509 8959
rect 17509 8925 17543 8959
rect 17543 8925 17552 8959
rect 17500 8916 17552 8925
rect 17960 8959 18012 8968
rect 17960 8925 17969 8959
rect 17969 8925 18003 8959
rect 18003 8925 18012 8959
rect 17960 8916 18012 8925
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 12716 8848 12768 8900
rect 13544 8780 13596 8832
rect 16488 8848 16540 8900
rect 14004 8780 14056 8832
rect 14188 8780 14240 8832
rect 14556 8823 14608 8832
rect 14556 8789 14565 8823
rect 14565 8789 14599 8823
rect 14599 8789 14608 8823
rect 14556 8780 14608 8789
rect 15200 8780 15252 8832
rect 15568 8780 15620 8832
rect 16212 8780 16264 8832
rect 17040 8823 17092 8832
rect 17040 8789 17049 8823
rect 17049 8789 17083 8823
rect 17083 8789 17092 8823
rect 17040 8780 17092 8789
rect 6880 8678 6932 8730
rect 6944 8678 6996 8730
rect 7008 8678 7060 8730
rect 7072 8678 7124 8730
rect 7136 8678 7188 8730
rect 12811 8678 12863 8730
rect 12875 8678 12927 8730
rect 12939 8678 12991 8730
rect 13003 8678 13055 8730
rect 13067 8678 13119 8730
rect 1492 8619 1544 8628
rect 1492 8585 1501 8619
rect 1501 8585 1535 8619
rect 1535 8585 1544 8619
rect 1492 8576 1544 8585
rect 2320 8576 2372 8628
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 7748 8619 7800 8628
rect 3424 8508 3476 8560
rect 4804 8508 4856 8560
rect 5632 8483 5684 8492
rect 2780 8372 2832 8424
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 7748 8585 7757 8619
rect 7757 8585 7791 8619
rect 7791 8585 7800 8619
rect 7748 8576 7800 8585
rect 8116 8576 8168 8628
rect 7288 8508 7340 8560
rect 8392 8551 8444 8560
rect 8392 8517 8401 8551
rect 8401 8517 8435 8551
rect 8435 8517 8444 8551
rect 8392 8508 8444 8517
rect 6460 8440 6512 8492
rect 7472 8440 7524 8492
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 10876 8576 10928 8628
rect 11704 8576 11756 8628
rect 10232 8508 10284 8560
rect 10508 8508 10560 8560
rect 10600 8508 10652 8560
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 12624 8576 12676 8628
rect 9128 8440 9180 8449
rect 1584 8304 1636 8356
rect 2228 8236 2280 8288
rect 9680 8372 9732 8424
rect 7380 8236 7432 8288
rect 9496 8304 9548 8356
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 12256 8483 12308 8492
rect 12256 8449 12260 8483
rect 12260 8449 12294 8483
rect 12294 8449 12308 8483
rect 12256 8440 12308 8449
rect 12716 8440 12768 8492
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 14096 8576 14148 8628
rect 13544 8508 13596 8560
rect 17684 8576 17736 8628
rect 17040 8551 17092 8560
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 14004 8440 14056 8492
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 14464 8483 14516 8492
rect 14464 8449 14473 8483
rect 14473 8449 14507 8483
rect 14507 8449 14516 8483
rect 14464 8440 14516 8449
rect 17040 8517 17074 8551
rect 17074 8517 17092 8551
rect 17040 8508 17092 8517
rect 14924 8483 14976 8492
rect 10416 8236 10468 8288
rect 12532 8304 12584 8356
rect 13820 8372 13872 8424
rect 12164 8236 12216 8288
rect 13360 8304 13412 8356
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 16764 8483 16816 8492
rect 16764 8449 16773 8483
rect 16773 8449 16807 8483
rect 16807 8449 16816 8483
rect 16764 8440 16816 8449
rect 13544 8236 13596 8288
rect 14464 8236 14516 8288
rect 17500 8236 17552 8288
rect 18144 8279 18196 8288
rect 18144 8245 18153 8279
rect 18153 8245 18187 8279
rect 18187 8245 18196 8279
rect 18144 8236 18196 8245
rect 3915 8134 3967 8186
rect 3979 8134 4031 8186
rect 4043 8134 4095 8186
rect 4107 8134 4159 8186
rect 4171 8134 4223 8186
rect 9846 8134 9898 8186
rect 9910 8134 9962 8186
rect 9974 8134 10026 8186
rect 10038 8134 10090 8186
rect 10102 8134 10154 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 15904 8134 15956 8186
rect 15968 8134 16020 8186
rect 16032 8134 16084 8186
rect 5632 8032 5684 8084
rect 6092 8032 6144 8084
rect 3148 7896 3200 7948
rect 4344 7896 4396 7948
rect 4712 7896 4764 7948
rect 5908 7896 5960 7948
rect 7748 7964 7800 8016
rect 7840 7939 7892 7948
rect 2044 7828 2096 7880
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 5172 7828 5224 7880
rect 5540 7760 5592 7812
rect 6552 7828 6604 7880
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 8484 7896 8536 7948
rect 9128 7896 9180 7948
rect 11060 7896 11112 7948
rect 7380 7828 7432 7880
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 7748 7803 7800 7812
rect 7748 7769 7757 7803
rect 7757 7769 7791 7803
rect 7791 7769 7800 7803
rect 7748 7760 7800 7769
rect 10508 7760 10560 7812
rect 10876 7828 10928 7880
rect 12348 8032 12400 8084
rect 14096 8075 14148 8084
rect 14096 8041 14105 8075
rect 14105 8041 14139 8075
rect 14139 8041 14148 8075
rect 14096 8032 14148 8041
rect 14924 8032 14976 8084
rect 16396 8032 16448 8084
rect 12348 7871 12400 7880
rect 1952 7735 2004 7744
rect 1952 7701 1961 7735
rect 1961 7701 1995 7735
rect 1995 7701 2004 7735
rect 1952 7692 2004 7701
rect 2136 7692 2188 7744
rect 3056 7692 3108 7744
rect 8944 7692 8996 7744
rect 11520 7760 11572 7812
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 14556 7964 14608 8016
rect 16488 7964 16540 8016
rect 13452 7896 13504 7948
rect 14372 7896 14424 7948
rect 12716 7828 12768 7837
rect 13268 7828 13320 7880
rect 14280 7871 14332 7880
rect 12256 7760 12308 7812
rect 14280 7837 14284 7871
rect 14284 7837 14318 7871
rect 14318 7837 14332 7871
rect 14280 7828 14332 7837
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 14648 7871 14700 7880
rect 14648 7837 14656 7871
rect 14656 7837 14690 7871
rect 14690 7837 14700 7871
rect 14648 7828 14700 7837
rect 14924 7828 14976 7880
rect 16120 7896 16172 7948
rect 16304 7828 16356 7880
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 17224 7828 17276 7880
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 14556 7760 14608 7812
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 11428 7735 11480 7744
rect 11428 7701 11437 7735
rect 11437 7701 11471 7735
rect 11471 7701 11480 7735
rect 11428 7692 11480 7701
rect 12716 7692 12768 7744
rect 14924 7692 14976 7744
rect 18144 7692 18196 7744
rect 6880 7590 6932 7642
rect 6944 7590 6996 7642
rect 7008 7590 7060 7642
rect 7072 7590 7124 7642
rect 7136 7590 7188 7642
rect 12811 7590 12863 7642
rect 12875 7590 12927 7642
rect 12939 7590 12991 7642
rect 13003 7590 13055 7642
rect 13067 7590 13119 7642
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 9680 7531 9732 7540
rect 9680 7497 9689 7531
rect 9689 7497 9723 7531
rect 9723 7497 9732 7531
rect 9680 7488 9732 7497
rect 1952 7463 2004 7472
rect 1952 7429 1986 7463
rect 1986 7429 2004 7463
rect 1952 7420 2004 7429
rect 1584 7352 1636 7404
rect 6644 7420 6696 7472
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 5356 7395 5408 7404
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 2688 7284 2740 7336
rect 4804 7284 4856 7336
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 5908 7216 5960 7268
rect 6644 7259 6696 7268
rect 6644 7225 6653 7259
rect 6653 7225 6687 7259
rect 6687 7225 6696 7259
rect 6644 7216 6696 7225
rect 7380 7216 7432 7268
rect 3056 7191 3108 7200
rect 3056 7157 3065 7191
rect 3065 7157 3099 7191
rect 3099 7157 3108 7191
rect 3056 7148 3108 7157
rect 6276 7148 6328 7200
rect 8944 7420 8996 7472
rect 11152 7488 11204 7540
rect 10324 7420 10376 7472
rect 8576 7284 8628 7336
rect 9496 7284 9548 7336
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 12624 7420 12676 7472
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 11796 7327 11848 7336
rect 11796 7293 11805 7327
rect 11805 7293 11839 7327
rect 11839 7293 11848 7327
rect 11796 7284 11848 7293
rect 12256 7284 12308 7336
rect 12348 7284 12400 7336
rect 12992 7284 13044 7336
rect 14464 7488 14516 7540
rect 13912 7395 13964 7404
rect 13912 7361 13921 7395
rect 13921 7361 13955 7395
rect 13955 7361 13964 7395
rect 13912 7352 13964 7361
rect 9772 7216 9824 7268
rect 10876 7216 10928 7268
rect 10968 7216 11020 7268
rect 11152 7216 11204 7268
rect 12716 7216 12768 7268
rect 12900 7259 12952 7268
rect 12900 7225 12909 7259
rect 12909 7225 12943 7259
rect 12943 7225 12952 7259
rect 12900 7216 12952 7225
rect 10600 7148 10652 7200
rect 12624 7148 12676 7200
rect 13268 7148 13320 7200
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 14648 7352 14700 7404
rect 15016 7420 15068 7472
rect 15384 7463 15436 7472
rect 15384 7429 15393 7463
rect 15393 7429 15427 7463
rect 15427 7429 15436 7463
rect 15384 7420 15436 7429
rect 16580 7420 16632 7472
rect 14924 7352 14976 7404
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 15016 7284 15068 7336
rect 16212 7352 16264 7404
rect 16764 7352 16816 7404
rect 16488 7284 16540 7336
rect 14556 7216 14608 7268
rect 15108 7148 15160 7200
rect 15384 7148 15436 7200
rect 16120 7148 16172 7200
rect 16856 7148 16908 7200
rect 3915 7046 3967 7098
rect 3979 7046 4031 7098
rect 4043 7046 4095 7098
rect 4107 7046 4159 7098
rect 4171 7046 4223 7098
rect 9846 7046 9898 7098
rect 9910 7046 9962 7098
rect 9974 7046 10026 7098
rect 10038 7046 10090 7098
rect 10102 7046 10154 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 15904 7046 15956 7098
rect 15968 7046 16020 7098
rect 16032 7046 16084 7098
rect 2044 6944 2096 6996
rect 4896 6987 4948 6996
rect 4896 6953 4905 6987
rect 4905 6953 4939 6987
rect 4939 6953 4948 6987
rect 4896 6944 4948 6953
rect 8944 6987 8996 6996
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 1768 6808 1820 6860
rect 2688 6808 2740 6860
rect 3516 6808 3568 6860
rect 4804 6876 4856 6928
rect 8944 6953 8953 6987
rect 8953 6953 8987 6987
rect 8987 6953 8996 6987
rect 8944 6944 8996 6953
rect 11428 6944 11480 6996
rect 8208 6876 8260 6928
rect 9404 6876 9456 6928
rect 4344 6851 4396 6860
rect 4344 6817 4353 6851
rect 4353 6817 4387 6851
rect 4387 6817 4396 6851
rect 4344 6808 4396 6817
rect 7288 6808 7340 6860
rect 13452 6944 13504 6996
rect 14556 6944 14608 6996
rect 14924 6987 14976 6996
rect 14924 6953 14933 6987
rect 14933 6953 14967 6987
rect 14967 6953 14976 6987
rect 14924 6944 14976 6953
rect 16212 6944 16264 6996
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 4160 6740 4212 6792
rect 6276 6783 6328 6792
rect 6276 6749 6294 6783
rect 6294 6749 6328 6783
rect 6276 6740 6328 6749
rect 7656 6740 7708 6792
rect 9680 6740 9732 6792
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 11704 6808 11756 6860
rect 12348 6851 12400 6860
rect 10232 6740 10284 6749
rect 11060 6740 11112 6792
rect 11336 6740 11388 6792
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 12348 6817 12357 6851
rect 12357 6817 12391 6851
rect 12391 6817 12400 6851
rect 12348 6808 12400 6817
rect 12440 6808 12492 6860
rect 12716 6808 12768 6860
rect 13820 6808 13872 6860
rect 13912 6808 13964 6860
rect 14280 6808 14332 6860
rect 15016 6808 15068 6860
rect 15568 6808 15620 6860
rect 13452 6740 13504 6792
rect 14556 6740 14608 6792
rect 14924 6740 14976 6792
rect 15384 6783 15436 6792
rect 5356 6672 5408 6724
rect 7564 6672 7616 6724
rect 10324 6672 10376 6724
rect 10508 6672 10560 6724
rect 2596 6647 2648 6656
rect 2596 6613 2605 6647
rect 2605 6613 2639 6647
rect 2639 6613 2648 6647
rect 2596 6604 2648 6613
rect 3056 6604 3108 6656
rect 4528 6647 4580 6656
rect 4528 6613 4537 6647
rect 4537 6613 4571 6647
rect 4571 6613 4580 6647
rect 5172 6647 5224 6656
rect 4528 6604 4580 6613
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 8116 6647 8168 6656
rect 8116 6613 8125 6647
rect 8125 6613 8159 6647
rect 8159 6613 8168 6647
rect 8116 6604 8168 6613
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 10140 6647 10192 6656
rect 10140 6613 10149 6647
rect 10149 6613 10183 6647
rect 10183 6613 10192 6647
rect 10140 6604 10192 6613
rect 10876 6647 10928 6656
rect 10876 6613 10885 6647
rect 10885 6613 10919 6647
rect 10919 6613 10928 6647
rect 10876 6604 10928 6613
rect 12992 6672 13044 6724
rect 13820 6672 13872 6724
rect 13912 6672 13964 6724
rect 15016 6672 15068 6724
rect 11796 6604 11848 6656
rect 11980 6647 12032 6656
rect 11980 6613 11989 6647
rect 11989 6613 12023 6647
rect 12023 6613 12032 6647
rect 11980 6604 12032 6613
rect 12256 6604 12308 6656
rect 12624 6604 12676 6656
rect 14556 6604 14608 6656
rect 15384 6749 15393 6783
rect 15393 6749 15427 6783
rect 15427 6749 15436 6783
rect 15384 6740 15436 6749
rect 16120 6740 16172 6792
rect 16672 6808 16724 6860
rect 16948 6808 17000 6860
rect 18236 6740 18288 6792
rect 15568 6672 15620 6724
rect 16212 6672 16264 6724
rect 15660 6604 15712 6656
rect 16580 6604 16632 6656
rect 16856 6604 16908 6656
rect 17868 6672 17920 6724
rect 6880 6502 6932 6554
rect 6944 6502 6996 6554
rect 7008 6502 7060 6554
rect 7072 6502 7124 6554
rect 7136 6502 7188 6554
rect 12811 6502 12863 6554
rect 12875 6502 12927 6554
rect 12939 6502 12991 6554
rect 13003 6502 13055 6554
rect 13067 6502 13119 6554
rect 3056 6400 3108 6452
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 5172 6400 5224 6452
rect 7288 6400 7340 6452
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 8300 6400 8352 6452
rect 10048 6400 10100 6452
rect 10232 6400 10284 6452
rect 11152 6443 11204 6452
rect 11152 6409 11161 6443
rect 11161 6409 11195 6443
rect 11195 6409 11204 6443
rect 11152 6400 11204 6409
rect 2964 6375 3016 6384
rect 2964 6341 2973 6375
rect 2973 6341 3007 6375
rect 3007 6341 3016 6375
rect 2964 6332 3016 6341
rect 5540 6332 5592 6384
rect 6920 6332 6972 6384
rect 8392 6375 8444 6384
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 3148 6239 3200 6248
rect 3148 6205 3157 6239
rect 3157 6205 3191 6239
rect 3191 6205 3200 6239
rect 3148 6196 3200 6205
rect 3516 6239 3568 6248
rect 3516 6205 3525 6239
rect 3525 6205 3559 6239
rect 3559 6205 3568 6239
rect 3516 6196 3568 6205
rect 3792 6264 3844 6316
rect 5908 6307 5960 6316
rect 4344 6196 4396 6248
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 8392 6341 8401 6375
rect 8401 6341 8435 6375
rect 8435 6341 8444 6375
rect 8392 6332 8444 6341
rect 8576 6332 8628 6384
rect 8024 6264 8076 6316
rect 7380 6196 7432 6248
rect 8208 6264 8260 6316
rect 8760 6264 8812 6316
rect 10508 6264 10560 6316
rect 10971 6307 11023 6316
rect 10971 6273 10980 6307
rect 10980 6273 11014 6307
rect 11014 6273 11023 6307
rect 10971 6264 11023 6273
rect 11152 6264 11204 6316
rect 12348 6400 12400 6452
rect 11612 6332 11664 6384
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 12256 6264 12308 6316
rect 12348 6264 12400 6316
rect 12532 6264 12584 6316
rect 15476 6400 15528 6452
rect 18236 6443 18288 6452
rect 13176 6375 13228 6384
rect 13176 6341 13185 6375
rect 13185 6341 13219 6375
rect 13219 6341 13228 6375
rect 13176 6332 13228 6341
rect 13912 6375 13964 6384
rect 13912 6341 13921 6375
rect 13921 6341 13955 6375
rect 13955 6341 13964 6375
rect 13912 6332 13964 6341
rect 13728 6307 13780 6316
rect 1584 6128 1636 6180
rect 5264 6128 5316 6180
rect 9680 6239 9732 6248
rect 9680 6205 9689 6239
rect 9689 6205 9723 6239
rect 9723 6205 9732 6239
rect 9680 6196 9732 6205
rect 13728 6273 13737 6307
rect 13737 6273 13771 6307
rect 13771 6273 13780 6307
rect 13728 6264 13780 6273
rect 14280 6264 14332 6316
rect 15108 6332 15160 6384
rect 15568 6332 15620 6384
rect 18236 6409 18245 6443
rect 18245 6409 18279 6443
rect 18279 6409 18288 6443
rect 18236 6400 18288 6409
rect 10140 6128 10192 6180
rect 1952 6060 2004 6112
rect 3792 6060 3844 6112
rect 5540 6060 5592 6112
rect 7656 6060 7708 6112
rect 10692 6128 10744 6180
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 14004 6196 14056 6248
rect 14740 6264 14792 6316
rect 14924 6307 14976 6316
rect 14924 6273 14933 6307
rect 14933 6273 14967 6307
rect 14967 6273 14976 6307
rect 14924 6264 14976 6273
rect 16212 6264 16264 6316
rect 16764 6264 16816 6316
rect 13360 6128 13412 6180
rect 15660 6196 15712 6248
rect 16488 6196 16540 6248
rect 11520 6103 11572 6112
rect 10508 6060 10560 6069
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 13728 6060 13780 6112
rect 14464 6060 14516 6112
rect 15568 6060 15620 6112
rect 3915 5958 3967 6010
rect 3979 5958 4031 6010
rect 4043 5958 4095 6010
rect 4107 5958 4159 6010
rect 4171 5958 4223 6010
rect 9846 5958 9898 6010
rect 9910 5958 9962 6010
rect 9974 5958 10026 6010
rect 10038 5958 10090 6010
rect 10102 5958 10154 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 15904 5958 15956 6010
rect 15968 5958 16020 6010
rect 16032 5958 16084 6010
rect 2964 5856 3016 5908
rect 3700 5856 3752 5908
rect 4528 5856 4580 5908
rect 10324 5899 10376 5908
rect 8852 5788 8904 5840
rect 9680 5788 9732 5840
rect 10324 5865 10333 5899
rect 10333 5865 10367 5899
rect 10367 5865 10376 5899
rect 10324 5856 10376 5865
rect 10692 5856 10744 5908
rect 10876 5856 10928 5908
rect 11888 5856 11940 5908
rect 12624 5856 12676 5908
rect 4344 5720 4396 5772
rect 5264 5763 5316 5772
rect 5264 5729 5273 5763
rect 5273 5729 5307 5763
rect 5307 5729 5316 5763
rect 5264 5720 5316 5729
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 1584 5652 1636 5704
rect 2596 5652 2648 5704
rect 4988 5652 5040 5704
rect 5540 5695 5592 5704
rect 5540 5661 5574 5695
rect 5574 5661 5592 5695
rect 5540 5652 5592 5661
rect 8392 5652 8444 5704
rect 10508 5720 10560 5772
rect 14648 5788 14700 5840
rect 7472 5584 7524 5636
rect 9680 5584 9732 5636
rect 9956 5627 10008 5636
rect 9956 5593 9965 5627
rect 9965 5593 9999 5627
rect 9999 5593 10008 5627
rect 9956 5584 10008 5593
rect 4344 5559 4396 5568
rect 4344 5525 4353 5559
rect 4353 5525 4387 5559
rect 4387 5525 4396 5559
rect 8300 5559 8352 5568
rect 4344 5516 4396 5525
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 8300 5516 8352 5525
rect 9864 5516 9916 5568
rect 10232 5584 10284 5636
rect 10692 5695 10744 5704
rect 10692 5661 10701 5695
rect 10701 5661 10735 5695
rect 10735 5661 10744 5695
rect 10692 5652 10744 5661
rect 12072 5720 12124 5772
rect 16948 5763 17000 5772
rect 16948 5729 16957 5763
rect 16957 5729 16991 5763
rect 16991 5729 17000 5763
rect 16948 5720 17000 5729
rect 10968 5695 11020 5704
rect 10968 5661 10985 5695
rect 10985 5661 11019 5695
rect 11019 5661 11020 5695
rect 10968 5652 11020 5661
rect 11152 5652 11204 5704
rect 11060 5584 11112 5636
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 13268 5695 13320 5704
rect 12440 5652 12492 5661
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 13728 5652 13780 5704
rect 13820 5652 13872 5704
rect 12164 5584 12216 5636
rect 14372 5652 14424 5704
rect 14832 5652 14884 5704
rect 16672 5652 16724 5704
rect 17132 5652 17184 5704
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 15108 5584 15160 5636
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 12624 5516 12676 5525
rect 13360 5559 13412 5568
rect 13360 5525 13369 5559
rect 13369 5525 13403 5559
rect 13403 5525 13412 5559
rect 13360 5516 13412 5525
rect 13728 5559 13780 5568
rect 13728 5525 13737 5559
rect 13737 5525 13771 5559
rect 13771 5525 13780 5559
rect 13728 5516 13780 5525
rect 15200 5516 15252 5568
rect 16212 5516 16264 5568
rect 16396 5559 16448 5568
rect 16396 5525 16405 5559
rect 16405 5525 16439 5559
rect 16439 5525 16448 5559
rect 16396 5516 16448 5525
rect 6880 5414 6932 5466
rect 6944 5414 6996 5466
rect 7008 5414 7060 5466
rect 7072 5414 7124 5466
rect 7136 5414 7188 5466
rect 12811 5414 12863 5466
rect 12875 5414 12927 5466
rect 12939 5414 12991 5466
rect 13003 5414 13055 5466
rect 13067 5414 13119 5466
rect 1400 5355 1452 5364
rect 1400 5321 1409 5355
rect 1409 5321 1443 5355
rect 1443 5321 1452 5355
rect 1400 5312 1452 5321
rect 2780 5312 2832 5364
rect 3056 5312 3108 5364
rect 4344 5312 4396 5364
rect 5448 5312 5500 5364
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 2964 5244 3016 5296
rect 3700 5176 3752 5228
rect 5356 5176 5408 5228
rect 3148 5108 3200 5160
rect 1584 5040 1636 5092
rect 5448 5108 5500 5160
rect 8300 5312 8352 5364
rect 11060 5312 11112 5364
rect 11980 5312 12032 5364
rect 13360 5312 13412 5364
rect 15108 5355 15160 5364
rect 15108 5321 15117 5355
rect 15117 5321 15151 5355
rect 15151 5321 15160 5355
rect 15108 5312 15160 5321
rect 16672 5312 16724 5364
rect 9864 5244 9916 5296
rect 10508 5244 10560 5296
rect 7564 5219 7616 5228
rect 6736 5108 6788 5160
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 7564 5176 7616 5185
rect 9772 5176 9824 5228
rect 10232 5176 10284 5228
rect 11520 5244 11572 5296
rect 11796 5244 11848 5296
rect 11336 5176 11388 5228
rect 12164 5219 12216 5228
rect 7288 5108 7340 5160
rect 11152 5108 11204 5160
rect 12164 5185 12173 5219
rect 12173 5185 12207 5219
rect 12207 5185 12216 5219
rect 12164 5176 12216 5185
rect 12256 5176 12308 5228
rect 14188 5176 14240 5228
rect 14372 5219 14424 5228
rect 14372 5185 14381 5219
rect 14381 5185 14415 5219
rect 14415 5185 14424 5219
rect 14372 5176 14424 5185
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 14648 5219 14700 5228
rect 14648 5185 14657 5219
rect 14657 5185 14691 5219
rect 14691 5185 14700 5219
rect 14648 5176 14700 5185
rect 15568 5219 15620 5228
rect 4988 5083 5040 5092
rect 4988 5049 4997 5083
rect 4997 5049 5031 5083
rect 5031 5049 5040 5083
rect 4988 5040 5040 5049
rect 7748 5040 7800 5092
rect 14096 5108 14148 5160
rect 15200 5108 15252 5160
rect 2412 5015 2464 5024
rect 2412 4981 2421 5015
rect 2421 4981 2455 5015
rect 2455 4981 2464 5015
rect 2412 4972 2464 4981
rect 6276 4972 6328 5024
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 9680 4972 9732 5024
rect 10416 5015 10468 5024
rect 10416 4981 10425 5015
rect 10425 4981 10459 5015
rect 10459 4981 10468 5015
rect 10416 4972 10468 4981
rect 14188 5040 14240 5092
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 14096 4972 14148 5024
rect 14464 4972 14516 5024
rect 16764 5176 16816 5228
rect 16948 5219 17000 5228
rect 16948 5185 16982 5219
rect 16982 5185 17000 5219
rect 16948 5176 17000 5185
rect 16120 4972 16172 5024
rect 3915 4870 3967 4922
rect 3979 4870 4031 4922
rect 4043 4870 4095 4922
rect 4107 4870 4159 4922
rect 4171 4870 4223 4922
rect 9846 4870 9898 4922
rect 9910 4870 9962 4922
rect 9974 4870 10026 4922
rect 10038 4870 10090 4922
rect 10102 4870 10154 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 15904 4870 15956 4922
rect 15968 4870 16020 4922
rect 16032 4870 16084 4922
rect 3056 4811 3108 4820
rect 3056 4777 3065 4811
rect 3065 4777 3099 4811
rect 3099 4777 3108 4811
rect 3056 4768 3108 4777
rect 3700 4768 3752 4820
rect 7472 4768 7524 4820
rect 7748 4768 7800 4820
rect 11796 4768 11848 4820
rect 12440 4768 12492 4820
rect 16212 4768 16264 4820
rect 9496 4743 9548 4752
rect 9496 4709 9505 4743
rect 9505 4709 9539 4743
rect 9539 4709 9548 4743
rect 9496 4700 9548 4709
rect 1584 4632 1636 4684
rect 5448 4632 5500 4684
rect 6552 4632 6604 4684
rect 9128 4675 9180 4684
rect 9128 4641 9137 4675
rect 9137 4641 9171 4675
rect 9171 4641 9180 4675
rect 9128 4632 9180 4641
rect 3792 4564 3844 4616
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 7196 4564 7248 4616
rect 7380 4607 7432 4616
rect 7380 4573 7414 4607
rect 7414 4573 7432 4607
rect 7380 4564 7432 4573
rect 11336 4632 11388 4684
rect 11428 4632 11480 4684
rect 10600 4607 10652 4616
rect 10600 4573 10609 4607
rect 10609 4573 10643 4607
rect 10643 4573 10652 4607
rect 10600 4564 10652 4573
rect 1676 4496 1728 4548
rect 2320 4428 2372 4480
rect 10508 4496 10560 4548
rect 4896 4428 4948 4480
rect 8484 4471 8536 4480
rect 8484 4437 8493 4471
rect 8493 4437 8527 4471
rect 8527 4437 8536 4471
rect 11980 4564 12032 4616
rect 14464 4564 14516 4616
rect 14004 4496 14056 4548
rect 8484 4428 8536 4437
rect 11888 4428 11940 4480
rect 12072 4471 12124 4480
rect 12072 4437 12081 4471
rect 12081 4437 12115 4471
rect 12115 4437 12124 4471
rect 12072 4428 12124 4437
rect 13820 4428 13872 4480
rect 14924 4496 14976 4548
rect 15660 4564 15712 4616
rect 16028 4564 16080 4616
rect 16396 4607 16448 4616
rect 16396 4573 16405 4607
rect 16405 4573 16439 4607
rect 16439 4573 16448 4607
rect 16396 4564 16448 4573
rect 16580 4564 16632 4616
rect 16764 4496 16816 4548
rect 17316 4496 17368 4548
rect 16672 4428 16724 4480
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 18328 4428 18380 4437
rect 6880 4326 6932 4378
rect 6944 4326 6996 4378
rect 7008 4326 7060 4378
rect 7072 4326 7124 4378
rect 7136 4326 7188 4378
rect 12811 4326 12863 4378
rect 12875 4326 12927 4378
rect 12939 4326 12991 4378
rect 13003 4326 13055 4378
rect 13067 4326 13119 4378
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 3056 4224 3108 4276
rect 8484 4224 8536 4276
rect 10968 4224 11020 4276
rect 12256 4267 12308 4276
rect 12256 4233 12265 4267
rect 12265 4233 12299 4267
rect 12299 4233 12308 4267
rect 12256 4224 12308 4233
rect 7288 4156 7340 4208
rect 2412 4088 2464 4140
rect 1768 4020 1820 4072
rect 2504 4020 2556 4072
rect 2780 4020 2832 4072
rect 3424 4063 3476 4072
rect 3424 4029 3433 4063
rect 3433 4029 3467 4063
rect 3467 4029 3476 4063
rect 3424 4020 3476 4029
rect 3608 4020 3660 4072
rect 4252 4088 4304 4140
rect 4896 4131 4948 4140
rect 4896 4097 4930 4131
rect 4930 4097 4948 4131
rect 4896 4088 4948 4097
rect 5356 4088 5408 4140
rect 7748 4131 7800 4140
rect 4528 4020 4580 4072
rect 7196 4063 7248 4072
rect 2044 3952 2096 4004
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 8944 4088 8996 4140
rect 9588 4088 9640 4140
rect 9772 4088 9824 4140
rect 5632 3952 5684 4004
rect 2688 3884 2740 3936
rect 4344 3927 4396 3936
rect 4344 3893 4353 3927
rect 4353 3893 4387 3927
rect 4387 3893 4396 3927
rect 4344 3884 4396 3893
rect 6920 3884 6972 3936
rect 10232 3952 10284 4004
rect 10416 4088 10468 4140
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 11244 4088 11296 4140
rect 11520 4020 11572 4072
rect 10784 3952 10836 4004
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 12624 4088 12676 4140
rect 14004 4156 14056 4208
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 16948 4224 17000 4276
rect 17316 4267 17368 4276
rect 17316 4233 17325 4267
rect 17325 4233 17359 4267
rect 17359 4233 17368 4267
rect 17316 4224 17368 4233
rect 16028 4156 16080 4208
rect 16304 4199 16356 4208
rect 16304 4165 16313 4199
rect 16313 4165 16347 4199
rect 16347 4165 16356 4199
rect 16304 4156 16356 4165
rect 14280 4131 14332 4140
rect 11980 4063 12032 4072
rect 11980 4029 11989 4063
rect 11989 4029 12023 4063
rect 12023 4029 12032 4063
rect 11980 4020 12032 4029
rect 11796 3952 11848 4004
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 17408 4088 17460 4140
rect 17684 4131 17736 4140
rect 17684 4097 17693 4131
rect 17693 4097 17727 4131
rect 17727 4097 17736 4131
rect 17684 4088 17736 4097
rect 18328 4088 18380 4140
rect 16856 4020 16908 4072
rect 17776 4063 17828 4072
rect 17776 4029 17785 4063
rect 17785 4029 17819 4063
rect 17819 4029 17828 4063
rect 17776 4020 17828 4029
rect 12900 3995 12952 4004
rect 12900 3961 12909 3995
rect 12909 3961 12943 3995
rect 12943 3961 12952 3995
rect 12900 3952 12952 3961
rect 15660 3952 15712 4004
rect 16120 3952 16172 4004
rect 18236 3995 18288 4004
rect 9036 3884 9088 3936
rect 9220 3884 9272 3936
rect 11428 3884 11480 3936
rect 12716 3884 12768 3936
rect 13176 3884 13228 3936
rect 14372 3884 14424 3936
rect 14556 3884 14608 3936
rect 14924 3927 14976 3936
rect 14924 3893 14933 3927
rect 14933 3893 14967 3927
rect 14967 3893 14976 3927
rect 14924 3884 14976 3893
rect 18236 3961 18245 3995
rect 18245 3961 18279 3995
rect 18279 3961 18288 3995
rect 18236 3952 18288 3961
rect 18696 3884 18748 3936
rect 3915 3782 3967 3834
rect 3979 3782 4031 3834
rect 4043 3782 4095 3834
rect 4107 3782 4159 3834
rect 4171 3782 4223 3834
rect 9846 3782 9898 3834
rect 9910 3782 9962 3834
rect 9974 3782 10026 3834
rect 10038 3782 10090 3834
rect 10102 3782 10154 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 15904 3782 15956 3834
rect 15968 3782 16020 3834
rect 16032 3782 16084 3834
rect 2412 3680 2464 3732
rect 3608 3680 3660 3732
rect 4252 3680 4304 3732
rect 5080 3680 5132 3732
rect 7564 3680 7616 3732
rect 8944 3723 8996 3732
rect 8944 3689 8953 3723
rect 8953 3689 8987 3723
rect 8987 3689 8996 3723
rect 8944 3680 8996 3689
rect 1584 3612 1636 3664
rect 3424 3655 3476 3664
rect 3424 3621 3433 3655
rect 3433 3621 3467 3655
rect 3467 3621 3476 3655
rect 3424 3612 3476 3621
rect 2044 3587 2096 3596
rect 2044 3553 2053 3587
rect 2053 3553 2087 3587
rect 2087 3553 2096 3587
rect 2044 3544 2096 3553
rect 2780 3476 2832 3528
rect 3240 3476 3292 3528
rect 5540 3612 5592 3664
rect 5724 3612 5776 3664
rect 6644 3612 6696 3664
rect 11796 3680 11848 3732
rect 11980 3723 12032 3732
rect 11980 3689 11989 3723
rect 11989 3689 12023 3723
rect 12023 3689 12032 3723
rect 11980 3680 12032 3689
rect 14280 3680 14332 3732
rect 14372 3680 14424 3732
rect 16856 3723 16908 3732
rect 12164 3612 12216 3664
rect 4620 3544 4672 3596
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 6552 3544 6604 3596
rect 9128 3544 9180 3596
rect 6920 3519 6972 3528
rect 6920 3485 6929 3519
rect 6929 3485 6963 3519
rect 6963 3485 6972 3519
rect 6920 3476 6972 3485
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 13176 3544 13228 3596
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 9588 3519 9640 3528
rect 9588 3485 9597 3519
rect 9597 3485 9631 3519
rect 9631 3485 9640 3519
rect 9588 3476 9640 3485
rect 11428 3519 11480 3528
rect 11428 3485 11446 3519
rect 11446 3485 11480 3519
rect 11428 3476 11480 3485
rect 12900 3519 12952 3528
rect 3148 3408 3200 3460
rect 10140 3408 10192 3460
rect 10968 3408 11020 3460
rect 5632 3340 5684 3392
rect 6092 3383 6144 3392
rect 6092 3349 6101 3383
rect 6101 3349 6135 3383
rect 6135 3349 6144 3383
rect 6092 3340 6144 3349
rect 10232 3340 10284 3392
rect 11060 3340 11112 3392
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 12440 3408 12492 3460
rect 13452 3408 13504 3460
rect 13636 3476 13688 3528
rect 13820 3476 13872 3528
rect 16120 3476 16172 3528
rect 16856 3689 16865 3723
rect 16865 3689 16899 3723
rect 16899 3689 16908 3723
rect 16856 3680 16908 3689
rect 17776 3723 17828 3732
rect 17776 3689 17785 3723
rect 17785 3689 17819 3723
rect 17819 3689 17828 3723
rect 17776 3680 17828 3689
rect 16488 3655 16540 3664
rect 16488 3621 16497 3655
rect 16497 3621 16531 3655
rect 16531 3621 16540 3655
rect 16488 3612 16540 3621
rect 18328 3544 18380 3596
rect 17040 3519 17092 3528
rect 17040 3485 17049 3519
rect 17049 3485 17083 3519
rect 17083 3485 17092 3519
rect 17040 3476 17092 3485
rect 17132 3519 17184 3528
rect 17132 3485 17141 3519
rect 17141 3485 17175 3519
rect 17175 3485 17184 3519
rect 17132 3476 17184 3485
rect 13912 3408 13964 3460
rect 14464 3451 14516 3460
rect 14464 3417 14473 3451
rect 14473 3417 14507 3451
rect 14507 3417 14516 3451
rect 14464 3408 14516 3417
rect 14648 3408 14700 3460
rect 15108 3383 15160 3392
rect 15108 3349 15117 3383
rect 15117 3349 15151 3383
rect 15151 3349 15160 3383
rect 15108 3340 15160 3349
rect 6880 3238 6932 3290
rect 6944 3238 6996 3290
rect 7008 3238 7060 3290
rect 7072 3238 7124 3290
rect 7136 3238 7188 3290
rect 12811 3238 12863 3290
rect 12875 3238 12927 3290
rect 12939 3238 12991 3290
rect 13003 3238 13055 3290
rect 13067 3238 13119 3290
rect 3148 3179 3200 3188
rect 3148 3145 3157 3179
rect 3157 3145 3191 3179
rect 3191 3145 3200 3179
rect 3148 3136 3200 3145
rect 2044 3068 2096 3120
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 2688 3043 2740 3052
rect 2688 3009 2697 3043
rect 2697 3009 2731 3043
rect 2731 3009 2740 3043
rect 2688 3000 2740 3009
rect 4620 3068 4672 3120
rect 7104 3068 7156 3120
rect 7840 3068 7892 3120
rect 4252 3043 4304 3052
rect 4252 3009 4286 3043
rect 4286 3009 4304 3043
rect 5724 3043 5776 3052
rect 4252 3000 4304 3009
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 6552 3000 6604 3052
rect 7748 3043 7800 3052
rect 7748 3009 7757 3043
rect 7757 3009 7791 3043
rect 7791 3009 7800 3043
rect 7748 3000 7800 3009
rect 9220 3136 9272 3188
rect 9588 3136 9640 3188
rect 10140 3136 10192 3188
rect 14004 3136 14056 3188
rect 15200 3136 15252 3188
rect 15384 3136 15436 3188
rect 17132 3136 17184 3188
rect 9036 3068 9088 3120
rect 9128 3000 9180 3052
rect 9404 3068 9456 3120
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 12164 3068 12216 3120
rect 12440 3000 12492 3052
rect 12716 3043 12768 3052
rect 14280 3068 14332 3120
rect 12716 3009 12734 3043
rect 12734 3009 12768 3043
rect 12716 3000 12768 3009
rect 13636 3000 13688 3052
rect 15108 3068 15160 3120
rect 16304 3068 16356 3120
rect 16580 3000 16632 3052
rect 16764 3000 16816 3052
rect 2044 2932 2096 2984
rect 2228 2975 2280 2984
rect 2228 2941 2237 2975
rect 2237 2941 2271 2975
rect 2271 2941 2280 2975
rect 2228 2932 2280 2941
rect 13176 2932 13228 2984
rect 5540 2864 5592 2916
rect 6736 2864 6788 2916
rect 7840 2864 7892 2916
rect 7380 2796 7432 2848
rect 11612 2839 11664 2848
rect 11612 2805 11621 2839
rect 11621 2805 11655 2839
rect 11655 2805 11664 2839
rect 11612 2796 11664 2805
rect 12624 2796 12676 2848
rect 13360 2839 13412 2848
rect 13360 2805 13369 2839
rect 13369 2805 13403 2839
rect 13403 2805 13412 2839
rect 13360 2796 13412 2805
rect 3915 2694 3967 2746
rect 3979 2694 4031 2746
rect 4043 2694 4095 2746
rect 4107 2694 4159 2746
rect 4171 2694 4223 2746
rect 9846 2694 9898 2746
rect 9910 2694 9962 2746
rect 9974 2694 10026 2746
rect 10038 2694 10090 2746
rect 10102 2694 10154 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 15904 2694 15956 2746
rect 15968 2694 16020 2746
rect 16032 2694 16084 2746
rect 3424 2592 3476 2644
rect 9312 2592 9364 2644
rect 11152 2592 11204 2644
rect 12716 2592 12768 2644
rect 13820 2592 13872 2644
rect 14648 2592 14700 2644
rect 4252 2524 4304 2576
rect 6552 2567 6604 2576
rect 6552 2533 6561 2567
rect 6561 2533 6595 2567
rect 6595 2533 6604 2567
rect 6552 2524 6604 2533
rect 1308 2456 1360 2508
rect 2320 2456 2372 2508
rect 8852 2524 8904 2576
rect 9128 2567 9180 2576
rect 9128 2533 9137 2567
rect 9137 2533 9171 2567
rect 9171 2533 9180 2567
rect 9128 2524 9180 2533
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 9588 2499 9640 2508
rect 9588 2465 9597 2499
rect 9597 2465 9631 2499
rect 9631 2465 9640 2499
rect 9588 2456 9640 2465
rect 11704 2524 11756 2576
rect 1952 2431 2004 2440
rect 1952 2397 1961 2431
rect 1961 2397 1995 2431
rect 1995 2397 2004 2431
rect 1952 2388 2004 2397
rect 2780 2388 2832 2440
rect 3884 2388 3936 2440
rect 4344 2388 4396 2440
rect 5540 2388 5592 2440
rect 6092 2388 6144 2440
rect 6736 2388 6788 2440
rect 7288 2388 7340 2440
rect 9036 2388 9088 2440
rect 9404 2388 9456 2440
rect 9496 2431 9548 2440
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 6460 2320 6512 2372
rect 10324 2388 10376 2440
rect 10232 2320 10284 2372
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11612 2456 11664 2508
rect 13176 2524 13228 2576
rect 15476 2524 15528 2576
rect 13912 2456 13964 2508
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 12624 2431 12676 2440
rect 11152 2388 11204 2397
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 13452 2388 13504 2440
rect 14556 2431 14608 2440
rect 14556 2397 14590 2431
rect 14590 2397 14608 2431
rect 14556 2388 14608 2397
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 17684 2388 17736 2440
rect 12716 2320 12768 2372
rect 13728 2320 13780 2372
rect 2044 2252 2096 2304
rect 7656 2252 7708 2304
rect 7748 2252 7800 2304
rect 11520 2252 11572 2304
rect 11980 2295 12032 2304
rect 11980 2261 11989 2295
rect 11989 2261 12023 2295
rect 12023 2261 12032 2295
rect 11980 2252 12032 2261
rect 16764 2252 16816 2304
rect 18052 2252 18104 2304
rect 6880 2150 6932 2202
rect 6944 2150 6996 2202
rect 7008 2150 7060 2202
rect 7072 2150 7124 2202
rect 7136 2150 7188 2202
rect 12811 2150 12863 2202
rect 12875 2150 12927 2202
rect 12939 2150 12991 2202
rect 13003 2150 13055 2202
rect 13067 2150 13119 2202
rect 1952 2048 2004 2100
rect 7472 2048 7524 2100
rect 7656 2048 7708 2100
rect 11980 2048 12032 2100
rect 9496 1980 9548 2032
rect 14188 1980 14240 2032
<< metal2 >>
rect 18 19200 74 20000
rect 1306 19200 1362 20000
rect 1950 19200 2006 20000
rect 2594 19200 2650 20000
rect 3882 19200 3938 20000
rect 4526 19200 4582 20000
rect 5170 19200 5226 20000
rect 6458 19200 6514 20000
rect 7102 19200 7158 20000
rect 7746 19200 7802 20000
rect 9034 19200 9090 20000
rect 9678 19200 9734 20000
rect 10322 19200 10378 20000
rect 11610 19200 11666 20000
rect 12254 19200 12310 20000
rect 12898 19200 12954 20000
rect 13004 19230 13216 19258
rect 32 16590 60 19200
rect 1320 17202 1348 19200
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2226 17776 2282 17785
rect 2226 17711 2282 17720
rect 1308 17196 1360 17202
rect 1308 17138 1360 17144
rect 1398 17096 1454 17105
rect 1398 17031 1454 17040
rect 20 16584 72 16590
rect 20 16526 72 16532
rect 1412 16114 1440 17031
rect 2240 16522 2268 17711
rect 2504 16720 2556 16726
rect 2504 16662 2556 16668
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2228 16516 2280 16522
rect 2228 16458 2280 16464
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 16250 1992 16390
rect 2240 16250 2268 16458
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1768 15972 1820 15978
rect 1768 15914 1820 15920
rect 1780 15434 1808 15914
rect 1768 15428 1820 15434
rect 1768 15370 1820 15376
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1398 15056 1454 15065
rect 1398 14991 1400 15000
rect 1452 14991 1454 15000
rect 1400 14962 1452 14968
rect 1872 14958 1900 15370
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 1400 14408 1452 14414
rect 1398 14376 1400 14385
rect 1452 14376 1454 14385
rect 1398 14311 1454 14320
rect 1872 13326 1900 14894
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1768 12232 1820 12238
rect 1872 12186 1900 13262
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1964 12238 1992 12582
rect 2424 12424 2452 16594
rect 2240 12396 2452 12424
rect 1820 12180 1900 12186
rect 1768 12174 1900 12180
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1780 12158 1900 12174
rect 1872 11762 1900 12158
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1398 11656 1454 11665
rect 1398 11591 1400 11600
rect 1452 11591 1454 11600
rect 1400 11562 1452 11568
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1872 10674 1900 11698
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2056 10266 2084 10610
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9625 1440 9998
rect 1398 9616 1454 9625
rect 2148 9586 2176 11154
rect 1398 9551 1454 9560
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1584 8968 1636 8974
rect 1490 8936 1546 8945
rect 1584 8910 1636 8916
rect 1490 8871 1546 8880
rect 1504 8634 1532 8871
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1596 8362 1624 8910
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 7410 1624 8298
rect 2240 8294 2268 12396
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2332 10062 2360 10950
rect 2424 10266 2452 11086
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2332 8634 2360 9522
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1964 7478 1992 7686
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1398 6896 1454 6905
rect 1398 6831 1400 6840
rect 1452 6831 1454 6840
rect 1400 6802 1452 6808
rect 1400 6248 1452 6254
rect 1398 6216 1400 6225
rect 1452 6216 1454 6225
rect 1596 6186 1624 7346
rect 2056 7002 2084 7822
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1398 6151 1454 6160
rect 1584 6180 1636 6186
rect 1412 5370 1440 6151
rect 1584 6122 1636 6128
rect 1596 5710 1624 6122
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1596 5098 1624 5646
rect 1780 5234 1808 6802
rect 2148 6798 2176 7686
rect 2516 6905 2544 16662
rect 2792 16454 2820 19071
rect 7116 17626 7144 19200
rect 7116 17598 7328 17626
rect 6880 17436 7188 17456
rect 6880 17434 6886 17436
rect 6942 17434 6966 17436
rect 7022 17434 7046 17436
rect 7102 17434 7126 17436
rect 7182 17434 7188 17436
rect 6942 17382 6944 17434
rect 7124 17382 7126 17434
rect 6880 17380 6886 17382
rect 6942 17380 6966 17382
rect 7022 17380 7046 17382
rect 7102 17380 7126 17382
rect 7182 17380 7188 17382
rect 6880 17360 7188 17380
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2884 16794 2912 17138
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2976 16590 3004 16934
rect 3915 16892 4223 16912
rect 3915 16890 3921 16892
rect 3977 16890 4001 16892
rect 4057 16890 4081 16892
rect 4137 16890 4161 16892
rect 4217 16890 4223 16892
rect 3977 16838 3979 16890
rect 4159 16838 4161 16890
rect 3915 16836 3921 16838
rect 3977 16836 4001 16838
rect 4057 16836 4081 16838
rect 4137 16836 4161 16838
rect 4217 16836 4223 16838
rect 3915 16816 4223 16836
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2792 15706 2820 16050
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 3160 15570 3188 16662
rect 4356 16590 4384 17274
rect 7300 17202 7328 17598
rect 7760 17338 7788 19200
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 9048 17202 9076 19200
rect 9692 17338 9720 19200
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 3344 16114 3372 16458
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3344 15706 3372 16050
rect 3528 16046 3556 16186
rect 3608 16176 3660 16182
rect 3608 16118 3660 16124
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 3436 15502 3464 15914
rect 3620 15706 3648 16118
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3712 14958 3740 16186
rect 3804 16046 3832 16390
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3804 15688 3832 15982
rect 3915 15804 4223 15824
rect 3915 15802 3921 15804
rect 3977 15802 4001 15804
rect 4057 15802 4081 15804
rect 4137 15802 4161 15804
rect 4217 15802 4223 15804
rect 3977 15750 3979 15802
rect 4159 15750 4161 15802
rect 3915 15748 3921 15750
rect 3977 15748 4001 15750
rect 4057 15748 4081 15750
rect 4137 15748 4161 15750
rect 4217 15748 4223 15750
rect 3915 15728 4223 15748
rect 3804 15660 3924 15688
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3804 15162 3832 15506
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14482 3740 14894
rect 3896 14890 3924 15660
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4080 14958 4108 15370
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3915 14716 4223 14736
rect 3915 14714 3921 14716
rect 3977 14714 4001 14716
rect 4057 14714 4081 14716
rect 4137 14714 4161 14716
rect 4217 14714 4223 14716
rect 3977 14662 3979 14714
rect 4159 14662 4161 14714
rect 3915 14660 3921 14662
rect 3977 14660 4001 14662
rect 4057 14660 4081 14662
rect 4137 14660 4161 14662
rect 4217 14660 4223 14662
rect 3915 14640 4223 14660
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 4264 14414 4292 16050
rect 5184 15570 5212 16526
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5276 15706 5304 15846
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4356 14346 4384 15438
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 14618 4936 14758
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4344 14340 4396 14346
rect 4344 14282 4396 14288
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 5000 13938 5028 14282
rect 5184 14006 5212 15506
rect 5356 15496 5408 15502
rect 5460 15484 5488 15982
rect 5552 15502 5580 16390
rect 6380 16250 6408 16526
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 5644 16114 5672 16186
rect 6564 16182 6592 17138
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6656 16454 6684 17070
rect 6748 16794 6776 17138
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6552 16176 6604 16182
rect 6552 16118 6604 16124
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5408 15456 5488 15484
rect 5540 15496 5592 15502
rect 5356 15438 5408 15444
rect 5540 15438 5592 15444
rect 5632 15088 5684 15094
rect 5684 15048 5764 15076
rect 5632 15030 5684 15036
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5276 14278 5304 14894
rect 5552 14346 5580 14894
rect 5736 14618 5764 15048
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6288 14618 6316 14894
rect 6564 14822 6592 16118
rect 6656 16114 6684 16390
rect 6748 16182 6776 16730
rect 7208 16697 7236 16934
rect 7748 16720 7800 16726
rect 7194 16688 7250 16697
rect 7194 16623 7250 16632
rect 7484 16680 7748 16708
rect 7484 16522 7512 16680
rect 7748 16662 7800 16668
rect 7944 16590 7972 17002
rect 9048 16794 9076 17138
rect 10336 17134 10364 19200
rect 12268 17252 12296 19200
rect 12912 19122 12940 19200
rect 13004 19122 13032 19230
rect 12912 19094 13032 19122
rect 12811 17436 13119 17456
rect 12811 17434 12817 17436
rect 12873 17434 12897 17436
rect 12953 17434 12977 17436
rect 13033 17434 13057 17436
rect 13113 17434 13119 17436
rect 12873 17382 12875 17434
rect 13055 17382 13057 17434
rect 12811 17380 12817 17382
rect 12873 17380 12897 17382
rect 12953 17380 12977 17382
rect 13033 17380 13057 17382
rect 13113 17380 13119 17382
rect 12811 17360 13119 17380
rect 12440 17264 12492 17270
rect 12268 17224 12440 17252
rect 12440 17206 12492 17212
rect 13188 17202 13216 19230
rect 14186 19200 14242 20000
rect 14830 19200 14886 20000
rect 15474 19200 15530 20000
rect 16762 19200 16818 20000
rect 17406 19200 17462 20000
rect 18050 19200 18106 20000
rect 19338 19200 19394 20000
rect 14200 17338 14228 19200
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 7472 16516 7524 16522
rect 7472 16458 7524 16464
rect 6880 16348 7188 16368
rect 6880 16346 6886 16348
rect 6942 16346 6966 16348
rect 7022 16346 7046 16348
rect 7102 16346 7126 16348
rect 7182 16346 7188 16348
rect 6942 16294 6944 16346
rect 7124 16294 7126 16346
rect 6880 16292 6886 16294
rect 6942 16292 6966 16294
rect 7022 16292 7046 16294
rect 7102 16292 7126 16294
rect 7182 16292 7188 16294
rect 6880 16272 7188 16292
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 7576 16114 7604 16526
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 7208 15706 7236 16050
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 6880 15260 7188 15280
rect 6880 15258 6886 15260
rect 6942 15258 6966 15260
rect 7022 15258 7046 15260
rect 7102 15258 7126 15260
rect 7182 15258 7188 15260
rect 6942 15206 6944 15258
rect 7124 15206 7126 15258
rect 6880 15204 6886 15206
rect 6942 15204 6966 15206
rect 7022 15204 7046 15206
rect 7102 15204 7126 15206
rect 7182 15204 7188 15206
rect 6880 15184 7188 15204
rect 7300 15026 7328 15846
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 15026 7512 15302
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7012 14952 7064 14958
rect 6932 14912 7012 14940
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 5736 14414 5764 14554
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 3620 13530 3648 13874
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 3915 13628 4223 13648
rect 3915 13626 3921 13628
rect 3977 13626 4001 13628
rect 4057 13626 4081 13628
rect 4137 13626 4161 13628
rect 4217 13626 4223 13628
rect 3977 13574 3979 13626
rect 4159 13574 4161 13626
rect 3915 13572 3921 13574
rect 3977 13572 4001 13574
rect 4057 13572 4081 13574
rect 4137 13572 4161 13574
rect 4217 13572 4223 13574
rect 3915 13552 4223 13572
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 2596 13252 2648 13258
rect 2596 13194 2648 13200
rect 2608 12986 2636 13194
rect 3804 12986 3832 13262
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 11830 3096 12582
rect 3712 12442 3740 12650
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3252 11354 3280 11494
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3712 11082 3740 12038
rect 3804 11694 3832 12922
rect 4264 12646 4292 13126
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 3915 12540 4223 12560
rect 3915 12538 3921 12540
rect 3977 12538 4001 12540
rect 4057 12538 4081 12540
rect 4137 12538 4161 12540
rect 4217 12538 4223 12540
rect 3977 12486 3979 12538
rect 4159 12486 4161 12538
rect 3915 12484 3921 12486
rect 3977 12484 4001 12486
rect 4057 12484 4081 12486
rect 4137 12484 4161 12486
rect 4217 12484 4223 12486
rect 3915 12464 4223 12484
rect 4264 12238 4292 12582
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3804 10742 3832 11630
rect 3915 11452 4223 11472
rect 3915 11450 3921 11452
rect 3977 11450 4001 11452
rect 4057 11450 4081 11452
rect 4137 11450 4161 11452
rect 4217 11450 4223 11452
rect 3977 11398 3979 11450
rect 4159 11398 4161 11450
rect 3915 11396 3921 11398
rect 3977 11396 4001 11398
rect 4057 11396 4081 11398
rect 4137 11396 4161 11398
rect 4217 11396 4223 11398
rect 3915 11376 4223 11396
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 4172 10674 4200 11222
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2884 9994 2912 10406
rect 3915 10364 4223 10384
rect 3915 10362 3921 10364
rect 3977 10362 4001 10364
rect 4057 10362 4081 10364
rect 4137 10362 4161 10364
rect 4217 10362 4223 10364
rect 3977 10310 3979 10362
rect 4159 10310 4161 10362
rect 3915 10308 3921 10310
rect 3977 10308 4001 10310
rect 4057 10308 4081 10310
rect 4137 10308 4161 10310
rect 4217 10308 4223 10310
rect 3915 10288 4223 10308
rect 3054 10160 3110 10169
rect 3054 10095 3110 10104
rect 3148 10124 3200 10130
rect 3068 10062 3096 10095
rect 3148 10066 3200 10072
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 8974 2820 9318
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2884 8906 2912 9930
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8430 2820 8774
rect 2884 8634 2912 8842
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3160 8430 3188 10066
rect 4356 10062 4384 13806
rect 4540 13326 4568 13874
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 13326 4752 13670
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 5184 12986 5212 13942
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 5276 13530 5304 13738
rect 5552 13734 5580 14282
rect 5736 13938 5764 14350
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5368 13326 5396 13466
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 5000 12434 5028 12786
rect 5276 12782 5304 13194
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5276 12646 5304 12718
rect 5368 12714 5396 13262
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5460 12646 5488 13262
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5552 12850 5580 13126
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5000 12406 5120 12434
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4540 10062 4568 12310
rect 5092 12238 5120 12406
rect 5276 12306 5304 12582
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 5000 11082 5028 11562
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 5092 10810 5120 12174
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 11286 5212 11494
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 5368 11218 5396 12378
rect 5460 12238 5488 12582
rect 5552 12442 5580 12582
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5644 12170 5672 12854
rect 5736 12850 5764 13874
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5736 12442 5764 12650
rect 5828 12646 5856 14282
rect 6012 14074 6040 14282
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6104 13530 6132 13942
rect 6564 13734 6592 14758
rect 6656 13734 6684 14758
rect 6734 14648 6790 14657
rect 6734 14583 6790 14592
rect 6748 14414 6776 14583
rect 6932 14550 6960 14912
rect 7012 14894 7064 14900
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7102 14784 7158 14793
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 7024 14414 7052 14758
rect 7102 14719 7158 14728
rect 6736 14408 6788 14414
rect 7012 14408 7064 14414
rect 6736 14350 6788 14356
rect 7010 14376 7012 14385
rect 7064 14376 7066 14385
rect 7116 14346 7144 14719
rect 7380 14544 7432 14550
rect 7286 14512 7342 14521
rect 7380 14486 7432 14492
rect 7286 14447 7288 14456
rect 7340 14447 7342 14456
rect 7288 14418 7340 14424
rect 7010 14311 7066 14320
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 6880 14172 7188 14192
rect 6880 14170 6886 14172
rect 6942 14170 6966 14172
rect 7022 14170 7046 14172
rect 7102 14170 7126 14172
rect 7182 14170 7188 14172
rect 6942 14118 6944 14170
rect 7124 14118 7126 14170
rect 6880 14116 6886 14118
rect 6942 14116 6966 14118
rect 7022 14116 7046 14118
rect 7102 14116 7126 14118
rect 7182 14116 7188 14118
rect 6880 14096 7188 14116
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6092 13524 6144 13530
rect 7300 13512 7328 14214
rect 7392 14074 7420 14486
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7392 13530 7420 14010
rect 7484 13938 7512 14214
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 6092 13466 6144 13472
rect 7208 13484 7328 13512
rect 7380 13524 7432 13530
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5816 12164 5868 12170
rect 5816 12106 5868 12112
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5552 11150 5580 12038
rect 5828 11898 5856 12106
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5920 11354 5948 11834
rect 6104 11694 6132 13466
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6288 11830 6316 12378
rect 6748 12374 6776 13194
rect 7208 13172 7236 13484
rect 7380 13466 7432 13472
rect 7288 13184 7340 13190
rect 7208 13144 7288 13172
rect 7288 13126 7340 13132
rect 6880 13084 7188 13104
rect 6880 13082 6886 13084
rect 6942 13082 6966 13084
rect 7022 13082 7046 13084
rect 7102 13082 7126 13084
rect 7182 13082 7188 13084
rect 6942 13030 6944 13082
rect 7124 13030 7126 13082
rect 6880 13028 6886 13030
rect 6942 13028 6966 13030
rect 7022 13028 7046 13030
rect 7102 13028 7126 13030
rect 7182 13028 7188 13030
rect 6880 13008 7188 13028
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7208 12442 7236 12786
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 7300 12306 7328 13126
rect 7576 12918 7604 16050
rect 7654 16008 7710 16017
rect 7654 15943 7710 15952
rect 7668 15502 7696 15943
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7840 15632 7892 15638
rect 7840 15574 7892 15580
rect 7656 15496 7708 15502
rect 7708 15456 7788 15484
rect 7656 15438 7708 15444
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7564 12912 7616 12918
rect 7564 12854 7616 12860
rect 7576 12442 7604 12854
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 6880 11996 7188 12016
rect 6880 11994 6886 11996
rect 6942 11994 6966 11996
rect 7022 11994 7046 11996
rect 7102 11994 7126 11996
rect 7182 11994 7188 11996
rect 6942 11942 6944 11994
rect 7124 11942 7126 11994
rect 6880 11940 6886 11942
rect 6942 11940 6966 11942
rect 7022 11940 7046 11942
rect 7102 11940 7126 11942
rect 7182 11940 7188 11942
rect 6880 11920 7188 11940
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 7472 11756 7524 11762
rect 7576 11744 7604 12378
rect 7668 12238 7696 14894
rect 7760 14532 7788 15456
rect 7852 15026 7880 15574
rect 7944 15434 7972 15846
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 8036 15162 8064 16050
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8312 15502 8340 15574
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8220 15026 8248 15302
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8220 14822 8248 14962
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8312 14550 8340 15438
rect 8496 15026 8524 15506
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 8680 15026 8708 15370
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8482 14784 8538 14793
rect 8482 14719 8538 14728
rect 8300 14544 8352 14550
rect 7760 14504 7972 14532
rect 7748 14408 7800 14414
rect 7746 14376 7748 14385
rect 7800 14376 7802 14385
rect 7746 14311 7802 14320
rect 7760 13938 7788 14311
rect 7944 14278 7972 14504
rect 8300 14486 8352 14492
rect 8312 14346 8340 14486
rect 8496 14346 8524 14719
rect 8942 14648 8998 14657
rect 8942 14583 8998 14592
rect 8956 14550 8984 14583
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 9036 14340 9088 14346
rect 9036 14282 9088 14288
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7944 13734 7972 13874
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7944 13326 7972 13670
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7656 12232 7708 12238
rect 7708 12192 7788 12220
rect 7656 12174 7708 12180
rect 7524 11716 7696 11744
rect 7472 11698 7524 11704
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5552 10674 5580 10950
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 3915 9276 4223 9296
rect 3915 9274 3921 9276
rect 3977 9274 4001 9276
rect 4057 9274 4081 9276
rect 4137 9274 4161 9276
rect 4217 9274 4223 9276
rect 3977 9222 3979 9274
rect 4159 9222 4161 9274
rect 3915 9220 3921 9222
rect 3977 9220 4001 9222
rect 4057 9220 4081 9222
rect 4137 9220 4161 9222
rect 4217 9220 4223 9222
rect 3915 9200 4223 9220
rect 4264 9178 4292 9522
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4448 8945 4476 9318
rect 4434 8936 4490 8945
rect 4434 8871 4490 8880
rect 4448 8838 4476 8871
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 3436 8566 3464 8774
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 2792 7886 2820 8366
rect 3160 7954 3188 8366
rect 3915 8188 4223 8208
rect 3915 8186 3921 8188
rect 3977 8186 4001 8188
rect 4057 8186 4081 8188
rect 4137 8186 4161 8188
rect 4217 8186 4223 8188
rect 3977 8134 3979 8186
rect 4159 8134 4161 8186
rect 3915 8132 3921 8134
rect 3977 8132 4001 8134
rect 4057 8132 4081 8134
rect 4137 8132 4161 8134
rect 4217 8132 4223 8134
rect 3915 8112 4223 8132
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2502 6896 2558 6905
rect 2700 6866 2728 7278
rect 3068 7206 3096 7686
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 2502 6831 2558 6840
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1964 5234 1992 6054
rect 2608 5710 2636 6598
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2792 5370 2820 6734
rect 3068 6662 3096 7142
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 6458 3096 6598
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2976 5914 3004 6326
rect 3160 6254 3188 7890
rect 3915 7100 4223 7120
rect 3915 7098 3921 7100
rect 3977 7098 4001 7100
rect 4057 7098 4081 7100
rect 4137 7098 4161 7100
rect 4217 7098 4223 7100
rect 3977 7046 3979 7098
rect 4159 7046 4161 7098
rect 3915 7044 3921 7046
rect 3977 7044 4001 7046
rect 4057 7044 4081 7046
rect 4137 7044 4161 7046
rect 4217 7044 4223 7046
rect 3915 7024 4223 7044
rect 4356 6866 4384 7890
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 3528 6254 3556 6802
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4172 6458 4200 6734
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3516 6248 3568 6254
rect 3804 6202 3832 6258
rect 4356 6254 4384 6802
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 3516 6190 3568 6196
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2976 5302 3004 5850
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1584 5092 1636 5098
rect 1584 5034 1636 5040
rect 1596 4690 1624 5034
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1596 3670 1624 4626
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1688 4282 1716 4490
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1780 4078 1808 5170
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 2044 4004 2096 4010
rect 2044 3946 2096 3952
rect 1584 3664 1636 3670
rect 1584 3606 1636 3612
rect 2056 3602 2084 3946
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2056 3126 2084 3538
rect 2044 3120 2096 3126
rect 2044 3062 2096 3068
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 1308 2508 1360 2514
rect 1308 2450 1360 2456
rect 1320 800 1348 2450
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 1964 2106 1992 2382
rect 2056 2310 2084 2926
rect 2240 2825 2268 2926
rect 2226 2816 2282 2825
rect 2226 2751 2282 2760
rect 2332 2514 2360 4422
rect 2424 4146 2452 4966
rect 3068 4826 3096 5306
rect 3160 5166 3188 6190
rect 3712 6174 3832 6202
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 3712 5914 3740 6174
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3712 4826 3740 5170
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3068 4282 3096 4762
rect 3804 4622 3832 6054
rect 3915 6012 4223 6032
rect 3915 6010 3921 6012
rect 3977 6010 4001 6012
rect 4057 6010 4081 6012
rect 4137 6010 4161 6012
rect 4217 6010 4223 6012
rect 3977 5958 3979 6010
rect 4159 5958 4161 6010
rect 3915 5956 3921 5958
rect 3977 5956 4001 5958
rect 4057 5956 4081 5958
rect 4137 5956 4161 5958
rect 4217 5956 4223 5958
rect 3915 5936 4223 5956
rect 4356 5778 4384 6190
rect 4540 5914 4568 6598
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4356 5370 4384 5510
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 3915 4924 4223 4944
rect 3915 4922 3921 4924
rect 3977 4922 4001 4924
rect 4057 4922 4081 4924
rect 4137 4922 4161 4924
rect 4217 4922 4223 4924
rect 3977 4870 3979 4922
rect 4159 4870 4161 4922
rect 3915 4868 3921 4870
rect 3977 4868 4001 4870
rect 4057 4868 4081 4870
rect 4137 4868 4161 4870
rect 4217 4868 4223 4870
rect 3915 4848 4223 4868
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 2516 3754 2544 4014
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2424 3738 2544 3754
rect 2412 3732 2544 3738
rect 2464 3726 2544 3732
rect 2412 3674 2464 3680
rect 2516 3058 2544 3726
rect 2700 3058 2728 3878
rect 2792 3534 2820 4014
rect 3436 3670 3464 4014
rect 3620 3738 3648 4014
rect 3915 3836 4223 3856
rect 3915 3834 3921 3836
rect 3977 3834 4001 3836
rect 4057 3834 4081 3836
rect 4137 3834 4161 3836
rect 4217 3834 4223 3836
rect 3977 3782 3979 3834
rect 4159 3782 4161 3834
rect 3915 3780 3921 3782
rect 3977 3780 4001 3782
rect 4057 3780 4081 3782
rect 4137 3780 4161 3782
rect 4217 3780 4223 3782
rect 3915 3760 4223 3780
rect 4264 3738 4292 4082
rect 4528 4072 4580 4078
rect 4632 4060 4660 9930
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9518 4752 9862
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4724 9194 4752 9454
rect 4724 9166 4844 9194
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4724 7954 4752 8978
rect 4816 8566 4844 9166
rect 5276 8906 5304 10406
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 4804 8560 4856 8566
rect 5184 8537 5212 8570
rect 4804 8502 4856 8508
rect 5170 8528 5226 8537
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4816 7342 4844 8502
rect 5170 8463 5226 8472
rect 5184 7886 5212 8463
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4816 6934 4844 7278
rect 4908 7002 4936 7346
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 6458 5212 6598
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5184 6361 5212 6394
rect 5170 6352 5226 6361
rect 5276 6338 5304 8842
rect 5368 7562 5396 10202
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5552 9654 5580 9998
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5736 9586 5764 9862
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5460 8634 5488 8910
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5644 8090 5672 8434
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5920 7954 5948 11290
rect 6012 11150 6040 11290
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 6012 9586 6040 10678
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6564 9110 6592 11698
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6656 10538 6684 11562
rect 6748 11354 6776 11698
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 10690 6776 11086
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 6880 10908 7188 10928
rect 6880 10906 6886 10908
rect 6942 10906 6966 10908
rect 7022 10906 7046 10908
rect 7102 10906 7126 10908
rect 7182 10906 7188 10908
rect 6942 10854 6944 10906
rect 7124 10854 7126 10906
rect 6880 10852 6886 10854
rect 6942 10852 6966 10854
rect 7022 10852 7046 10854
rect 7102 10852 7126 10854
rect 7182 10852 7188 10854
rect 6880 10832 7188 10852
rect 6748 10662 6960 10690
rect 7300 10674 7328 10950
rect 7484 10742 7512 11222
rect 7576 11218 7604 11494
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7668 11150 7696 11716
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 6932 10554 6960 10662
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7472 10600 7524 10606
rect 6644 10532 6696 10538
rect 6932 10526 7328 10554
rect 7472 10542 7524 10548
rect 6644 10474 6696 10480
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6104 8090 6132 8910
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6472 8498 6500 8774
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 6564 7886 6592 9046
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5368 7534 5488 7562
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5368 6730 5396 7346
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5276 6310 5396 6338
rect 5170 6287 5226 6296
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5276 5778 5304 6122
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5000 5098 5028 5646
rect 5368 5234 5396 6310
rect 5460 5370 5488 7534
rect 5552 6390 5580 7754
rect 6656 7478 6684 10474
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6748 9722 6776 9930
rect 6880 9820 7188 9840
rect 6880 9818 6886 9820
rect 6942 9818 6966 9820
rect 7022 9818 7046 9820
rect 7102 9818 7126 9820
rect 7182 9818 7188 9820
rect 6942 9766 6944 9818
rect 7124 9766 7126 9818
rect 6880 9764 6886 9766
rect 6942 9764 6966 9766
rect 7022 9764 7046 9766
rect 7102 9764 7126 9766
rect 7182 9764 7188 9766
rect 6880 9744 7188 9764
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 7300 9586 7328 10526
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7484 9518 7512 10542
rect 7576 10538 7604 11018
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7668 10062 7696 11086
rect 7760 10742 7788 12192
rect 7852 11830 7880 13262
rect 8128 13258 8156 14214
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8864 13870 8892 13942
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8220 13530 8248 13670
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 8864 12306 8892 13806
rect 9048 13326 9076 14282
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9048 12374 9076 12718
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 8864 11286 8892 12242
rect 9048 12170 9076 12310
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9140 11762 9168 16594
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 16250 9444 16458
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9218 16008 9274 16017
rect 9218 15943 9220 15952
rect 9272 15943 9274 15952
rect 9220 15914 9272 15920
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9324 14618 9352 14894
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9324 14278 9352 14554
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9416 14006 9444 14758
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9232 12782 9260 13126
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9232 12306 9260 12718
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9324 12102 9352 12786
rect 9508 12434 9536 17070
rect 9846 16892 10154 16912
rect 9846 16890 9852 16892
rect 9908 16890 9932 16892
rect 9988 16890 10012 16892
rect 10068 16890 10092 16892
rect 10148 16890 10154 16892
rect 9908 16838 9910 16890
rect 10090 16838 10092 16890
rect 9846 16836 9852 16838
rect 9908 16836 9932 16838
rect 9988 16836 10012 16838
rect 10068 16836 10092 16838
rect 10148 16836 10154 16838
rect 9846 16816 10154 16836
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10244 16250 10272 16526
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10336 16114 10364 16594
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 9846 15804 10154 15824
rect 9846 15802 9852 15804
rect 9908 15802 9932 15804
rect 9988 15802 10012 15804
rect 10068 15802 10092 15804
rect 10148 15802 10154 15804
rect 9908 15750 9910 15802
rect 10090 15750 10092 15802
rect 9846 15748 9852 15750
rect 9908 15748 9932 15750
rect 9988 15748 10012 15750
rect 10068 15748 10092 15750
rect 10148 15748 10154 15750
rect 9846 15728 10154 15748
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9600 15026 9628 15438
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9692 14618 9720 14894
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9600 13734 9628 14350
rect 9784 14346 9812 15438
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 9846 14716 10154 14736
rect 9846 14714 9852 14716
rect 9908 14714 9932 14716
rect 9988 14714 10012 14716
rect 10068 14714 10092 14716
rect 10148 14714 10154 14716
rect 9908 14662 9910 14714
rect 10090 14662 10092 14714
rect 9846 14660 9852 14662
rect 9908 14660 9932 14662
rect 9988 14660 10012 14662
rect 10068 14660 10092 14662
rect 10148 14660 10154 14662
rect 9846 14640 10154 14660
rect 10140 14544 10192 14550
rect 10138 14512 10140 14521
rect 10192 14512 10194 14521
rect 10138 14447 10194 14456
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 13938 9720 14214
rect 10152 13938 10180 14447
rect 10244 14278 10272 14962
rect 10428 14770 10456 17138
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10336 14742 10456 14770
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9846 13628 10154 13648
rect 9846 13626 9852 13628
rect 9908 13626 9932 13628
rect 9988 13626 10012 13628
rect 10068 13626 10092 13628
rect 10148 13626 10154 13628
rect 9908 13574 9910 13626
rect 10090 13574 10092 13626
rect 9846 13572 9852 13574
rect 9908 13572 9932 13574
rect 9988 13572 10012 13574
rect 10068 13572 10092 13574
rect 10148 13572 10154 13574
rect 9846 13552 10154 13572
rect 9846 12540 10154 12560
rect 9846 12538 9852 12540
rect 9908 12538 9932 12540
rect 9988 12538 10012 12540
rect 10068 12538 10092 12540
rect 10148 12538 10154 12540
rect 9908 12486 9910 12538
rect 10090 12486 10092 12538
rect 9846 12484 9852 12486
rect 9908 12484 9932 12486
rect 9988 12484 10012 12486
rect 10068 12484 10092 12486
rect 10148 12484 10154 12486
rect 9846 12464 10154 12484
rect 9416 12406 9536 12434
rect 10336 12434 10364 14742
rect 10520 13802 10548 14758
rect 10508 13796 10560 13802
rect 10508 13738 10560 13744
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10428 12986 10456 13194
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10336 12406 10548 12434
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9324 11354 9352 11698
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7760 10198 7788 10678
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 9722 7604 9862
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 6880 8732 7188 8752
rect 6880 8730 6886 8732
rect 6942 8730 6966 8732
rect 7022 8730 7046 8732
rect 7102 8730 7126 8732
rect 7182 8730 7188 8732
rect 6942 8678 6944 8730
rect 7124 8678 7126 8730
rect 6880 8676 6886 8678
rect 6942 8676 6966 8678
rect 7022 8676 7046 8678
rect 7102 8676 7126 8678
rect 7182 8676 7188 8678
rect 6880 8656 7188 8676
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 6880 7644 7188 7664
rect 6880 7642 6886 7644
rect 6942 7642 6966 7644
rect 7022 7642 7046 7644
rect 7102 7642 7126 7644
rect 7182 7642 7188 7644
rect 6942 7590 6944 7642
rect 7124 7590 7126 7642
rect 6880 7588 6886 7590
rect 6942 7588 6966 7590
rect 7022 7588 7046 7590
rect 7102 7588 7126 7590
rect 7182 7588 7188 7590
rect 6880 7568 7188 7588
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5920 6322 5948 7210
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 6798 6316 7142
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 5710 5580 6054
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4908 4146 4936 4422
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4580 4032 4660 4060
rect 4528 4014 4580 4020
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3148 3460 3200 3466
rect 3148 3402 3200 3408
rect 3160 3194 3188 3402
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 1952 2100 2004 2106
rect 1952 2042 2004 2048
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 2792 785 2820 2382
rect 3252 800 3280 3470
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 3915 2748 4223 2768
rect 3915 2746 3921 2748
rect 3977 2746 4001 2748
rect 4057 2746 4081 2748
rect 4137 2746 4161 2748
rect 4217 2746 4223 2748
rect 3977 2694 3979 2746
rect 4159 2694 4161 2746
rect 3915 2692 3921 2694
rect 3977 2692 4001 2694
rect 4057 2692 4081 2694
rect 4137 2692 4161 2694
rect 4217 2692 4223 2694
rect 3915 2672 4223 2692
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3436 1465 3464 2586
rect 4264 2582 4292 2994
rect 4252 2576 4304 2582
rect 4252 2518 4304 2524
rect 4356 2446 4384 3878
rect 4632 3602 4660 4032
rect 5092 3738 5120 4558
rect 5368 4146 5396 5170
rect 5460 5166 5488 5306
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5460 4690 5488 5102
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 6288 4622 6316 4966
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 5356 4140 5408 4146
rect 5408 4100 5488 4128
rect 5356 4082 5408 4088
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5460 3602 5488 4100
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 4632 3126 4660 3538
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 5552 2922 5580 3606
rect 5644 3398 5672 3946
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5736 3058 5764 3606
rect 6564 3602 6592 4626
rect 6656 3670 6684 7210
rect 7300 6866 7328 8502
rect 7484 8498 7512 9454
rect 7576 8974 7604 9658
rect 7668 9586 7696 9998
rect 7760 9654 7788 10134
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7852 9178 7880 10610
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 9586 7972 10406
rect 8128 10062 8156 11086
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8128 9722 8156 9998
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 9324 9586 9352 9930
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8128 8634 8156 8910
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7392 7886 7420 8230
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7410 7420 7822
rect 7484 7546 7512 8434
rect 7760 8022 7788 8570
rect 8220 8498 8248 8910
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8404 8566 8432 8774
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7838 7984 7894 7993
rect 7760 7818 7788 7958
rect 8496 7954 8524 8774
rect 7838 7919 7840 7928
rect 7892 7919 7894 7928
rect 8484 7948 8536 7954
rect 7840 7890 7892 7896
rect 8484 7890 8536 7896
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 6880 6556 7188 6576
rect 6880 6554 6886 6556
rect 6942 6554 6966 6556
rect 7022 6554 7046 6556
rect 7102 6554 7126 6556
rect 7182 6554 7188 6556
rect 6942 6502 6944 6554
rect 7124 6502 7126 6554
rect 6880 6500 6886 6502
rect 6942 6500 6966 6502
rect 7022 6500 7046 6502
rect 7102 6500 7126 6502
rect 7182 6500 7188 6502
rect 6880 6480 7188 6500
rect 7300 6458 7328 6802
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6932 5778 6960 6326
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6880 5468 7188 5488
rect 6880 5466 6886 5468
rect 6942 5466 6966 5468
rect 7022 5466 7046 5468
rect 7102 5466 7126 5468
rect 7182 5466 7188 5468
rect 6942 5414 6944 5466
rect 7124 5414 7126 5466
rect 6880 5412 6886 5414
rect 6942 5412 6966 5414
rect 7022 5412 7046 5414
rect 7102 5412 7126 5414
rect 7182 5412 7188 5414
rect 6880 5392 7188 5412
rect 7300 5166 7328 6394
rect 7392 6254 7420 7210
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 8114 6760 8170 6769
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7576 6458 7604 6666
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7668 6118 7696 6734
rect 8114 6695 8170 6704
rect 8128 6662 8156 6695
rect 8116 6656 8168 6662
rect 8036 6616 8116 6644
rect 8036 6322 8064 6616
rect 8116 6598 8168 6604
rect 8220 6322 8248 6870
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6458 8340 6598
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8588 6390 8616 7278
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 6104 2446 6132 3334
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6564 2582 6592 2994
rect 6748 2922 6776 5102
rect 7196 4616 7248 4622
rect 7300 4604 7328 5102
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4622 7420 4966
rect 7484 4826 7512 5578
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7248 4576 7328 4604
rect 7196 4558 7248 4564
rect 6880 4380 7188 4400
rect 6880 4378 6886 4380
rect 6942 4378 6966 4380
rect 7022 4378 7046 4380
rect 7102 4378 7126 4380
rect 7182 4378 7188 4380
rect 6942 4326 6944 4378
rect 7124 4326 7126 4378
rect 6880 4324 6886 4326
rect 6942 4324 6966 4326
rect 7022 4324 7046 4326
rect 7102 4324 7126 4326
rect 7182 4324 7188 4326
rect 6880 4304 7188 4324
rect 7300 4214 7328 4576
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7196 4072 7248 4078
rect 7248 4032 7328 4060
rect 7196 4014 7248 4020
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6932 3534 6960 3878
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6880 3292 7188 3312
rect 6880 3290 6886 3292
rect 6942 3290 6966 3292
rect 7022 3290 7046 3292
rect 7102 3290 7126 3292
rect 7182 3290 7188 3292
rect 6942 3238 6944 3290
rect 7124 3238 7126 3290
rect 6880 3236 6886 3238
rect 6942 3236 6966 3238
rect 7022 3236 7046 3238
rect 7102 3236 7126 3238
rect 7182 3236 7188 3238
rect 6880 3216 7188 3236
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 6748 2446 6776 2858
rect 7116 2514 7144 3062
rect 7300 2836 7328 4032
rect 7576 3738 7604 5170
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7380 2848 7432 2854
rect 7300 2808 7380 2836
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7300 2446 7328 2808
rect 7380 2790 7432 2796
rect 7668 2774 7696 6054
rect 8404 5710 8432 6326
rect 8772 6322 8800 8910
rect 9140 8498 9168 9114
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9140 7954 9168 8434
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 7478 8984 7686
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 8956 7002 8984 7414
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 5370 8340 5510
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7760 4826 7788 5034
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8496 4282 8524 4422
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7760 3058 7788 4082
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7852 2922 7880 3062
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7484 2746 7696 2774
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4344 2440 4396 2446
rect 5540 2440 5592 2446
rect 4344 2382 4396 2388
rect 5460 2388 5540 2394
rect 5460 2382 5592 2388
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 3422 1456 3478 1465
rect 3422 1391 3478 1400
rect 3896 800 3924 2382
rect 5460 2366 5580 2382
rect 6460 2372 6512 2378
rect 5184 870 5304 898
rect 5184 800 5212 870
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 5276 762 5304 870
rect 5460 762 5488 2366
rect 6460 2314 6512 2320
rect 6472 800 6500 2314
rect 6880 2204 7188 2224
rect 6880 2202 6886 2204
rect 6942 2202 6966 2204
rect 7022 2202 7046 2204
rect 7102 2202 7126 2204
rect 7182 2202 7188 2204
rect 6942 2150 6944 2202
rect 7124 2150 7126 2202
rect 6880 2148 6886 2150
rect 6942 2148 6966 2150
rect 7022 2148 7046 2150
rect 7102 2148 7126 2150
rect 7182 2148 7188 2150
rect 6880 2128 7188 2148
rect 7484 2106 7512 2746
rect 8864 2582 8892 5782
rect 9140 4690 9168 7890
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8956 3738 8984 4082
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9140 3924 9168 4626
rect 9220 3936 9272 3942
rect 9140 3896 9220 3924
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9048 3126 9076 3878
rect 9140 3602 9168 3896
rect 9220 3878 9272 3884
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9232 3194 9260 3470
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 9048 2446 9076 3062
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9140 2582 9168 2994
rect 9324 2650 9352 9522
rect 9416 6934 9444 12406
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9600 11150 9628 11698
rect 10336 11558 10364 12106
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 9846 11452 10154 11472
rect 9846 11450 9852 11452
rect 9908 11450 9932 11452
rect 9988 11450 10012 11452
rect 10068 11450 10092 11452
rect 10148 11450 10154 11452
rect 9908 11398 9910 11450
rect 10090 11398 10092 11450
rect 9846 11396 9852 11398
rect 9908 11396 9932 11398
rect 9988 11396 10012 11398
rect 10068 11396 10092 11398
rect 10148 11396 10154 11398
rect 9846 11376 10154 11396
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9784 10810 9812 11086
rect 10336 11082 10364 11494
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 8974 9628 10406
rect 9692 9926 9720 10610
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9692 8974 9720 9658
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9508 8362 9536 8842
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9508 7342 9536 8298
rect 9692 7546 9720 8366
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9404 6928 9456 6934
rect 9404 6870 9456 6876
rect 9508 4758 9536 7278
rect 9784 7274 9812 10542
rect 9846 10364 10154 10384
rect 9846 10362 9852 10364
rect 9908 10362 9932 10364
rect 9988 10362 10012 10364
rect 10068 10362 10092 10364
rect 10148 10362 10154 10364
rect 9908 10310 9910 10362
rect 10090 10310 10092 10362
rect 9846 10308 9852 10310
rect 9908 10308 9932 10310
rect 9988 10308 10012 10310
rect 10068 10308 10092 10310
rect 10148 10308 10154 10310
rect 9846 10288 10154 10308
rect 9846 9276 10154 9296
rect 9846 9274 9852 9276
rect 9908 9274 9932 9276
rect 9988 9274 10012 9276
rect 10068 9274 10092 9276
rect 10148 9274 10154 9276
rect 9908 9222 9910 9274
rect 10090 9222 10092 9274
rect 9846 9220 9852 9222
rect 9908 9220 9932 9222
rect 9988 9220 10012 9222
rect 10068 9220 10092 9222
rect 10148 9220 10154 9222
rect 9846 9200 10154 9220
rect 10244 9178 10272 10610
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 9846 8188 10154 8208
rect 9846 8186 9852 8188
rect 9908 8186 9932 8188
rect 9988 8186 10012 8188
rect 10068 8186 10092 8188
rect 10148 8186 10154 8188
rect 9908 8134 9910 8186
rect 10090 8134 10092 8186
rect 9846 8132 9852 8134
rect 9908 8132 9932 8134
rect 9988 8132 10012 8134
rect 10068 8132 10092 8134
rect 10148 8132 10154 8134
rect 9846 8112 10154 8132
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9846 7100 10154 7120
rect 9846 7098 9852 7100
rect 9908 7098 9932 7100
rect 9988 7098 10012 7100
rect 10068 7098 10092 7100
rect 10148 7098 10154 7100
rect 9908 7046 9910 7098
rect 10090 7046 10092 7098
rect 9846 7044 9852 7046
rect 9908 7044 9932 7046
rect 9988 7044 10012 7046
rect 10068 7044 10092 7046
rect 10148 7044 10154 7046
rect 9846 7024 10154 7044
rect 10244 6882 10272 8502
rect 10336 7478 10364 11018
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10428 10062 10456 10406
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10428 9178 10456 9318
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10520 8566 10548 12406
rect 10612 11150 10640 16934
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10782 16144 10838 16153
rect 10782 16079 10838 16088
rect 10876 16108 10928 16114
rect 10796 15910 10824 16079
rect 10876 16050 10928 16056
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10888 15706 10916 16050
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 14346 10732 15302
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10888 14822 10916 14962
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10796 14006 10824 14554
rect 10888 14482 10916 14758
rect 10980 14618 11008 16594
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10704 12889 10732 13738
rect 11072 13462 11100 17002
rect 11624 16726 11652 17138
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11900 16590 11928 16934
rect 12268 16658 12572 16674
rect 12256 16652 12572 16658
rect 12308 16646 12572 16652
rect 12256 16594 12308 16600
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11256 15638 11284 16390
rect 11716 16046 11744 16526
rect 12164 16448 12216 16454
rect 11992 16396 12164 16402
rect 11992 16390 12216 16396
rect 11992 16374 12204 16390
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11992 15910 12020 16374
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11244 15632 11296 15638
rect 11244 15574 11296 15580
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11164 14346 11192 15438
rect 11256 14414 11284 15574
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11348 14890 11376 15506
rect 11992 15366 12020 15846
rect 12084 15502 12112 15982
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11336 14884 11388 14890
rect 11336 14826 11388 14832
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11348 14346 11376 14826
rect 11716 14822 11744 15302
rect 11992 15162 12020 15302
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11992 14618 12020 15098
rect 12084 15026 12112 15438
rect 12360 15094 12388 15846
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 12452 14958 12480 16526
rect 12544 16250 12572 16646
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12636 16153 12664 17070
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 14844 16590 14872 16934
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 12811 16348 13119 16368
rect 12811 16346 12817 16348
rect 12873 16346 12897 16348
rect 12953 16346 12977 16348
rect 13033 16346 13057 16348
rect 13113 16346 13119 16348
rect 12873 16294 12875 16346
rect 13055 16294 13057 16346
rect 12811 16292 12817 16294
rect 12873 16292 12897 16294
rect 12953 16292 12977 16294
rect 13033 16292 13057 16294
rect 13113 16292 13119 16294
rect 12811 16272 13119 16292
rect 13464 16250 13492 16390
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 12716 16176 12768 16182
rect 12622 16144 12678 16153
rect 12716 16118 12768 16124
rect 12990 16144 13046 16153
rect 12622 16079 12678 16088
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12636 15706 12664 15914
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12544 15094 12572 15438
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 12636 14550 12664 15302
rect 12728 15162 12756 16118
rect 13740 16114 13768 16390
rect 15028 16250 15056 17138
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 12990 16079 13046 16088
rect 13268 16108 13320 16114
rect 13004 15910 13032 16079
rect 13268 16050 13320 16056
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 13004 15638 13032 15846
rect 12992 15632 13044 15638
rect 12992 15574 13044 15580
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 12811 15260 13119 15280
rect 12811 15258 12817 15260
rect 12873 15258 12897 15260
rect 12953 15258 12977 15260
rect 13033 15258 13057 15260
rect 13113 15258 13119 15260
rect 12873 15206 12875 15258
rect 13055 15206 13057 15258
rect 12811 15204 12817 15206
rect 12873 15204 12897 15206
rect 12953 15204 12977 15206
rect 13033 15204 13057 15206
rect 13113 15204 13119 15206
rect 12811 15184 13119 15204
rect 13188 15162 13216 15370
rect 13280 15366 13308 16050
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13556 15502 13584 15846
rect 14016 15502 14044 15846
rect 15212 15706 15240 16118
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15304 15570 15332 16186
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13464 15094 13492 15302
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 11164 14074 11192 14282
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 10690 12880 10746 12889
rect 11256 12850 11284 13398
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 10690 12815 10692 12824
rect 10744 12815 10746 12824
rect 10876 12844 10928 12850
rect 10692 12786 10744 12792
rect 10876 12786 10928 12792
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 10704 12755 10732 12786
rect 10888 12442 10916 12786
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10796 11150 10824 11494
rect 10980 11354 11008 11698
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10968 11008 11020 11014
rect 11072 10996 11100 12786
rect 11440 11694 11468 13262
rect 11808 13258 11836 13670
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11348 11354 11376 11630
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11020 10968 11100 10996
rect 10968 10950 11020 10956
rect 10692 10736 10744 10742
rect 10612 10684 10692 10690
rect 10612 10678 10744 10684
rect 10612 10662 10732 10678
rect 10612 9382 10640 10662
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 9042 10640 9318
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 8566 10640 8774
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 7886 10456 8230
rect 10704 7886 10732 9862
rect 10796 9722 10824 9930
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 9722 10916 9862
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10874 9072 10930 9081
rect 10874 9007 10930 9016
rect 10888 8634 10916 9007
rect 10980 8974 11008 10950
rect 11164 10810 11192 11018
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11348 10062 11376 10678
rect 11440 10130 11468 11630
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11532 10062 11560 10610
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11348 9382 11376 9998
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11532 9178 11560 9998
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10876 8628 10928 8634
rect 10796 8588 10876 8616
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 9784 6854 10272 6882
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9692 6254 9720 6734
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9692 5846 9720 6190
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9692 5642 9720 5782
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9784 5386 9812 6854
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10060 6458 10088 6734
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10152 6186 10180 6598
rect 10244 6458 10272 6734
rect 10520 6730 10548 7754
rect 10690 7712 10746 7721
rect 10690 7647 10746 7656
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 9846 6012 10154 6032
rect 9846 6010 9852 6012
rect 9908 6010 9932 6012
rect 9988 6010 10012 6012
rect 10068 6010 10092 6012
rect 10148 6010 10154 6012
rect 9908 5958 9910 6010
rect 10090 5958 10092 6010
rect 9846 5956 9852 5958
rect 9908 5956 9932 5958
rect 9988 5956 10012 5958
rect 10068 5956 10092 5958
rect 10148 5956 10154 5958
rect 9846 5936 10154 5956
rect 10244 5642 10272 6394
rect 10336 5914 10364 6666
rect 10506 6624 10562 6633
rect 10506 6559 10562 6568
rect 10520 6322 10548 6559
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10520 5778 10548 6054
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9692 5358 9812 5386
rect 9692 5030 9720 5358
rect 9876 5302 9904 5510
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9508 4128 9536 4694
rect 9784 4146 9812 5170
rect 9968 5137 9996 5578
rect 10506 5400 10562 5409
rect 10506 5335 10562 5344
rect 10520 5302 10548 5335
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 9954 5128 10010 5137
rect 9954 5063 10010 5072
rect 9846 4924 10154 4944
rect 9846 4922 9852 4924
rect 9908 4922 9932 4924
rect 9988 4922 10012 4924
rect 10068 4922 10092 4924
rect 10148 4922 10154 4924
rect 9908 4870 9910 4922
rect 10090 4870 10092 4922
rect 9846 4868 9852 4870
rect 9908 4868 9932 4870
rect 9988 4868 10012 4870
rect 10068 4868 10092 4870
rect 10148 4868 10154 4870
rect 9846 4848 10154 4868
rect 9588 4140 9640 4146
rect 9508 4100 9588 4128
rect 9588 4082 9640 4088
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9600 3534 9628 4082
rect 10244 4010 10272 5170
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10428 4146 10456 4966
rect 10520 4554 10548 5238
rect 10612 4622 10640 7142
rect 10704 6474 10732 7647
rect 10796 6644 10824 8588
rect 10876 8570 10928 8576
rect 10876 7880 10928 7886
rect 10980 7857 11008 8910
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 11072 7954 11100 8842
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 10876 7822 10928 7828
rect 10966 7848 11022 7857
rect 10888 7274 10916 7822
rect 10966 7783 11022 7792
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 7410 11008 7686
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10876 6656 10928 6662
rect 10796 6616 10876 6644
rect 10980 6644 11008 7210
rect 11072 6798 11100 7890
rect 11164 7546 11192 9114
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10980 6616 11100 6644
rect 10876 6598 10928 6604
rect 10704 6446 10824 6474
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10704 5914 10732 6122
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10692 5704 10744 5710
rect 10690 5672 10692 5681
rect 10744 5672 10746 5681
rect 10690 5607 10746 5616
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10796 4010 10824 6446
rect 10888 6225 10916 6598
rect 10971 6316 11023 6322
rect 11072 6304 11100 6616
rect 11164 6458 11192 7210
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11152 6316 11204 6322
rect 11072 6276 11152 6304
rect 10971 6258 11023 6264
rect 11152 6258 11204 6264
rect 10874 6216 10930 6225
rect 10874 6151 10930 6160
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10888 5137 10916 5850
rect 10980 5710 11008 6258
rect 10968 5704 11020 5710
rect 11152 5704 11204 5710
rect 10968 5646 11020 5652
rect 11150 5672 11152 5681
rect 11204 5672 11206 5681
rect 11060 5636 11112 5642
rect 11150 5607 11206 5616
rect 11060 5578 11112 5584
rect 11072 5370 11100 5578
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11164 5250 11192 5607
rect 10980 5222 11192 5250
rect 10874 5128 10930 5137
rect 10874 5063 10930 5072
rect 10980 4282 11008 5222
rect 11164 5166 11192 5222
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10980 4146 11008 4218
rect 11256 4146 11284 8978
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11440 7002 11468 7686
rect 11532 7410 11560 7754
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11348 6633 11376 6734
rect 11334 6624 11390 6633
rect 11334 6559 11390 6568
rect 11334 5264 11390 5273
rect 11334 5199 11336 5208
rect 11388 5199 11390 5208
rect 11336 5170 11388 5176
rect 11348 4690 11376 5170
rect 11440 4690 11468 6938
rect 11624 6390 11652 12106
rect 11900 10674 11928 13466
rect 12268 12374 12296 13874
rect 12360 12918 12388 13942
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12452 12442 12480 14282
rect 12544 12850 12572 14350
rect 12728 13938 12756 14894
rect 14016 14550 14044 15438
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 15212 15162 15240 15370
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15396 14770 15424 17002
rect 15488 16538 15516 19200
rect 16302 17776 16358 17785
rect 16302 17711 16358 17720
rect 16316 17134 16344 17711
rect 16776 17202 16804 19200
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 15776 16892 16084 16912
rect 15776 16890 15782 16892
rect 15838 16890 15862 16892
rect 15918 16890 15942 16892
rect 15998 16890 16022 16892
rect 16078 16890 16084 16892
rect 15838 16838 15840 16890
rect 16020 16838 16022 16890
rect 15776 16836 15782 16838
rect 15838 16836 15862 16838
rect 15918 16836 15942 16838
rect 15998 16836 16022 16838
rect 16078 16836 16084 16838
rect 15776 16816 16084 16836
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 15488 16510 15608 16538
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 16182 15516 16390
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 15488 15502 15516 16118
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15488 15026 15516 15438
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15396 14742 15516 14770
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 12811 14172 13119 14192
rect 12811 14170 12817 14172
rect 12873 14170 12897 14172
rect 12953 14170 12977 14172
rect 13033 14170 13057 14172
rect 13113 14170 13119 14172
rect 12873 14118 12875 14170
rect 13055 14118 13057 14170
rect 12811 14116 12817 14118
rect 12873 14116 12897 14118
rect 12953 14116 12977 14118
rect 13033 14116 13057 14118
rect 13113 14116 13119 14118
rect 12811 14096 13119 14116
rect 13280 14074 13308 14350
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12256 12368 12308 12374
rect 12256 12310 12308 12316
rect 12544 12306 12572 12786
rect 12636 12714 12664 13806
rect 12728 13462 12756 13874
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 12811 13084 13119 13104
rect 12811 13082 12817 13084
rect 12873 13082 12897 13084
rect 12953 13082 12977 13084
rect 13033 13082 13057 13084
rect 13113 13082 13119 13084
rect 12873 13030 12875 13082
rect 13055 13030 13057 13082
rect 12811 13028 12817 13030
rect 12873 13028 12897 13030
rect 12953 13028 12977 13030
rect 13033 13028 13057 13030
rect 13113 13028 13119 13030
rect 12811 13008 13119 13028
rect 13188 12986 13216 13126
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 13280 12238 13308 14010
rect 13372 14006 13400 14214
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 14108 13734 14136 14350
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 14476 14074 14504 14214
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 12084 11082 12112 12174
rect 12636 11762 12664 12174
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11992 10062 12020 10542
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11716 8906 11744 9998
rect 11886 9480 11942 9489
rect 11886 9415 11942 9424
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11704 8628 11756 8634
rect 11808 8616 11836 9114
rect 11900 8974 11928 9415
rect 11992 9110 12020 9998
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11888 8968 11940 8974
rect 12084 8922 12112 11018
rect 12176 9110 12204 11154
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12268 10674 12296 10950
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12636 10606 12664 11698
rect 12728 11558 12756 12038
rect 12811 11996 13119 12016
rect 12811 11994 12817 11996
rect 12873 11994 12897 11996
rect 12953 11994 12977 11996
rect 13033 11994 13057 11996
rect 13113 11994 13119 11996
rect 12873 11942 12875 11994
rect 13055 11942 13057 11994
rect 12811 11940 12817 11942
rect 12873 11940 12897 11942
rect 12953 11940 12977 11942
rect 13033 11940 13057 11942
rect 13113 11940 13119 11942
rect 12811 11920 13119 11940
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12728 11082 12756 11494
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12268 8974 12296 10406
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12360 9178 12388 9930
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12636 9654 12664 9862
rect 12532 9648 12584 9654
rect 12530 9616 12532 9625
rect 12624 9648 12676 9654
rect 12584 9616 12586 9625
rect 12624 9590 12676 9596
rect 12530 9551 12586 9560
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 11888 8910 11940 8916
rect 11756 8588 11836 8616
rect 11992 8894 12112 8922
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 11704 8570 11756 8576
rect 11992 8242 12020 8894
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12084 8401 12112 8434
rect 12070 8392 12126 8401
rect 12070 8327 12126 8336
rect 12268 8294 12296 8434
rect 12544 8362 12572 8978
rect 12622 8936 12678 8945
rect 12728 8906 12756 11018
rect 12811 10908 13119 10928
rect 12811 10906 12817 10908
rect 12873 10906 12897 10908
rect 12953 10906 12977 10908
rect 13033 10906 13057 10908
rect 13113 10906 13119 10908
rect 12873 10854 12875 10906
rect 13055 10854 13057 10906
rect 12811 10852 12817 10854
rect 12873 10852 12897 10854
rect 12953 10852 12977 10854
rect 13033 10852 13057 10854
rect 13113 10852 13119 10854
rect 12811 10832 13119 10852
rect 13188 10810 13216 12038
rect 13464 11082 13492 13194
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12714 13768 13126
rect 14108 12918 14136 13670
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 14384 12782 14412 13194
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13740 12238 13768 12650
rect 14660 12434 14688 13874
rect 15212 13394 15240 14010
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15028 12918 15056 13126
rect 15304 12986 15332 13874
rect 15396 13462 15424 14214
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15016 12912 15068 12918
rect 14922 12880 14978 12889
rect 15016 12854 15068 12860
rect 14922 12815 14924 12824
rect 14976 12815 14978 12824
rect 14924 12786 14976 12792
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14752 12442 14780 12650
rect 14568 12406 14688 12434
rect 14740 12436 14792 12442
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13280 10538 13308 11018
rect 13464 10742 13492 11018
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13556 10606 13584 11766
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 12811 9820 13119 9840
rect 12811 9818 12817 9820
rect 12873 9818 12897 9820
rect 12953 9818 12977 9820
rect 13033 9818 13057 9820
rect 13113 9818 13119 9820
rect 12873 9766 12875 9818
rect 13055 9766 13057 9818
rect 12811 9764 12817 9766
rect 12873 9764 12897 9766
rect 12953 9764 12977 9766
rect 13033 9764 13057 9766
rect 13113 9764 13119 9766
rect 12811 9744 13119 9764
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12990 9072 13046 9081
rect 13096 9058 13124 9318
rect 13096 9042 13216 9058
rect 12990 9007 13046 9016
rect 13084 9036 13216 9042
rect 13004 8974 13032 9007
rect 13136 9030 13216 9036
rect 13084 8978 13136 8984
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 12622 8871 12678 8880
rect 12716 8900 12768 8906
rect 12636 8786 12664 8871
rect 12716 8842 12768 8848
rect 12636 8758 12756 8786
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12164 8288 12216 8294
rect 11992 8214 12112 8242
rect 12268 8266 12388 8294
rect 12164 8230 12216 8236
rect 11886 7848 11942 7857
rect 11886 7783 11942 7792
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11532 5302 11560 6054
rect 11520 5296 11572 5302
rect 11520 5238 11572 5244
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 9846 3836 10154 3856
rect 9846 3834 9852 3836
rect 9908 3834 9932 3836
rect 9988 3834 10012 3836
rect 10068 3834 10092 3836
rect 10148 3834 10154 3836
rect 9908 3782 9910 3834
rect 10090 3782 10092 3834
rect 9846 3780 9852 3782
rect 9908 3780 9932 3782
rect 9988 3780 10012 3782
rect 10068 3780 10092 3782
rect 10148 3780 10154 3782
rect 9846 3760 10154 3780
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9416 3126 9444 3470
rect 10980 3466 11008 4082
rect 11256 3505 11284 4082
rect 11532 4078 11560 4966
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3534 11468 3878
rect 11428 3528 11480 3534
rect 11242 3496 11298 3505
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 10968 3460 11020 3466
rect 11428 3470 11480 3476
rect 11242 3431 11298 3440
rect 10968 3402 11020 3408
rect 10152 3194 10180 3402
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 9416 2446 9444 3062
rect 9600 2514 9628 3130
rect 9846 2748 10154 2768
rect 9846 2746 9852 2748
rect 9908 2746 9932 2748
rect 9988 2746 10012 2748
rect 10068 2746 10092 2748
rect 10148 2746 10154 2748
rect 9908 2694 9910 2746
rect 10090 2694 10092 2746
rect 9846 2692 9852 2694
rect 9908 2692 9932 2694
rect 9988 2692 10012 2694
rect 10068 2692 10092 2694
rect 10148 2692 10154 2694
rect 9846 2672 10154 2692
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7668 2106 7696 2246
rect 7472 2100 7524 2106
rect 7472 2042 7524 2048
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7760 800 7788 2246
rect 9508 2038 9536 2382
rect 10244 2378 10272 3334
rect 10324 2440 10376 2446
rect 11072 2428 11100 3334
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11164 2650 11192 2994
rect 11624 2854 11652 6326
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11624 2514 11652 2790
rect 11716 2582 11744 6802
rect 11808 6798 11836 7278
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 5386 11836 6598
rect 11900 5914 11928 7783
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11992 6322 12020 6598
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 12084 5778 12112 8214
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12176 5642 12204 8230
rect 12360 8090 12388 8266
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12636 7970 12664 8570
rect 12728 8498 12756 8758
rect 12811 8732 13119 8752
rect 12811 8730 12817 8732
rect 12873 8730 12897 8732
rect 12953 8730 12977 8732
rect 13033 8730 13057 8732
rect 13113 8730 13119 8732
rect 12873 8678 12875 8730
rect 13055 8678 13057 8730
rect 12811 8676 12817 8678
rect 12873 8676 12897 8678
rect 12953 8676 12977 8678
rect 13033 8676 13057 8678
rect 13113 8676 13119 8678
rect 12811 8656 13119 8676
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 8401 13032 8434
rect 12990 8392 13046 8401
rect 12990 8327 13046 8336
rect 12544 7942 12664 7970
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12268 7342 12296 7754
rect 12360 7342 12388 7822
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12254 6896 12310 6905
rect 12348 6860 12400 6866
rect 12310 6840 12348 6848
rect 12254 6831 12348 6840
rect 12268 6820 12348 6831
rect 12268 6662 12296 6820
rect 12348 6802 12400 6808
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12452 6746 12480 6802
rect 12360 6718 12480 6746
rect 12544 6746 12572 7942
rect 12716 7880 12768 7886
rect 12636 7840 12716 7868
rect 12636 7478 12664 7840
rect 12716 7822 12768 7828
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12636 7206 12664 7414
rect 12728 7410 12756 7686
rect 12811 7644 13119 7664
rect 12811 7642 12817 7644
rect 12873 7642 12897 7644
rect 12953 7642 12977 7644
rect 13033 7642 13057 7644
rect 13113 7642 13119 7644
rect 12873 7590 12875 7642
rect 13055 7590 13057 7642
rect 12811 7588 12817 7590
rect 12873 7588 12897 7590
rect 12953 7588 12977 7590
rect 13033 7588 13057 7590
rect 13113 7588 13119 7590
rect 12811 7568 13119 7588
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12728 7274 12756 7346
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12912 7041 12940 7210
rect 12898 7032 12954 7041
rect 12898 6967 12954 6976
rect 12716 6860 12768 6866
rect 12768 6820 12848 6848
rect 12716 6802 12768 6808
rect 12820 6769 12848 6820
rect 12806 6760 12862 6769
rect 12544 6718 12756 6746
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12254 6488 12310 6497
rect 12360 6458 12388 6718
rect 12624 6656 12676 6662
rect 12530 6624 12586 6633
rect 12624 6598 12676 6604
rect 12530 6559 12586 6568
rect 12254 6423 12310 6432
rect 12348 6452 12400 6458
rect 12268 6322 12296 6423
rect 12348 6394 12400 6400
rect 12544 6322 12572 6559
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 11808 5370 12020 5386
rect 11808 5364 12032 5370
rect 11808 5358 11980 5364
rect 11980 5306 12032 5312
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11808 4826 11836 5238
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11992 4622 12020 5306
rect 12176 5234 12204 5578
rect 12360 5409 12388 6258
rect 12636 5914 12664 6598
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12346 5400 12402 5409
rect 12346 5335 12402 5344
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 11900 4146 11928 4422
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 11808 3738 11836 3946
rect 11992 3738 12020 4014
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11152 2440 11204 2446
rect 11072 2400 11152 2428
rect 10324 2382 10376 2388
rect 11152 2382 11204 2388
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 9496 2032 9548 2038
rect 9496 1974 9548 1980
rect 10336 800 10364 2382
rect 11520 2304 11572 2310
rect 11980 2304 12032 2310
rect 11572 2264 11652 2292
rect 11520 2246 11572 2252
rect 11624 800 11652 2264
rect 12084 2292 12112 4422
rect 12176 3670 12204 5170
rect 12268 4282 12296 5170
rect 12452 4826 12480 5646
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12636 4146 12664 5510
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12728 3942 12756 6718
rect 13004 6730 13032 7278
rect 12806 6695 12862 6704
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 12811 6556 13119 6576
rect 12811 6554 12817 6556
rect 12873 6554 12897 6556
rect 12953 6554 12977 6556
rect 13033 6554 13057 6556
rect 13113 6554 13119 6556
rect 12873 6502 12875 6554
rect 13055 6502 13057 6554
rect 12811 6500 12817 6502
rect 12873 6500 12897 6502
rect 12953 6500 12977 6502
rect 13033 6500 13057 6502
rect 13113 6500 13119 6502
rect 12811 6480 13119 6500
rect 13188 6390 13216 9030
rect 13280 7886 13308 10474
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13358 8528 13414 8537
rect 13358 8463 13360 8472
rect 13412 8463 13414 8472
rect 13360 8434 13412 8440
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 13280 5710 13308 7142
rect 13372 6186 13400 8298
rect 13464 7954 13492 8910
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13556 8566 13584 8774
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7002 13492 7890
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13464 6798 13492 6938
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13556 6202 13584 8230
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 13464 6174 13584 6202
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 12811 5468 13119 5488
rect 12811 5466 12817 5468
rect 12873 5466 12897 5468
rect 12953 5466 12977 5468
rect 13033 5466 13057 5468
rect 13113 5466 13119 5468
rect 12873 5414 12875 5466
rect 13055 5414 13057 5466
rect 12811 5412 12817 5414
rect 12873 5412 12897 5414
rect 12953 5412 12977 5414
rect 13033 5412 13057 5414
rect 13113 5412 13119 5414
rect 12811 5392 13119 5412
rect 13372 5370 13400 5510
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 12811 4380 13119 4400
rect 12811 4378 12817 4380
rect 12873 4378 12897 4380
rect 12953 4378 12977 4380
rect 13033 4378 13057 4380
rect 13113 4378 13119 4380
rect 12873 4326 12875 4378
rect 13055 4326 13057 4378
rect 12811 4324 12817 4326
rect 12873 4324 12897 4326
rect 12953 4324 12977 4326
rect 13033 4324 13057 4326
rect 13113 4324 13119 4326
rect 12811 4304 13119 4324
rect 13464 4049 13492 6174
rect 13450 4040 13506 4049
rect 12900 4004 12952 4010
rect 13450 3975 13506 3984
rect 12900 3946 12952 3952
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 12176 3126 12204 3606
rect 12912 3534 12940 3946
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13188 3602 13216 3878
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 12452 3058 12480 3402
rect 12811 3292 13119 3312
rect 12811 3290 12817 3292
rect 12873 3290 12897 3292
rect 12953 3290 12977 3292
rect 13033 3290 13057 3292
rect 13113 3290 13119 3292
rect 12873 3238 12875 3290
rect 13055 3238 13057 3290
rect 12811 3236 12817 3238
rect 12873 3236 12897 3238
rect 12953 3236 12977 3238
rect 13033 3236 13057 3238
rect 13113 3236 13119 3238
rect 12811 3216 13119 3236
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12636 2446 12664 2790
rect 12728 2650 12756 2994
rect 13188 2990 13216 3538
rect 13648 3534 13676 9658
rect 13740 6322 13768 11834
rect 14476 11558 14504 12038
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13832 9450 13860 9930
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13832 7857 13860 8366
rect 13818 7848 13874 7857
rect 13818 7783 13874 7792
rect 13818 7712 13874 7721
rect 13818 7647 13874 7656
rect 13832 6866 13860 7647
rect 13924 7410 13952 9862
rect 14016 8838 14044 11018
rect 14292 10810 14320 11494
rect 14568 11082 14596 12406
rect 14740 12378 14792 12384
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14292 10674 14320 10746
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14108 9926 14136 10610
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14200 9586 14228 10202
rect 14292 10062 14320 10610
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 9602 14504 9862
rect 14568 9722 14596 10610
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14188 9580 14240 9586
rect 14476 9574 14596 9602
rect 14188 9522 14240 9528
rect 14108 9178 14136 9522
rect 14200 9178 14228 9522
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14568 8838 14596 9574
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14016 8537 14044 8774
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14002 8528 14058 8537
rect 14002 8463 14004 8472
rect 14056 8463 14058 8472
rect 14004 8434 14056 8440
rect 14002 8392 14058 8401
rect 14002 8327 14058 8336
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13924 6866 13952 7346
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5710 13768 6054
rect 13832 5710 13860 6666
rect 13924 6390 13952 6666
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 14016 6338 14044 8327
rect 14108 8090 14136 8570
rect 14200 8537 14228 8774
rect 14186 8528 14242 8537
rect 14186 8463 14242 8472
rect 14280 8492 14332 8498
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14200 7993 14228 8463
rect 14280 8434 14332 8440
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14292 8401 14320 8434
rect 14278 8392 14334 8401
rect 14278 8327 14334 8336
rect 14476 8294 14504 8434
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14568 8022 14596 8774
rect 14556 8016 14608 8022
rect 14186 7984 14242 7993
rect 14556 7958 14608 7964
rect 14186 7919 14242 7928
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 13924 6225 13952 6326
rect 14016 6310 14136 6338
rect 14004 6248 14056 6254
rect 13910 6216 13966 6225
rect 14004 6190 14056 6196
rect 13910 6151 13966 6160
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 13188 2582 13216 2926
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13372 2446 13400 2790
rect 13464 2446 13492 3402
rect 13634 3088 13690 3097
rect 13634 3023 13636 3032
rect 13688 3023 13690 3032
rect 13636 2994 13688 3000
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 13740 2378 13768 5510
rect 14016 4554 14044 6190
rect 14108 5166 14136 6310
rect 14200 5273 14228 7346
rect 14292 6866 14320 7822
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14292 6322 14320 6802
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14384 5710 14412 7890
rect 14660 7886 14688 11630
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14476 7721 14504 7822
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14462 7712 14518 7721
rect 14462 7647 14518 7656
rect 14464 7540 14516 7546
rect 14568 7528 14596 7754
rect 14516 7500 14596 7528
rect 14464 7482 14516 7488
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14476 6118 14504 7346
rect 14568 7274 14596 7500
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14568 6798 14596 6938
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6338 14596 6598
rect 14660 6361 14688 7346
rect 14559 6310 14596 6338
rect 14646 6352 14702 6361
rect 14559 6236 14587 6310
rect 14752 6322 14780 12106
rect 14936 11830 14964 12786
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15396 12442 15424 12718
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15028 11082 15056 11698
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 14936 9722 14964 11018
rect 15304 9926 15332 12106
rect 15488 10538 15516 14742
rect 15580 14414 15608 16510
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 16120 16516 16172 16522
rect 16120 16458 16172 16464
rect 15948 16250 15976 16458
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15366 15700 15846
rect 15776 15804 16084 15824
rect 15776 15802 15782 15804
rect 15838 15802 15862 15804
rect 15918 15802 15942 15804
rect 15998 15802 16022 15804
rect 16078 15802 16084 15804
rect 15838 15750 15840 15802
rect 16020 15750 16022 15802
rect 15776 15748 15782 15750
rect 15838 15748 15862 15750
rect 15918 15748 15942 15750
rect 15998 15748 16022 15750
rect 16078 15748 16084 15750
rect 15776 15728 16084 15748
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 16040 14906 16068 15438
rect 16132 15094 16160 16458
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16224 15706 16252 16050
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 16040 14878 16160 14906
rect 16224 14890 16252 15642
rect 16592 15570 16620 16594
rect 16684 16590 16712 16934
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16684 15638 16712 16118
rect 16868 15910 16896 16390
rect 17052 16250 17080 17138
rect 17224 17060 17276 17066
rect 17224 17002 17276 17008
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16672 15632 16724 15638
rect 16672 15574 16724 15580
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 16316 15026 16344 15370
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 15776 14716 16084 14736
rect 15776 14714 15782 14716
rect 15838 14714 15862 14716
rect 15918 14714 15942 14716
rect 15998 14714 16022 14716
rect 16078 14714 16084 14716
rect 15838 14662 15840 14714
rect 16020 14662 16022 14714
rect 15776 14660 15782 14662
rect 15838 14660 15862 14662
rect 15918 14660 15942 14662
rect 15998 14660 16022 14662
rect 16078 14660 16084 14662
rect 15776 14640 16084 14660
rect 16132 14414 16160 14878
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16316 14414 16344 14962
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15580 11150 15608 14214
rect 16592 13938 16620 15506
rect 16684 15094 16712 15574
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 16776 14618 16804 15030
rect 16868 14822 16896 15302
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 15776 13628 16084 13648
rect 15776 13626 15782 13628
rect 15838 13626 15862 13628
rect 15918 13626 15942 13628
rect 15998 13626 16022 13628
rect 16078 13626 16084 13628
rect 15838 13574 15840 13626
rect 16020 13574 16022 13626
rect 15776 13572 15782 13574
rect 15838 13572 15862 13574
rect 15918 13572 15942 13574
rect 15998 13572 16022 13574
rect 16078 13572 16084 13574
rect 15776 13552 16084 13572
rect 16592 13394 16620 13874
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16500 13258 16528 13330
rect 16684 13326 16712 14010
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15672 12238 15700 12786
rect 15948 12714 15976 13126
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 15776 12540 16084 12560
rect 15776 12538 15782 12540
rect 15838 12538 15862 12540
rect 15918 12538 15942 12540
rect 15998 12538 16022 12540
rect 16078 12538 16084 12540
rect 15838 12486 15840 12538
rect 16020 12486 16022 12538
rect 15776 12484 15782 12486
rect 15838 12484 15862 12486
rect 15918 12484 15942 12486
rect 15998 12484 16022 12486
rect 16078 12484 16084 12486
rect 15776 12464 16084 12484
rect 16408 12238 16436 12786
rect 16500 12782 16528 13194
rect 16776 12986 16804 13874
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 15672 11762 15700 12174
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 15776 11452 16084 11472
rect 15776 11450 15782 11452
rect 15838 11450 15862 11452
rect 15918 11450 15942 11452
rect 15998 11450 16022 11452
rect 16078 11450 16084 11452
rect 15838 11398 15840 11450
rect 16020 11398 16022 11450
rect 15776 11396 15782 11398
rect 15838 11396 15862 11398
rect 15918 11396 15942 11398
rect 15998 11396 16022 11398
rect 16078 11396 16084 11398
rect 15776 11376 16084 11396
rect 16132 11354 16160 11630
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16224 11286 16252 12174
rect 16408 11762 16436 12174
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15658 11112 15714 11121
rect 16316 11082 16344 11494
rect 16500 11218 16528 12718
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16684 12306 16712 12582
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16776 11694 16804 12174
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16592 11150 16620 11494
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 15658 11047 15660 11056
rect 15712 11047 15714 11056
rect 16304 11076 16356 11082
rect 15660 11018 15712 11024
rect 16304 11018 16356 11024
rect 16776 10674 16804 11630
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14936 8498 14964 9454
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14936 8090 14964 8434
rect 14924 8084 14976 8090
rect 14844 8044 14924 8072
rect 14646 6287 14702 6296
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14559 6208 14596 6236
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14370 5536 14426 5545
rect 14370 5471 14426 5480
rect 14186 5264 14242 5273
rect 14384 5234 14412 5471
rect 14186 5199 14188 5208
rect 14240 5199 14242 5208
rect 14372 5228 14424 5234
rect 14188 5170 14240 5176
rect 14372 5170 14424 5176
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14108 5030 14136 5102
rect 14200 5098 14228 5170
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14476 5030 14504 6054
rect 14568 5234 14596 6208
rect 14648 5840 14700 5846
rect 14648 5782 14700 5788
rect 14660 5234 14688 5782
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13832 4146 13860 4422
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13832 2650 13860 3470
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13924 2514 13952 3402
rect 14016 3194 14044 4150
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14108 2774 14136 4966
rect 14752 4706 14780 6258
rect 14844 5710 14872 8044
rect 14924 8026 14976 8032
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14936 7750 14964 7822
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 15028 7478 15056 9318
rect 15396 8956 15424 10406
rect 15672 10146 15700 10474
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 15776 10364 16084 10384
rect 15776 10362 15782 10364
rect 15838 10362 15862 10364
rect 15918 10362 15942 10364
rect 15998 10362 16022 10364
rect 16078 10362 16084 10364
rect 15838 10310 15840 10362
rect 16020 10310 16022 10362
rect 15776 10308 15782 10310
rect 15838 10308 15862 10310
rect 15918 10308 15942 10310
rect 15998 10308 16022 10310
rect 16078 10308 16084 10310
rect 15776 10288 16084 10308
rect 15672 10118 15792 10146
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15580 9489 15608 9522
rect 15566 9480 15622 9489
rect 15566 9415 15622 9424
rect 15568 8968 15620 8974
rect 15396 8928 15568 8956
rect 15568 8910 15620 8916
rect 15580 8838 15608 8910
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 14936 7002 14964 7346
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 15028 6866 15056 7278
rect 15120 7206 15148 7346
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15106 7032 15162 7041
rect 15106 6967 15162 6976
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14936 6322 14964 6734
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 15028 6633 15056 6666
rect 15014 6624 15070 6633
rect 15014 6559 15070 6568
rect 15120 6390 15148 6967
rect 15212 6769 15240 8774
rect 15384 7472 15436 7478
rect 15436 7420 15516 7426
rect 15384 7414 15516 7420
rect 15292 7404 15344 7410
rect 15396 7398 15516 7414
rect 15292 7346 15344 7352
rect 15198 6760 15254 6769
rect 15198 6695 15254 6704
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 15304 6225 15332 7346
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 6798 15424 7142
rect 15488 6848 15516 7398
rect 15568 6860 15620 6866
rect 15488 6820 15568 6848
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15382 6624 15438 6633
rect 15382 6559 15438 6568
rect 15290 6216 15346 6225
rect 15290 6151 15346 6160
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15120 5370 15148 5578
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15212 5166 15240 5510
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 14660 4678 14780 4706
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14292 3738 14320 4082
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14384 3738 14412 3878
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14476 3466 14504 4558
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14108 2746 14228 2774
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 12032 2264 12112 2292
rect 11980 2246 12032 2252
rect 11992 2106 12020 2246
rect 11980 2100 12032 2106
rect 11980 2042 12032 2048
rect 12728 1986 12756 2314
rect 12811 2204 13119 2224
rect 12811 2202 12817 2204
rect 12873 2202 12897 2204
rect 12953 2202 12977 2204
rect 13033 2202 13057 2204
rect 13113 2202 13119 2204
rect 12873 2150 12875 2202
rect 13055 2150 13057 2202
rect 12811 2148 12817 2150
rect 12873 2148 12897 2150
rect 12953 2148 12977 2150
rect 13033 2148 13057 2150
rect 13113 2148 13119 2150
rect 12811 2128 13119 2148
rect 14200 2038 14228 2746
rect 14292 2514 14320 3062
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14568 2446 14596 3878
rect 14660 3466 14688 4678
rect 14924 4548 14976 4554
rect 14924 4490 14976 4496
rect 14936 3942 14964 4490
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 14660 2650 14688 3402
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15198 3360 15254 3369
rect 15120 3126 15148 3334
rect 15198 3295 15254 3304
rect 15212 3194 15240 3295
rect 15396 3194 15424 6559
rect 15488 6458 15516 6820
rect 15568 6802 15620 6808
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15580 6390 15608 6666
rect 15672 6662 15700 9862
rect 15764 9586 15792 10118
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15776 9276 16084 9296
rect 15776 9274 15782 9276
rect 15838 9274 15862 9276
rect 15918 9274 15942 9276
rect 15998 9274 16022 9276
rect 16078 9274 16084 9276
rect 15838 9222 15840 9274
rect 16020 9222 16022 9274
rect 15776 9220 15782 9222
rect 15838 9220 15862 9222
rect 15918 9220 15942 9222
rect 15998 9220 16022 9222
rect 16078 9220 16084 9222
rect 15776 9200 16084 9220
rect 16132 8974 16160 10066
rect 16224 9926 16252 10406
rect 16776 10130 16804 10610
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16868 10010 16896 13194
rect 16960 12238 16988 13330
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 17052 12986 17080 13126
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17052 12434 17080 12922
rect 17132 12436 17184 12442
rect 17052 12406 17132 12434
rect 17132 12378 17184 12384
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16776 9982 16896 10010
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16776 9654 16804 9982
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16868 9586 16896 9862
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16960 9450 16988 10610
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 17052 9042 17080 9454
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 15776 8188 16084 8208
rect 15776 8186 15782 8188
rect 15838 8186 15862 8188
rect 15918 8186 15942 8188
rect 15998 8186 16022 8188
rect 16078 8186 16084 8188
rect 15838 8134 15840 8186
rect 16020 8134 16022 8186
rect 15776 8132 15782 8134
rect 15838 8132 15862 8134
rect 15918 8132 15942 8134
rect 15998 8132 16022 8134
rect 16078 8132 16084 8134
rect 15776 8112 16084 8132
rect 16132 7954 16160 8910
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 7970 16252 8774
rect 16408 8090 16436 8910
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16500 8022 16528 8842
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 17052 8566 17080 8774
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 17130 8528 17186 8537
rect 16764 8492 16816 8498
rect 17130 8463 17186 8472
rect 16764 8434 16816 8440
rect 16488 8016 16540 8022
rect 16120 7948 16172 7954
rect 16224 7942 16436 7970
rect 16488 7958 16540 7964
rect 16120 7890 16172 7896
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15776 7100 16084 7120
rect 15776 7098 15782 7100
rect 15838 7098 15862 7100
rect 15918 7098 15942 7100
rect 15998 7098 16022 7100
rect 16078 7098 16084 7100
rect 15838 7046 15840 7098
rect 16020 7046 16022 7098
rect 15776 7044 15782 7046
rect 15838 7044 15862 7046
rect 15918 7044 15942 7046
rect 15998 7044 16022 7046
rect 16078 7044 16084 7046
rect 15776 7024 16084 7044
rect 16132 6798 16160 7142
rect 16224 7002 16252 7346
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16212 6724 16264 6730
rect 16212 6666 16264 6672
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 16224 6322 16252 6666
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 15660 6248 15712 6254
rect 16316 6225 16344 7822
rect 16408 6769 16436 7942
rect 16500 7585 16528 7958
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16486 7576 16542 7585
rect 16486 7511 16542 7520
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16394 6760 16450 6769
rect 16394 6695 16450 6704
rect 16500 6254 16528 7278
rect 16592 6662 16620 7414
rect 16684 6866 16712 7822
rect 16776 7410 16804 8434
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16776 6322 16804 7346
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16868 6662 16896 7142
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16488 6248 16540 6254
rect 15660 6190 15712 6196
rect 16302 6216 16358 6225
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5234 15608 6054
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15672 4622 15700 6190
rect 16488 6190 16540 6196
rect 16302 6151 16358 6160
rect 15776 6012 16084 6032
rect 15776 6010 15782 6012
rect 15838 6010 15862 6012
rect 15918 6010 15942 6012
rect 15998 6010 16022 6012
rect 16078 6010 16084 6012
rect 15838 5958 15840 6010
rect 16020 5958 16022 6010
rect 15776 5956 15782 5958
rect 15838 5956 15862 5958
rect 15918 5956 15942 5958
rect 15998 5956 16022 5958
rect 16078 5956 16084 5958
rect 15776 5936 16084 5956
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16212 5568 16264 5574
rect 16396 5568 16448 5574
rect 16264 5516 16344 5522
rect 16212 5510 16344 5516
rect 16396 5510 16448 5516
rect 16224 5494 16344 5510
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 15776 4924 16084 4944
rect 15776 4922 15782 4924
rect 15838 4922 15862 4924
rect 15918 4922 15942 4924
rect 15998 4922 16022 4924
rect 16078 4922 16084 4924
rect 15838 4870 15840 4922
rect 16020 4870 16022 4922
rect 15776 4868 15782 4870
rect 15838 4868 15862 4870
rect 15918 4868 15942 4870
rect 15998 4868 16022 4870
rect 16078 4868 16084 4870
rect 15776 4848 16084 4868
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 16040 4214 16068 4558
rect 16028 4208 16080 4214
rect 16028 4150 16080 4156
rect 16132 4010 16160 4966
rect 16210 4856 16266 4865
rect 16210 4791 16212 4800
rect 16264 4791 16266 4800
rect 16212 4762 16264 4768
rect 16316 4706 16344 5494
rect 16224 4678 16344 4706
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15108 3120 15160 3126
rect 15396 3097 15424 3130
rect 15108 3062 15160 3068
rect 15382 3088 15438 3097
rect 15382 3023 15438 3032
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 15476 2576 15528 2582
rect 15476 2518 15528 2524
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14188 2032 14240 2038
rect 12728 1958 12940 1986
rect 14188 1974 14240 1980
rect 12912 800 12940 1958
rect 15488 800 15516 2518
rect 5276 734 5488 762
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 15672 762 15700 3946
rect 15776 3836 16084 3856
rect 15776 3834 15782 3836
rect 15838 3834 15862 3836
rect 15918 3834 15942 3836
rect 15998 3834 16022 3836
rect 16078 3834 16084 3836
rect 15838 3782 15840 3834
rect 16020 3782 16022 3834
rect 15776 3780 15782 3782
rect 15838 3780 15862 3782
rect 15918 3780 15942 3782
rect 15998 3780 16022 3782
rect 16078 3780 16084 3782
rect 15776 3760 16084 3780
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 15776 2748 16084 2768
rect 15776 2746 15782 2748
rect 15838 2746 15862 2748
rect 15918 2746 15942 2748
rect 15998 2746 16022 2748
rect 16078 2746 16084 2748
rect 15838 2694 15840 2746
rect 16020 2694 16022 2746
rect 15776 2692 15782 2694
rect 15838 2692 15862 2694
rect 15918 2692 15942 2694
rect 15998 2692 16022 2694
rect 16078 2692 16084 2694
rect 15776 2672 16084 2692
rect 16132 2145 16160 3470
rect 16224 2446 16252 4678
rect 16408 4622 16436 5510
rect 16684 5370 16712 5646
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16776 5234 16804 6258
rect 16960 5778 16988 6802
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 17144 5710 17172 8463
rect 17236 7886 17264 17002
rect 17420 16046 17448 19200
rect 18064 17338 18092 19200
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17512 16114 17540 16390
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17328 15162 17356 15370
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17604 12434 17632 17138
rect 17682 17096 17738 17105
rect 17682 17031 17684 17040
rect 17736 17031 17738 17040
rect 17684 17002 17736 17008
rect 18064 16017 18092 17138
rect 18050 16008 18106 16017
rect 18050 15943 18106 15952
rect 18326 15736 18382 15745
rect 18326 15671 18382 15680
rect 17866 15056 17922 15065
rect 18340 15026 18368 15671
rect 17866 14991 17922 15000
rect 18328 15020 18380 15026
rect 17880 14618 17908 14991
rect 18328 14962 18380 14968
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 18328 14408 18380 14414
rect 18326 14376 18328 14385
rect 18380 14376 18382 14385
rect 18236 14340 18288 14346
rect 18326 14311 18382 14320
rect 18236 14282 18288 14288
rect 18248 13530 18276 14282
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18234 13016 18290 13025
rect 18234 12951 18236 12960
rect 18288 12951 18290 12960
rect 18236 12922 18288 12928
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17512 12406 17632 12434
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17328 9722 17356 9930
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16486 5128 16542 5137
rect 16486 5063 16542 5072
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 16316 3126 16344 4150
rect 16500 3670 16528 5063
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16592 3058 16620 4558
rect 16776 4554 16804 5170
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16684 4146 16712 4422
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16776 3058 16804 4490
rect 16960 4282 16988 5170
rect 17316 4548 17368 4554
rect 17316 4490 17368 4496
rect 17328 4282 17356 4490
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 17420 4146 17448 9522
rect 17512 9058 17540 12406
rect 17788 11558 17816 12786
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17604 9654 17632 11018
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17776 10056 17828 10062
rect 17880 10044 17908 10950
rect 18064 10266 18092 12786
rect 18326 11656 18382 11665
rect 18326 11591 18382 11600
rect 18340 11150 18368 11591
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17828 10016 17908 10044
rect 17776 9998 17828 10004
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17512 9030 17632 9058
rect 17500 8968 17552 8974
rect 17498 8936 17500 8945
rect 17552 8936 17554 8945
rect 17498 8871 17554 8880
rect 17500 8288 17552 8294
rect 17604 8276 17632 9030
rect 17696 8634 17724 9318
rect 17788 9178 17816 9454
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17552 8248 17632 8276
rect 17500 8230 17552 8236
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17788 6905 17816 7822
rect 17774 6896 17830 6905
rect 17774 6831 17830 6840
rect 17880 6730 17908 10016
rect 17958 9616 18014 9625
rect 17958 9551 17960 9560
rect 18012 9551 18014 9560
rect 17960 9522 18012 9528
rect 17958 9480 18014 9489
rect 17958 9415 18014 9424
rect 17972 8974 18000 9415
rect 18064 8974 18092 10202
rect 18236 9648 18288 9654
rect 18234 9616 18236 9625
rect 18288 9616 18290 9625
rect 18234 9551 18290 9560
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18156 7750 18184 8230
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 18248 6458 18276 6734
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17512 4865 17540 5646
rect 17498 4856 17554 4865
rect 17498 4791 17554 4800
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18234 4176 18290 4185
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17684 4140 17736 4146
rect 18340 4146 18368 4422
rect 18234 4111 18290 4120
rect 18328 4140 18380 4146
rect 17684 4082 17736 4088
rect 16856 4072 16908 4078
rect 17696 4049 17724 4082
rect 17776 4072 17828 4078
rect 16856 4014 16908 4020
rect 17682 4040 17738 4049
rect 16868 3738 16896 4014
rect 17776 4014 17828 4020
rect 17682 3975 17738 3984
rect 17788 3738 17816 4014
rect 18248 4010 18276 4111
rect 18328 4082 18380 4088
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 18340 3602 18368 4082
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 17040 3528 17092 3534
rect 17038 3496 17040 3505
rect 17132 3528 17184 3534
rect 17092 3496 17094 3505
rect 17132 3470 17184 3476
rect 17038 3431 17094 3440
rect 17144 3194 17172 3470
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 17144 2446 17172 3130
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16118 2136 16174 2145
rect 16118 2071 16174 2080
rect 16040 870 16160 898
rect 16040 762 16068 870
rect 16132 800 16160 870
rect 16776 800 16804 2246
rect 15672 734 16068 762
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17696 785 17724 2382
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 800 18092 2246
rect 18708 800 18736 3878
rect 17682 776 17738 785
rect 17682 711 17738 720
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
<< via2 >>
rect 2778 19080 2834 19136
rect 2226 17720 2282 17776
rect 1398 17040 1454 17096
rect 1398 15020 1454 15056
rect 1398 15000 1400 15020
rect 1400 15000 1452 15020
rect 1452 15000 1454 15020
rect 1398 14356 1400 14376
rect 1400 14356 1452 14376
rect 1452 14356 1454 14376
rect 1398 14320 1454 14356
rect 1398 11620 1454 11656
rect 1398 11600 1400 11620
rect 1400 11600 1452 11620
rect 1452 11600 1454 11620
rect 1398 10920 1454 10976
rect 1398 9560 1454 9616
rect 1490 8880 1546 8936
rect 1398 6860 1454 6896
rect 1398 6840 1400 6860
rect 1400 6840 1452 6860
rect 1452 6840 1454 6860
rect 1398 6196 1400 6216
rect 1400 6196 1452 6216
rect 1452 6196 1454 6216
rect 1398 6160 1454 6196
rect 6886 17434 6942 17436
rect 6966 17434 7022 17436
rect 7046 17434 7102 17436
rect 7126 17434 7182 17436
rect 6886 17382 6932 17434
rect 6932 17382 6942 17434
rect 6966 17382 6996 17434
rect 6996 17382 7008 17434
rect 7008 17382 7022 17434
rect 7046 17382 7060 17434
rect 7060 17382 7072 17434
rect 7072 17382 7102 17434
rect 7126 17382 7136 17434
rect 7136 17382 7182 17434
rect 6886 17380 6942 17382
rect 6966 17380 7022 17382
rect 7046 17380 7102 17382
rect 7126 17380 7182 17382
rect 3921 16890 3977 16892
rect 4001 16890 4057 16892
rect 4081 16890 4137 16892
rect 4161 16890 4217 16892
rect 3921 16838 3967 16890
rect 3967 16838 3977 16890
rect 4001 16838 4031 16890
rect 4031 16838 4043 16890
rect 4043 16838 4057 16890
rect 4081 16838 4095 16890
rect 4095 16838 4107 16890
rect 4107 16838 4137 16890
rect 4161 16838 4171 16890
rect 4171 16838 4217 16890
rect 3921 16836 3977 16838
rect 4001 16836 4057 16838
rect 4081 16836 4137 16838
rect 4161 16836 4217 16838
rect 3921 15802 3977 15804
rect 4001 15802 4057 15804
rect 4081 15802 4137 15804
rect 4161 15802 4217 15804
rect 3921 15750 3967 15802
rect 3967 15750 3977 15802
rect 4001 15750 4031 15802
rect 4031 15750 4043 15802
rect 4043 15750 4057 15802
rect 4081 15750 4095 15802
rect 4095 15750 4107 15802
rect 4107 15750 4137 15802
rect 4161 15750 4171 15802
rect 4171 15750 4217 15802
rect 3921 15748 3977 15750
rect 4001 15748 4057 15750
rect 4081 15748 4137 15750
rect 4161 15748 4217 15750
rect 3921 14714 3977 14716
rect 4001 14714 4057 14716
rect 4081 14714 4137 14716
rect 4161 14714 4217 14716
rect 3921 14662 3967 14714
rect 3967 14662 3977 14714
rect 4001 14662 4031 14714
rect 4031 14662 4043 14714
rect 4043 14662 4057 14714
rect 4081 14662 4095 14714
rect 4095 14662 4107 14714
rect 4107 14662 4137 14714
rect 4161 14662 4171 14714
rect 4171 14662 4217 14714
rect 3921 14660 3977 14662
rect 4001 14660 4057 14662
rect 4081 14660 4137 14662
rect 4161 14660 4217 14662
rect 7194 16632 7250 16688
rect 12817 17434 12873 17436
rect 12897 17434 12953 17436
rect 12977 17434 13033 17436
rect 13057 17434 13113 17436
rect 12817 17382 12863 17434
rect 12863 17382 12873 17434
rect 12897 17382 12927 17434
rect 12927 17382 12939 17434
rect 12939 17382 12953 17434
rect 12977 17382 12991 17434
rect 12991 17382 13003 17434
rect 13003 17382 13033 17434
rect 13057 17382 13067 17434
rect 13067 17382 13113 17434
rect 12817 17380 12873 17382
rect 12897 17380 12953 17382
rect 12977 17380 13033 17382
rect 13057 17380 13113 17382
rect 6886 16346 6942 16348
rect 6966 16346 7022 16348
rect 7046 16346 7102 16348
rect 7126 16346 7182 16348
rect 6886 16294 6932 16346
rect 6932 16294 6942 16346
rect 6966 16294 6996 16346
rect 6996 16294 7008 16346
rect 7008 16294 7022 16346
rect 7046 16294 7060 16346
rect 7060 16294 7072 16346
rect 7072 16294 7102 16346
rect 7126 16294 7136 16346
rect 7136 16294 7182 16346
rect 6886 16292 6942 16294
rect 6966 16292 7022 16294
rect 7046 16292 7102 16294
rect 7126 16292 7182 16294
rect 6886 15258 6942 15260
rect 6966 15258 7022 15260
rect 7046 15258 7102 15260
rect 7126 15258 7182 15260
rect 6886 15206 6932 15258
rect 6932 15206 6942 15258
rect 6966 15206 6996 15258
rect 6996 15206 7008 15258
rect 7008 15206 7022 15258
rect 7046 15206 7060 15258
rect 7060 15206 7072 15258
rect 7072 15206 7102 15258
rect 7126 15206 7136 15258
rect 7136 15206 7182 15258
rect 6886 15204 6942 15206
rect 6966 15204 7022 15206
rect 7046 15204 7102 15206
rect 7126 15204 7182 15206
rect 3921 13626 3977 13628
rect 4001 13626 4057 13628
rect 4081 13626 4137 13628
rect 4161 13626 4217 13628
rect 3921 13574 3967 13626
rect 3967 13574 3977 13626
rect 4001 13574 4031 13626
rect 4031 13574 4043 13626
rect 4043 13574 4057 13626
rect 4081 13574 4095 13626
rect 4095 13574 4107 13626
rect 4107 13574 4137 13626
rect 4161 13574 4171 13626
rect 4171 13574 4217 13626
rect 3921 13572 3977 13574
rect 4001 13572 4057 13574
rect 4081 13572 4137 13574
rect 4161 13572 4217 13574
rect 3921 12538 3977 12540
rect 4001 12538 4057 12540
rect 4081 12538 4137 12540
rect 4161 12538 4217 12540
rect 3921 12486 3967 12538
rect 3967 12486 3977 12538
rect 4001 12486 4031 12538
rect 4031 12486 4043 12538
rect 4043 12486 4057 12538
rect 4081 12486 4095 12538
rect 4095 12486 4107 12538
rect 4107 12486 4137 12538
rect 4161 12486 4171 12538
rect 4171 12486 4217 12538
rect 3921 12484 3977 12486
rect 4001 12484 4057 12486
rect 4081 12484 4137 12486
rect 4161 12484 4217 12486
rect 3921 11450 3977 11452
rect 4001 11450 4057 11452
rect 4081 11450 4137 11452
rect 4161 11450 4217 11452
rect 3921 11398 3967 11450
rect 3967 11398 3977 11450
rect 4001 11398 4031 11450
rect 4031 11398 4043 11450
rect 4043 11398 4057 11450
rect 4081 11398 4095 11450
rect 4095 11398 4107 11450
rect 4107 11398 4137 11450
rect 4161 11398 4171 11450
rect 4171 11398 4217 11450
rect 3921 11396 3977 11398
rect 4001 11396 4057 11398
rect 4081 11396 4137 11398
rect 4161 11396 4217 11398
rect 3921 10362 3977 10364
rect 4001 10362 4057 10364
rect 4081 10362 4137 10364
rect 4161 10362 4217 10364
rect 3921 10310 3967 10362
rect 3967 10310 3977 10362
rect 4001 10310 4031 10362
rect 4031 10310 4043 10362
rect 4043 10310 4057 10362
rect 4081 10310 4095 10362
rect 4095 10310 4107 10362
rect 4107 10310 4137 10362
rect 4161 10310 4171 10362
rect 4171 10310 4217 10362
rect 3921 10308 3977 10310
rect 4001 10308 4057 10310
rect 4081 10308 4137 10310
rect 4161 10308 4217 10310
rect 3054 10104 3110 10160
rect 6734 14592 6790 14648
rect 7102 14728 7158 14784
rect 7010 14356 7012 14376
rect 7012 14356 7064 14376
rect 7064 14356 7066 14376
rect 7010 14320 7066 14356
rect 7286 14476 7342 14512
rect 7286 14456 7288 14476
rect 7288 14456 7340 14476
rect 7340 14456 7342 14476
rect 6886 14170 6942 14172
rect 6966 14170 7022 14172
rect 7046 14170 7102 14172
rect 7126 14170 7182 14172
rect 6886 14118 6932 14170
rect 6932 14118 6942 14170
rect 6966 14118 6996 14170
rect 6996 14118 7008 14170
rect 7008 14118 7022 14170
rect 7046 14118 7060 14170
rect 7060 14118 7072 14170
rect 7072 14118 7102 14170
rect 7126 14118 7136 14170
rect 7136 14118 7182 14170
rect 6886 14116 6942 14118
rect 6966 14116 7022 14118
rect 7046 14116 7102 14118
rect 7126 14116 7182 14118
rect 6886 13082 6942 13084
rect 6966 13082 7022 13084
rect 7046 13082 7102 13084
rect 7126 13082 7182 13084
rect 6886 13030 6932 13082
rect 6932 13030 6942 13082
rect 6966 13030 6996 13082
rect 6996 13030 7008 13082
rect 7008 13030 7022 13082
rect 7046 13030 7060 13082
rect 7060 13030 7072 13082
rect 7072 13030 7102 13082
rect 7126 13030 7136 13082
rect 7136 13030 7182 13082
rect 6886 13028 6942 13030
rect 6966 13028 7022 13030
rect 7046 13028 7102 13030
rect 7126 13028 7182 13030
rect 7654 15952 7710 16008
rect 6886 11994 6942 11996
rect 6966 11994 7022 11996
rect 7046 11994 7102 11996
rect 7126 11994 7182 11996
rect 6886 11942 6932 11994
rect 6932 11942 6942 11994
rect 6966 11942 6996 11994
rect 6996 11942 7008 11994
rect 7008 11942 7022 11994
rect 7046 11942 7060 11994
rect 7060 11942 7072 11994
rect 7072 11942 7102 11994
rect 7126 11942 7136 11994
rect 7136 11942 7182 11994
rect 6886 11940 6942 11942
rect 6966 11940 7022 11942
rect 7046 11940 7102 11942
rect 7126 11940 7182 11942
rect 8482 14728 8538 14784
rect 7746 14356 7748 14376
rect 7748 14356 7800 14376
rect 7800 14356 7802 14376
rect 7746 14320 7802 14356
rect 8942 14592 8998 14648
rect 3921 9274 3977 9276
rect 4001 9274 4057 9276
rect 4081 9274 4137 9276
rect 4161 9274 4217 9276
rect 3921 9222 3967 9274
rect 3967 9222 3977 9274
rect 4001 9222 4031 9274
rect 4031 9222 4043 9274
rect 4043 9222 4057 9274
rect 4081 9222 4095 9274
rect 4095 9222 4107 9274
rect 4107 9222 4137 9274
rect 4161 9222 4171 9274
rect 4171 9222 4217 9274
rect 3921 9220 3977 9222
rect 4001 9220 4057 9222
rect 4081 9220 4137 9222
rect 4161 9220 4217 9222
rect 4434 8880 4490 8936
rect 3921 8186 3977 8188
rect 4001 8186 4057 8188
rect 4081 8186 4137 8188
rect 4161 8186 4217 8188
rect 3921 8134 3967 8186
rect 3967 8134 3977 8186
rect 4001 8134 4031 8186
rect 4031 8134 4043 8186
rect 4043 8134 4057 8186
rect 4081 8134 4095 8186
rect 4095 8134 4107 8186
rect 4107 8134 4137 8186
rect 4161 8134 4171 8186
rect 4171 8134 4217 8186
rect 3921 8132 3977 8134
rect 4001 8132 4057 8134
rect 4081 8132 4137 8134
rect 4161 8132 4217 8134
rect 2502 6840 2558 6896
rect 3921 7098 3977 7100
rect 4001 7098 4057 7100
rect 4081 7098 4137 7100
rect 4161 7098 4217 7100
rect 3921 7046 3967 7098
rect 3967 7046 3977 7098
rect 4001 7046 4031 7098
rect 4031 7046 4043 7098
rect 4043 7046 4057 7098
rect 4081 7046 4095 7098
rect 4095 7046 4107 7098
rect 4107 7046 4137 7098
rect 4161 7046 4171 7098
rect 4171 7046 4217 7098
rect 3921 7044 3977 7046
rect 4001 7044 4057 7046
rect 4081 7044 4137 7046
rect 4161 7044 4217 7046
rect 2226 2760 2282 2816
rect 3921 6010 3977 6012
rect 4001 6010 4057 6012
rect 4081 6010 4137 6012
rect 4161 6010 4217 6012
rect 3921 5958 3967 6010
rect 3967 5958 3977 6010
rect 4001 5958 4031 6010
rect 4031 5958 4043 6010
rect 4043 5958 4057 6010
rect 4081 5958 4095 6010
rect 4095 5958 4107 6010
rect 4107 5958 4137 6010
rect 4161 5958 4171 6010
rect 4171 5958 4217 6010
rect 3921 5956 3977 5958
rect 4001 5956 4057 5958
rect 4081 5956 4137 5958
rect 4161 5956 4217 5958
rect 3921 4922 3977 4924
rect 4001 4922 4057 4924
rect 4081 4922 4137 4924
rect 4161 4922 4217 4924
rect 3921 4870 3967 4922
rect 3967 4870 3977 4922
rect 4001 4870 4031 4922
rect 4031 4870 4043 4922
rect 4043 4870 4057 4922
rect 4081 4870 4095 4922
rect 4095 4870 4107 4922
rect 4107 4870 4137 4922
rect 4161 4870 4171 4922
rect 4171 4870 4217 4922
rect 3921 4868 3977 4870
rect 4001 4868 4057 4870
rect 4081 4868 4137 4870
rect 4161 4868 4217 4870
rect 3921 3834 3977 3836
rect 4001 3834 4057 3836
rect 4081 3834 4137 3836
rect 4161 3834 4217 3836
rect 3921 3782 3967 3834
rect 3967 3782 3977 3834
rect 4001 3782 4031 3834
rect 4031 3782 4043 3834
rect 4043 3782 4057 3834
rect 4081 3782 4095 3834
rect 4095 3782 4107 3834
rect 4107 3782 4137 3834
rect 4161 3782 4171 3834
rect 4171 3782 4217 3834
rect 3921 3780 3977 3782
rect 4001 3780 4057 3782
rect 4081 3780 4137 3782
rect 4161 3780 4217 3782
rect 5170 8472 5226 8528
rect 5170 6296 5226 6352
rect 6886 10906 6942 10908
rect 6966 10906 7022 10908
rect 7046 10906 7102 10908
rect 7126 10906 7182 10908
rect 6886 10854 6932 10906
rect 6932 10854 6942 10906
rect 6966 10854 6996 10906
rect 6996 10854 7008 10906
rect 7008 10854 7022 10906
rect 7046 10854 7060 10906
rect 7060 10854 7072 10906
rect 7072 10854 7102 10906
rect 7126 10854 7136 10906
rect 7136 10854 7182 10906
rect 6886 10852 6942 10854
rect 6966 10852 7022 10854
rect 7046 10852 7102 10854
rect 7126 10852 7182 10854
rect 6886 9818 6942 9820
rect 6966 9818 7022 9820
rect 7046 9818 7102 9820
rect 7126 9818 7182 9820
rect 6886 9766 6932 9818
rect 6932 9766 6942 9818
rect 6966 9766 6996 9818
rect 6996 9766 7008 9818
rect 7008 9766 7022 9818
rect 7046 9766 7060 9818
rect 7060 9766 7072 9818
rect 7072 9766 7102 9818
rect 7126 9766 7136 9818
rect 7136 9766 7182 9818
rect 6886 9764 6942 9766
rect 6966 9764 7022 9766
rect 7046 9764 7102 9766
rect 7126 9764 7182 9766
rect 9218 15972 9274 16008
rect 9218 15952 9220 15972
rect 9220 15952 9272 15972
rect 9272 15952 9274 15972
rect 9852 16890 9908 16892
rect 9932 16890 9988 16892
rect 10012 16890 10068 16892
rect 10092 16890 10148 16892
rect 9852 16838 9898 16890
rect 9898 16838 9908 16890
rect 9932 16838 9962 16890
rect 9962 16838 9974 16890
rect 9974 16838 9988 16890
rect 10012 16838 10026 16890
rect 10026 16838 10038 16890
rect 10038 16838 10068 16890
rect 10092 16838 10102 16890
rect 10102 16838 10148 16890
rect 9852 16836 9908 16838
rect 9932 16836 9988 16838
rect 10012 16836 10068 16838
rect 10092 16836 10148 16838
rect 9852 15802 9908 15804
rect 9932 15802 9988 15804
rect 10012 15802 10068 15804
rect 10092 15802 10148 15804
rect 9852 15750 9898 15802
rect 9898 15750 9908 15802
rect 9932 15750 9962 15802
rect 9962 15750 9974 15802
rect 9974 15750 9988 15802
rect 10012 15750 10026 15802
rect 10026 15750 10038 15802
rect 10038 15750 10068 15802
rect 10092 15750 10102 15802
rect 10102 15750 10148 15802
rect 9852 15748 9908 15750
rect 9932 15748 9988 15750
rect 10012 15748 10068 15750
rect 10092 15748 10148 15750
rect 9852 14714 9908 14716
rect 9932 14714 9988 14716
rect 10012 14714 10068 14716
rect 10092 14714 10148 14716
rect 9852 14662 9898 14714
rect 9898 14662 9908 14714
rect 9932 14662 9962 14714
rect 9962 14662 9974 14714
rect 9974 14662 9988 14714
rect 10012 14662 10026 14714
rect 10026 14662 10038 14714
rect 10038 14662 10068 14714
rect 10092 14662 10102 14714
rect 10102 14662 10148 14714
rect 9852 14660 9908 14662
rect 9932 14660 9988 14662
rect 10012 14660 10068 14662
rect 10092 14660 10148 14662
rect 10138 14492 10140 14512
rect 10140 14492 10192 14512
rect 10192 14492 10194 14512
rect 10138 14456 10194 14492
rect 9852 13626 9908 13628
rect 9932 13626 9988 13628
rect 10012 13626 10068 13628
rect 10092 13626 10148 13628
rect 9852 13574 9898 13626
rect 9898 13574 9908 13626
rect 9932 13574 9962 13626
rect 9962 13574 9974 13626
rect 9974 13574 9988 13626
rect 10012 13574 10026 13626
rect 10026 13574 10038 13626
rect 10038 13574 10068 13626
rect 10092 13574 10102 13626
rect 10102 13574 10148 13626
rect 9852 13572 9908 13574
rect 9932 13572 9988 13574
rect 10012 13572 10068 13574
rect 10092 13572 10148 13574
rect 9852 12538 9908 12540
rect 9932 12538 9988 12540
rect 10012 12538 10068 12540
rect 10092 12538 10148 12540
rect 9852 12486 9898 12538
rect 9898 12486 9908 12538
rect 9932 12486 9962 12538
rect 9962 12486 9974 12538
rect 9974 12486 9988 12538
rect 10012 12486 10026 12538
rect 10026 12486 10038 12538
rect 10038 12486 10068 12538
rect 10092 12486 10102 12538
rect 10102 12486 10148 12538
rect 9852 12484 9908 12486
rect 9932 12484 9988 12486
rect 10012 12484 10068 12486
rect 10092 12484 10148 12486
rect 6886 8730 6942 8732
rect 6966 8730 7022 8732
rect 7046 8730 7102 8732
rect 7126 8730 7182 8732
rect 6886 8678 6932 8730
rect 6932 8678 6942 8730
rect 6966 8678 6996 8730
rect 6996 8678 7008 8730
rect 7008 8678 7022 8730
rect 7046 8678 7060 8730
rect 7060 8678 7072 8730
rect 7072 8678 7102 8730
rect 7126 8678 7136 8730
rect 7136 8678 7182 8730
rect 6886 8676 6942 8678
rect 6966 8676 7022 8678
rect 7046 8676 7102 8678
rect 7126 8676 7182 8678
rect 6886 7642 6942 7644
rect 6966 7642 7022 7644
rect 7046 7642 7102 7644
rect 7126 7642 7182 7644
rect 6886 7590 6932 7642
rect 6932 7590 6942 7642
rect 6966 7590 6996 7642
rect 6996 7590 7008 7642
rect 7008 7590 7022 7642
rect 7046 7590 7060 7642
rect 7060 7590 7072 7642
rect 7072 7590 7102 7642
rect 7126 7590 7136 7642
rect 7136 7590 7182 7642
rect 6886 7588 6942 7590
rect 6966 7588 7022 7590
rect 7046 7588 7102 7590
rect 7126 7588 7182 7590
rect 3921 2746 3977 2748
rect 4001 2746 4057 2748
rect 4081 2746 4137 2748
rect 4161 2746 4217 2748
rect 3921 2694 3967 2746
rect 3967 2694 3977 2746
rect 4001 2694 4031 2746
rect 4031 2694 4043 2746
rect 4043 2694 4057 2746
rect 4081 2694 4095 2746
rect 4095 2694 4107 2746
rect 4107 2694 4137 2746
rect 4161 2694 4171 2746
rect 4171 2694 4217 2746
rect 3921 2692 3977 2694
rect 4001 2692 4057 2694
rect 4081 2692 4137 2694
rect 4161 2692 4217 2694
rect 7838 7948 7894 7984
rect 7838 7928 7840 7948
rect 7840 7928 7892 7948
rect 7892 7928 7894 7948
rect 6886 6554 6942 6556
rect 6966 6554 7022 6556
rect 7046 6554 7102 6556
rect 7126 6554 7182 6556
rect 6886 6502 6932 6554
rect 6932 6502 6942 6554
rect 6966 6502 6996 6554
rect 6996 6502 7008 6554
rect 7008 6502 7022 6554
rect 7046 6502 7060 6554
rect 7060 6502 7072 6554
rect 7072 6502 7102 6554
rect 7126 6502 7136 6554
rect 7136 6502 7182 6554
rect 6886 6500 6942 6502
rect 6966 6500 7022 6502
rect 7046 6500 7102 6502
rect 7126 6500 7182 6502
rect 6886 5466 6942 5468
rect 6966 5466 7022 5468
rect 7046 5466 7102 5468
rect 7126 5466 7182 5468
rect 6886 5414 6932 5466
rect 6932 5414 6942 5466
rect 6966 5414 6996 5466
rect 6996 5414 7008 5466
rect 7008 5414 7022 5466
rect 7046 5414 7060 5466
rect 7060 5414 7072 5466
rect 7072 5414 7102 5466
rect 7126 5414 7136 5466
rect 7136 5414 7182 5466
rect 6886 5412 6942 5414
rect 6966 5412 7022 5414
rect 7046 5412 7102 5414
rect 7126 5412 7182 5414
rect 8114 6704 8170 6760
rect 6886 4378 6942 4380
rect 6966 4378 7022 4380
rect 7046 4378 7102 4380
rect 7126 4378 7182 4380
rect 6886 4326 6932 4378
rect 6932 4326 6942 4378
rect 6966 4326 6996 4378
rect 6996 4326 7008 4378
rect 7008 4326 7022 4378
rect 7046 4326 7060 4378
rect 7060 4326 7072 4378
rect 7072 4326 7102 4378
rect 7126 4326 7136 4378
rect 7136 4326 7182 4378
rect 6886 4324 6942 4326
rect 6966 4324 7022 4326
rect 7046 4324 7102 4326
rect 7126 4324 7182 4326
rect 6886 3290 6942 3292
rect 6966 3290 7022 3292
rect 7046 3290 7102 3292
rect 7126 3290 7182 3292
rect 6886 3238 6932 3290
rect 6932 3238 6942 3290
rect 6966 3238 6996 3290
rect 6996 3238 7008 3290
rect 7008 3238 7022 3290
rect 7046 3238 7060 3290
rect 7060 3238 7072 3290
rect 7072 3238 7102 3290
rect 7126 3238 7136 3290
rect 7136 3238 7182 3290
rect 6886 3236 6942 3238
rect 6966 3236 7022 3238
rect 7046 3236 7102 3238
rect 7126 3236 7182 3238
rect 3422 1400 3478 1456
rect 2778 720 2834 776
rect 6886 2202 6942 2204
rect 6966 2202 7022 2204
rect 7046 2202 7102 2204
rect 7126 2202 7182 2204
rect 6886 2150 6932 2202
rect 6932 2150 6942 2202
rect 6966 2150 6996 2202
rect 6996 2150 7008 2202
rect 7008 2150 7022 2202
rect 7046 2150 7060 2202
rect 7060 2150 7072 2202
rect 7072 2150 7102 2202
rect 7126 2150 7136 2202
rect 7136 2150 7182 2202
rect 6886 2148 6942 2150
rect 6966 2148 7022 2150
rect 7046 2148 7102 2150
rect 7126 2148 7182 2150
rect 9852 11450 9908 11452
rect 9932 11450 9988 11452
rect 10012 11450 10068 11452
rect 10092 11450 10148 11452
rect 9852 11398 9898 11450
rect 9898 11398 9908 11450
rect 9932 11398 9962 11450
rect 9962 11398 9974 11450
rect 9974 11398 9988 11450
rect 10012 11398 10026 11450
rect 10026 11398 10038 11450
rect 10038 11398 10068 11450
rect 10092 11398 10102 11450
rect 10102 11398 10148 11450
rect 9852 11396 9908 11398
rect 9932 11396 9988 11398
rect 10012 11396 10068 11398
rect 10092 11396 10148 11398
rect 9852 10362 9908 10364
rect 9932 10362 9988 10364
rect 10012 10362 10068 10364
rect 10092 10362 10148 10364
rect 9852 10310 9898 10362
rect 9898 10310 9908 10362
rect 9932 10310 9962 10362
rect 9962 10310 9974 10362
rect 9974 10310 9988 10362
rect 10012 10310 10026 10362
rect 10026 10310 10038 10362
rect 10038 10310 10068 10362
rect 10092 10310 10102 10362
rect 10102 10310 10148 10362
rect 9852 10308 9908 10310
rect 9932 10308 9988 10310
rect 10012 10308 10068 10310
rect 10092 10308 10148 10310
rect 9852 9274 9908 9276
rect 9932 9274 9988 9276
rect 10012 9274 10068 9276
rect 10092 9274 10148 9276
rect 9852 9222 9898 9274
rect 9898 9222 9908 9274
rect 9932 9222 9962 9274
rect 9962 9222 9974 9274
rect 9974 9222 9988 9274
rect 10012 9222 10026 9274
rect 10026 9222 10038 9274
rect 10038 9222 10068 9274
rect 10092 9222 10102 9274
rect 10102 9222 10148 9274
rect 9852 9220 9908 9222
rect 9932 9220 9988 9222
rect 10012 9220 10068 9222
rect 10092 9220 10148 9222
rect 9852 8186 9908 8188
rect 9932 8186 9988 8188
rect 10012 8186 10068 8188
rect 10092 8186 10148 8188
rect 9852 8134 9898 8186
rect 9898 8134 9908 8186
rect 9932 8134 9962 8186
rect 9962 8134 9974 8186
rect 9974 8134 9988 8186
rect 10012 8134 10026 8186
rect 10026 8134 10038 8186
rect 10038 8134 10068 8186
rect 10092 8134 10102 8186
rect 10102 8134 10148 8186
rect 9852 8132 9908 8134
rect 9932 8132 9988 8134
rect 10012 8132 10068 8134
rect 10092 8132 10148 8134
rect 9852 7098 9908 7100
rect 9932 7098 9988 7100
rect 10012 7098 10068 7100
rect 10092 7098 10148 7100
rect 9852 7046 9898 7098
rect 9898 7046 9908 7098
rect 9932 7046 9962 7098
rect 9962 7046 9974 7098
rect 9974 7046 9988 7098
rect 10012 7046 10026 7098
rect 10026 7046 10038 7098
rect 10038 7046 10068 7098
rect 10092 7046 10102 7098
rect 10102 7046 10148 7098
rect 9852 7044 9908 7046
rect 9932 7044 9988 7046
rect 10012 7044 10068 7046
rect 10092 7044 10148 7046
rect 10782 16088 10838 16144
rect 12817 16346 12873 16348
rect 12897 16346 12953 16348
rect 12977 16346 13033 16348
rect 13057 16346 13113 16348
rect 12817 16294 12863 16346
rect 12863 16294 12873 16346
rect 12897 16294 12927 16346
rect 12927 16294 12939 16346
rect 12939 16294 12953 16346
rect 12977 16294 12991 16346
rect 12991 16294 13003 16346
rect 13003 16294 13033 16346
rect 13057 16294 13067 16346
rect 13067 16294 13113 16346
rect 12817 16292 12873 16294
rect 12897 16292 12953 16294
rect 12977 16292 13033 16294
rect 13057 16292 13113 16294
rect 12622 16088 12678 16144
rect 12990 16088 13046 16144
rect 12817 15258 12873 15260
rect 12897 15258 12953 15260
rect 12977 15258 13033 15260
rect 13057 15258 13113 15260
rect 12817 15206 12863 15258
rect 12863 15206 12873 15258
rect 12897 15206 12927 15258
rect 12927 15206 12939 15258
rect 12939 15206 12953 15258
rect 12977 15206 12991 15258
rect 12991 15206 13003 15258
rect 13003 15206 13033 15258
rect 13057 15206 13067 15258
rect 13067 15206 13113 15258
rect 12817 15204 12873 15206
rect 12897 15204 12953 15206
rect 12977 15204 13033 15206
rect 13057 15204 13113 15206
rect 10690 12844 10746 12880
rect 10690 12824 10692 12844
rect 10692 12824 10744 12844
rect 10744 12824 10746 12844
rect 10874 9016 10930 9072
rect 10690 7656 10746 7712
rect 9852 6010 9908 6012
rect 9932 6010 9988 6012
rect 10012 6010 10068 6012
rect 10092 6010 10148 6012
rect 9852 5958 9898 6010
rect 9898 5958 9908 6010
rect 9932 5958 9962 6010
rect 9962 5958 9974 6010
rect 9974 5958 9988 6010
rect 10012 5958 10026 6010
rect 10026 5958 10038 6010
rect 10038 5958 10068 6010
rect 10092 5958 10102 6010
rect 10102 5958 10148 6010
rect 9852 5956 9908 5958
rect 9932 5956 9988 5958
rect 10012 5956 10068 5958
rect 10092 5956 10148 5958
rect 10506 6568 10562 6624
rect 10506 5344 10562 5400
rect 9954 5072 10010 5128
rect 9852 4922 9908 4924
rect 9932 4922 9988 4924
rect 10012 4922 10068 4924
rect 10092 4922 10148 4924
rect 9852 4870 9898 4922
rect 9898 4870 9908 4922
rect 9932 4870 9962 4922
rect 9962 4870 9974 4922
rect 9974 4870 9988 4922
rect 10012 4870 10026 4922
rect 10026 4870 10038 4922
rect 10038 4870 10068 4922
rect 10092 4870 10102 4922
rect 10102 4870 10148 4922
rect 9852 4868 9908 4870
rect 9932 4868 9988 4870
rect 10012 4868 10068 4870
rect 10092 4868 10148 4870
rect 10966 7792 11022 7848
rect 10690 5652 10692 5672
rect 10692 5652 10744 5672
rect 10744 5652 10746 5672
rect 10690 5616 10746 5652
rect 10874 6160 10930 6216
rect 11150 5652 11152 5672
rect 11152 5652 11204 5672
rect 11204 5652 11206 5672
rect 11150 5616 11206 5652
rect 10874 5072 10930 5128
rect 11334 6568 11390 6624
rect 11334 5228 11390 5264
rect 11334 5208 11336 5228
rect 11336 5208 11388 5228
rect 11388 5208 11390 5228
rect 16302 17720 16358 17776
rect 15782 16890 15838 16892
rect 15862 16890 15918 16892
rect 15942 16890 15998 16892
rect 16022 16890 16078 16892
rect 15782 16838 15828 16890
rect 15828 16838 15838 16890
rect 15862 16838 15892 16890
rect 15892 16838 15904 16890
rect 15904 16838 15918 16890
rect 15942 16838 15956 16890
rect 15956 16838 15968 16890
rect 15968 16838 15998 16890
rect 16022 16838 16032 16890
rect 16032 16838 16078 16890
rect 15782 16836 15838 16838
rect 15862 16836 15918 16838
rect 15942 16836 15998 16838
rect 16022 16836 16078 16838
rect 12817 14170 12873 14172
rect 12897 14170 12953 14172
rect 12977 14170 13033 14172
rect 13057 14170 13113 14172
rect 12817 14118 12863 14170
rect 12863 14118 12873 14170
rect 12897 14118 12927 14170
rect 12927 14118 12939 14170
rect 12939 14118 12953 14170
rect 12977 14118 12991 14170
rect 12991 14118 13003 14170
rect 13003 14118 13033 14170
rect 13057 14118 13067 14170
rect 13067 14118 13113 14170
rect 12817 14116 12873 14118
rect 12897 14116 12953 14118
rect 12977 14116 13033 14118
rect 13057 14116 13113 14118
rect 12817 13082 12873 13084
rect 12897 13082 12953 13084
rect 12977 13082 13033 13084
rect 13057 13082 13113 13084
rect 12817 13030 12863 13082
rect 12863 13030 12873 13082
rect 12897 13030 12927 13082
rect 12927 13030 12939 13082
rect 12939 13030 12953 13082
rect 12977 13030 12991 13082
rect 12991 13030 13003 13082
rect 13003 13030 13033 13082
rect 13057 13030 13067 13082
rect 13067 13030 13113 13082
rect 12817 13028 12873 13030
rect 12897 13028 12953 13030
rect 12977 13028 13033 13030
rect 13057 13028 13113 13030
rect 11886 9424 11942 9480
rect 12817 11994 12873 11996
rect 12897 11994 12953 11996
rect 12977 11994 13033 11996
rect 13057 11994 13113 11996
rect 12817 11942 12863 11994
rect 12863 11942 12873 11994
rect 12897 11942 12927 11994
rect 12927 11942 12939 11994
rect 12939 11942 12953 11994
rect 12977 11942 12991 11994
rect 12991 11942 13003 11994
rect 13003 11942 13033 11994
rect 13057 11942 13067 11994
rect 13067 11942 13113 11994
rect 12817 11940 12873 11942
rect 12897 11940 12953 11942
rect 12977 11940 13033 11942
rect 13057 11940 13113 11942
rect 12530 9596 12532 9616
rect 12532 9596 12584 9616
rect 12584 9596 12586 9616
rect 12530 9560 12586 9596
rect 12070 8336 12126 8392
rect 12622 8880 12678 8936
rect 12817 10906 12873 10908
rect 12897 10906 12953 10908
rect 12977 10906 13033 10908
rect 13057 10906 13113 10908
rect 12817 10854 12863 10906
rect 12863 10854 12873 10906
rect 12897 10854 12927 10906
rect 12927 10854 12939 10906
rect 12939 10854 12953 10906
rect 12977 10854 12991 10906
rect 12991 10854 13003 10906
rect 13003 10854 13033 10906
rect 13057 10854 13067 10906
rect 13067 10854 13113 10906
rect 12817 10852 12873 10854
rect 12897 10852 12953 10854
rect 12977 10852 13033 10854
rect 13057 10852 13113 10854
rect 14922 12844 14978 12880
rect 14922 12824 14924 12844
rect 14924 12824 14976 12844
rect 14976 12824 14978 12844
rect 12817 9818 12873 9820
rect 12897 9818 12953 9820
rect 12977 9818 13033 9820
rect 13057 9818 13113 9820
rect 12817 9766 12863 9818
rect 12863 9766 12873 9818
rect 12897 9766 12927 9818
rect 12927 9766 12939 9818
rect 12939 9766 12953 9818
rect 12977 9766 12991 9818
rect 12991 9766 13003 9818
rect 13003 9766 13033 9818
rect 13057 9766 13067 9818
rect 13067 9766 13113 9818
rect 12817 9764 12873 9766
rect 12897 9764 12953 9766
rect 12977 9764 13033 9766
rect 13057 9764 13113 9766
rect 12990 9016 13046 9072
rect 11886 7792 11942 7848
rect 9852 3834 9908 3836
rect 9932 3834 9988 3836
rect 10012 3834 10068 3836
rect 10092 3834 10148 3836
rect 9852 3782 9898 3834
rect 9898 3782 9908 3834
rect 9932 3782 9962 3834
rect 9962 3782 9974 3834
rect 9974 3782 9988 3834
rect 10012 3782 10026 3834
rect 10026 3782 10038 3834
rect 10038 3782 10068 3834
rect 10092 3782 10102 3834
rect 10102 3782 10148 3834
rect 9852 3780 9908 3782
rect 9932 3780 9988 3782
rect 10012 3780 10068 3782
rect 10092 3780 10148 3782
rect 11242 3440 11298 3496
rect 9852 2746 9908 2748
rect 9932 2746 9988 2748
rect 10012 2746 10068 2748
rect 10092 2746 10148 2748
rect 9852 2694 9898 2746
rect 9898 2694 9908 2746
rect 9932 2694 9962 2746
rect 9962 2694 9974 2746
rect 9974 2694 9988 2746
rect 10012 2694 10026 2746
rect 10026 2694 10038 2746
rect 10038 2694 10068 2746
rect 10092 2694 10102 2746
rect 10102 2694 10148 2746
rect 9852 2692 9908 2694
rect 9932 2692 9988 2694
rect 10012 2692 10068 2694
rect 10092 2692 10148 2694
rect 12817 8730 12873 8732
rect 12897 8730 12953 8732
rect 12977 8730 13033 8732
rect 13057 8730 13113 8732
rect 12817 8678 12863 8730
rect 12863 8678 12873 8730
rect 12897 8678 12927 8730
rect 12927 8678 12939 8730
rect 12939 8678 12953 8730
rect 12977 8678 12991 8730
rect 12991 8678 13003 8730
rect 13003 8678 13033 8730
rect 13057 8678 13067 8730
rect 13067 8678 13113 8730
rect 12817 8676 12873 8678
rect 12897 8676 12953 8678
rect 12977 8676 13033 8678
rect 13057 8676 13113 8678
rect 12990 8336 13046 8392
rect 12254 6840 12310 6896
rect 12817 7642 12873 7644
rect 12897 7642 12953 7644
rect 12977 7642 13033 7644
rect 13057 7642 13113 7644
rect 12817 7590 12863 7642
rect 12863 7590 12873 7642
rect 12897 7590 12927 7642
rect 12927 7590 12939 7642
rect 12939 7590 12953 7642
rect 12977 7590 12991 7642
rect 12991 7590 13003 7642
rect 13003 7590 13033 7642
rect 13057 7590 13067 7642
rect 13067 7590 13113 7642
rect 12817 7588 12873 7590
rect 12897 7588 12953 7590
rect 12977 7588 13033 7590
rect 13057 7588 13113 7590
rect 12898 6976 12954 7032
rect 12254 6432 12310 6488
rect 12530 6568 12586 6624
rect 12346 5344 12402 5400
rect 12806 6704 12862 6760
rect 12817 6554 12873 6556
rect 12897 6554 12953 6556
rect 12977 6554 13033 6556
rect 13057 6554 13113 6556
rect 12817 6502 12863 6554
rect 12863 6502 12873 6554
rect 12897 6502 12927 6554
rect 12927 6502 12939 6554
rect 12939 6502 12953 6554
rect 12977 6502 12991 6554
rect 12991 6502 13003 6554
rect 13003 6502 13033 6554
rect 13057 6502 13067 6554
rect 13067 6502 13113 6554
rect 12817 6500 12873 6502
rect 12897 6500 12953 6502
rect 12977 6500 13033 6502
rect 13057 6500 13113 6502
rect 13358 8492 13414 8528
rect 13358 8472 13360 8492
rect 13360 8472 13412 8492
rect 13412 8472 13414 8492
rect 12817 5466 12873 5468
rect 12897 5466 12953 5468
rect 12977 5466 13033 5468
rect 13057 5466 13113 5468
rect 12817 5414 12863 5466
rect 12863 5414 12873 5466
rect 12897 5414 12927 5466
rect 12927 5414 12939 5466
rect 12939 5414 12953 5466
rect 12977 5414 12991 5466
rect 12991 5414 13003 5466
rect 13003 5414 13033 5466
rect 13057 5414 13067 5466
rect 13067 5414 13113 5466
rect 12817 5412 12873 5414
rect 12897 5412 12953 5414
rect 12977 5412 13033 5414
rect 13057 5412 13113 5414
rect 12817 4378 12873 4380
rect 12897 4378 12953 4380
rect 12977 4378 13033 4380
rect 13057 4378 13113 4380
rect 12817 4326 12863 4378
rect 12863 4326 12873 4378
rect 12897 4326 12927 4378
rect 12927 4326 12939 4378
rect 12939 4326 12953 4378
rect 12977 4326 12991 4378
rect 12991 4326 13003 4378
rect 13003 4326 13033 4378
rect 13057 4326 13067 4378
rect 13067 4326 13113 4378
rect 12817 4324 12873 4326
rect 12897 4324 12953 4326
rect 12977 4324 13033 4326
rect 13057 4324 13113 4326
rect 13450 3984 13506 4040
rect 12817 3290 12873 3292
rect 12897 3290 12953 3292
rect 12977 3290 13033 3292
rect 13057 3290 13113 3292
rect 12817 3238 12863 3290
rect 12863 3238 12873 3290
rect 12897 3238 12927 3290
rect 12927 3238 12939 3290
rect 12939 3238 12953 3290
rect 12977 3238 12991 3290
rect 12991 3238 13003 3290
rect 13003 3238 13033 3290
rect 13057 3238 13067 3290
rect 13067 3238 13113 3290
rect 12817 3236 12873 3238
rect 12897 3236 12953 3238
rect 12977 3236 13033 3238
rect 13057 3236 13113 3238
rect 13818 7792 13874 7848
rect 13818 7656 13874 7712
rect 14002 8492 14058 8528
rect 14002 8472 14004 8492
rect 14004 8472 14056 8492
rect 14056 8472 14058 8492
rect 14002 8336 14058 8392
rect 14186 8472 14242 8528
rect 14278 8336 14334 8392
rect 14186 7928 14242 7984
rect 13910 6160 13966 6216
rect 13634 3052 13690 3088
rect 13634 3032 13636 3052
rect 13636 3032 13688 3052
rect 13688 3032 13690 3052
rect 14462 7656 14518 7712
rect 14646 6296 14702 6352
rect 15782 15802 15838 15804
rect 15862 15802 15918 15804
rect 15942 15802 15998 15804
rect 16022 15802 16078 15804
rect 15782 15750 15828 15802
rect 15828 15750 15838 15802
rect 15862 15750 15892 15802
rect 15892 15750 15904 15802
rect 15904 15750 15918 15802
rect 15942 15750 15956 15802
rect 15956 15750 15968 15802
rect 15968 15750 15998 15802
rect 16022 15750 16032 15802
rect 16032 15750 16078 15802
rect 15782 15748 15838 15750
rect 15862 15748 15918 15750
rect 15942 15748 15998 15750
rect 16022 15748 16078 15750
rect 15782 14714 15838 14716
rect 15862 14714 15918 14716
rect 15942 14714 15998 14716
rect 16022 14714 16078 14716
rect 15782 14662 15828 14714
rect 15828 14662 15838 14714
rect 15862 14662 15892 14714
rect 15892 14662 15904 14714
rect 15904 14662 15918 14714
rect 15942 14662 15956 14714
rect 15956 14662 15968 14714
rect 15968 14662 15998 14714
rect 16022 14662 16032 14714
rect 16032 14662 16078 14714
rect 15782 14660 15838 14662
rect 15862 14660 15918 14662
rect 15942 14660 15998 14662
rect 16022 14660 16078 14662
rect 15782 13626 15838 13628
rect 15862 13626 15918 13628
rect 15942 13626 15998 13628
rect 16022 13626 16078 13628
rect 15782 13574 15828 13626
rect 15828 13574 15838 13626
rect 15862 13574 15892 13626
rect 15892 13574 15904 13626
rect 15904 13574 15918 13626
rect 15942 13574 15956 13626
rect 15956 13574 15968 13626
rect 15968 13574 15998 13626
rect 16022 13574 16032 13626
rect 16032 13574 16078 13626
rect 15782 13572 15838 13574
rect 15862 13572 15918 13574
rect 15942 13572 15998 13574
rect 16022 13572 16078 13574
rect 15782 12538 15838 12540
rect 15862 12538 15918 12540
rect 15942 12538 15998 12540
rect 16022 12538 16078 12540
rect 15782 12486 15828 12538
rect 15828 12486 15838 12538
rect 15862 12486 15892 12538
rect 15892 12486 15904 12538
rect 15904 12486 15918 12538
rect 15942 12486 15956 12538
rect 15956 12486 15968 12538
rect 15968 12486 15998 12538
rect 16022 12486 16032 12538
rect 16032 12486 16078 12538
rect 15782 12484 15838 12486
rect 15862 12484 15918 12486
rect 15942 12484 15998 12486
rect 16022 12484 16078 12486
rect 15782 11450 15838 11452
rect 15862 11450 15918 11452
rect 15942 11450 15998 11452
rect 16022 11450 16078 11452
rect 15782 11398 15828 11450
rect 15828 11398 15838 11450
rect 15862 11398 15892 11450
rect 15892 11398 15904 11450
rect 15904 11398 15918 11450
rect 15942 11398 15956 11450
rect 15956 11398 15968 11450
rect 15968 11398 15998 11450
rect 16022 11398 16032 11450
rect 16032 11398 16078 11450
rect 15782 11396 15838 11398
rect 15862 11396 15918 11398
rect 15942 11396 15998 11398
rect 16022 11396 16078 11398
rect 15658 11076 15714 11112
rect 15658 11056 15660 11076
rect 15660 11056 15712 11076
rect 15712 11056 15714 11076
rect 14370 5480 14426 5536
rect 14186 5228 14242 5264
rect 14186 5208 14188 5228
rect 14188 5208 14240 5228
rect 14240 5208 14242 5228
rect 15782 10362 15838 10364
rect 15862 10362 15918 10364
rect 15942 10362 15998 10364
rect 16022 10362 16078 10364
rect 15782 10310 15828 10362
rect 15828 10310 15838 10362
rect 15862 10310 15892 10362
rect 15892 10310 15904 10362
rect 15904 10310 15918 10362
rect 15942 10310 15956 10362
rect 15956 10310 15968 10362
rect 15968 10310 15998 10362
rect 16022 10310 16032 10362
rect 16032 10310 16078 10362
rect 15782 10308 15838 10310
rect 15862 10308 15918 10310
rect 15942 10308 15998 10310
rect 16022 10308 16078 10310
rect 15566 9424 15622 9480
rect 15106 6976 15162 7032
rect 15014 6568 15070 6624
rect 15198 6704 15254 6760
rect 15382 6568 15438 6624
rect 15290 6160 15346 6216
rect 12817 2202 12873 2204
rect 12897 2202 12953 2204
rect 12977 2202 13033 2204
rect 13057 2202 13113 2204
rect 12817 2150 12863 2202
rect 12863 2150 12873 2202
rect 12897 2150 12927 2202
rect 12927 2150 12939 2202
rect 12939 2150 12953 2202
rect 12977 2150 12991 2202
rect 12991 2150 13003 2202
rect 13003 2150 13033 2202
rect 13057 2150 13067 2202
rect 13067 2150 13113 2202
rect 12817 2148 12873 2150
rect 12897 2148 12953 2150
rect 12977 2148 13033 2150
rect 13057 2148 13113 2150
rect 15198 3304 15254 3360
rect 15782 9274 15838 9276
rect 15862 9274 15918 9276
rect 15942 9274 15998 9276
rect 16022 9274 16078 9276
rect 15782 9222 15828 9274
rect 15828 9222 15838 9274
rect 15862 9222 15892 9274
rect 15892 9222 15904 9274
rect 15904 9222 15918 9274
rect 15942 9222 15956 9274
rect 15956 9222 15968 9274
rect 15968 9222 15998 9274
rect 16022 9222 16032 9274
rect 16032 9222 16078 9274
rect 15782 9220 15838 9222
rect 15862 9220 15918 9222
rect 15942 9220 15998 9222
rect 16022 9220 16078 9222
rect 15782 8186 15838 8188
rect 15862 8186 15918 8188
rect 15942 8186 15998 8188
rect 16022 8186 16078 8188
rect 15782 8134 15828 8186
rect 15828 8134 15838 8186
rect 15862 8134 15892 8186
rect 15892 8134 15904 8186
rect 15904 8134 15918 8186
rect 15942 8134 15956 8186
rect 15956 8134 15968 8186
rect 15968 8134 15998 8186
rect 16022 8134 16032 8186
rect 16032 8134 16078 8186
rect 15782 8132 15838 8134
rect 15862 8132 15918 8134
rect 15942 8132 15998 8134
rect 16022 8132 16078 8134
rect 17130 8472 17186 8528
rect 15782 7098 15838 7100
rect 15862 7098 15918 7100
rect 15942 7098 15998 7100
rect 16022 7098 16078 7100
rect 15782 7046 15828 7098
rect 15828 7046 15838 7098
rect 15862 7046 15892 7098
rect 15892 7046 15904 7098
rect 15904 7046 15918 7098
rect 15942 7046 15956 7098
rect 15956 7046 15968 7098
rect 15968 7046 15998 7098
rect 16022 7046 16032 7098
rect 16032 7046 16078 7098
rect 15782 7044 15838 7046
rect 15862 7044 15918 7046
rect 15942 7044 15998 7046
rect 16022 7044 16078 7046
rect 16486 7520 16542 7576
rect 16394 6704 16450 6760
rect 16302 6160 16358 6216
rect 15782 6010 15838 6012
rect 15862 6010 15918 6012
rect 15942 6010 15998 6012
rect 16022 6010 16078 6012
rect 15782 5958 15828 6010
rect 15828 5958 15838 6010
rect 15862 5958 15892 6010
rect 15892 5958 15904 6010
rect 15904 5958 15918 6010
rect 15942 5958 15956 6010
rect 15956 5958 15968 6010
rect 15968 5958 15998 6010
rect 16022 5958 16032 6010
rect 16032 5958 16078 6010
rect 15782 5956 15838 5958
rect 15862 5956 15918 5958
rect 15942 5956 15998 5958
rect 16022 5956 16078 5958
rect 15782 4922 15838 4924
rect 15862 4922 15918 4924
rect 15942 4922 15998 4924
rect 16022 4922 16078 4924
rect 15782 4870 15828 4922
rect 15828 4870 15838 4922
rect 15862 4870 15892 4922
rect 15892 4870 15904 4922
rect 15904 4870 15918 4922
rect 15942 4870 15956 4922
rect 15956 4870 15968 4922
rect 15968 4870 15998 4922
rect 16022 4870 16032 4922
rect 16032 4870 16078 4922
rect 15782 4868 15838 4870
rect 15862 4868 15918 4870
rect 15942 4868 15998 4870
rect 16022 4868 16078 4870
rect 16210 4820 16266 4856
rect 16210 4800 16212 4820
rect 16212 4800 16264 4820
rect 16264 4800 16266 4820
rect 15382 3032 15438 3088
rect 15782 3834 15838 3836
rect 15862 3834 15918 3836
rect 15942 3834 15998 3836
rect 16022 3834 16078 3836
rect 15782 3782 15828 3834
rect 15828 3782 15838 3834
rect 15862 3782 15892 3834
rect 15892 3782 15904 3834
rect 15904 3782 15918 3834
rect 15942 3782 15956 3834
rect 15956 3782 15968 3834
rect 15968 3782 15998 3834
rect 16022 3782 16032 3834
rect 16032 3782 16078 3834
rect 15782 3780 15838 3782
rect 15862 3780 15918 3782
rect 15942 3780 15998 3782
rect 16022 3780 16078 3782
rect 15782 2746 15838 2748
rect 15862 2746 15918 2748
rect 15942 2746 15998 2748
rect 16022 2746 16078 2748
rect 15782 2694 15828 2746
rect 15828 2694 15838 2746
rect 15862 2694 15892 2746
rect 15892 2694 15904 2746
rect 15904 2694 15918 2746
rect 15942 2694 15956 2746
rect 15956 2694 15968 2746
rect 15968 2694 15998 2746
rect 16022 2694 16032 2746
rect 16032 2694 16078 2746
rect 15782 2692 15838 2694
rect 15862 2692 15918 2694
rect 15942 2692 15998 2694
rect 16022 2692 16078 2694
rect 17682 17060 17738 17096
rect 17682 17040 17684 17060
rect 17684 17040 17736 17060
rect 17736 17040 17738 17060
rect 18050 15952 18106 16008
rect 18326 15680 18382 15736
rect 17866 15000 17922 15056
rect 18326 14356 18328 14376
rect 18328 14356 18380 14376
rect 18380 14356 18382 14376
rect 18326 14320 18382 14356
rect 18234 12980 18290 13016
rect 18234 12960 18236 12980
rect 18236 12960 18288 12980
rect 18288 12960 18290 12980
rect 16486 5072 16542 5128
rect 18326 11600 18382 11656
rect 17498 8916 17500 8936
rect 17500 8916 17552 8936
rect 17552 8916 17554 8936
rect 17498 8880 17554 8916
rect 17774 6840 17830 6896
rect 17958 9580 18014 9616
rect 17958 9560 17960 9580
rect 17960 9560 18012 9580
rect 18012 9560 18014 9580
rect 17958 9424 18014 9480
rect 18234 9596 18236 9616
rect 18236 9596 18288 9616
rect 18288 9596 18290 9616
rect 18234 9560 18290 9596
rect 17498 4800 17554 4856
rect 18234 4120 18290 4176
rect 17682 3984 17738 4040
rect 17038 3476 17040 3496
rect 17040 3476 17092 3496
rect 17092 3476 17094 3496
rect 17038 3440 17094 3476
rect 16118 2080 16174 2136
rect 17682 720 17738 776
<< metal3 >>
rect 0 19728 800 19848
rect 19200 19728 20000 19848
rect 0 19138 800 19168
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 19200 18368 20000 18488
rect 0 17778 800 17808
rect 2221 17778 2287 17781
rect 0 17776 2287 17778
rect 0 17720 2226 17776
rect 2282 17720 2287 17776
rect 0 17718 2287 17720
rect 0 17688 800 17718
rect 2221 17715 2287 17718
rect 16297 17778 16363 17781
rect 19200 17778 20000 17808
rect 16297 17776 20000 17778
rect 16297 17720 16302 17776
rect 16358 17720 20000 17776
rect 16297 17718 20000 17720
rect 16297 17715 16363 17718
rect 19200 17688 20000 17718
rect 6874 17440 7194 17441
rect 6874 17376 6882 17440
rect 6946 17376 6962 17440
rect 7026 17376 7042 17440
rect 7106 17376 7122 17440
rect 7186 17376 7194 17440
rect 6874 17375 7194 17376
rect 12805 17440 13125 17441
rect 12805 17376 12813 17440
rect 12877 17376 12893 17440
rect 12957 17376 12973 17440
rect 13037 17376 13053 17440
rect 13117 17376 13125 17440
rect 12805 17375 13125 17376
rect 0 17098 800 17128
rect 1393 17098 1459 17101
rect 0 17096 1459 17098
rect 0 17040 1398 17096
rect 1454 17040 1459 17096
rect 0 17038 1459 17040
rect 0 17008 800 17038
rect 1393 17035 1459 17038
rect 17677 17098 17743 17101
rect 19200 17098 20000 17128
rect 17677 17096 20000 17098
rect 17677 17040 17682 17096
rect 17738 17040 20000 17096
rect 17677 17038 20000 17040
rect 17677 17035 17743 17038
rect 19200 17008 20000 17038
rect 3909 16896 4229 16897
rect 3909 16832 3917 16896
rect 3981 16832 3997 16896
rect 4061 16832 4077 16896
rect 4141 16832 4157 16896
rect 4221 16832 4229 16896
rect 3909 16831 4229 16832
rect 9840 16896 10160 16897
rect 9840 16832 9848 16896
rect 9912 16832 9928 16896
rect 9992 16832 10008 16896
rect 10072 16832 10088 16896
rect 10152 16832 10160 16896
rect 9840 16831 10160 16832
rect 15770 16896 16090 16897
rect 15770 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15938 16896
rect 16002 16832 16018 16896
rect 16082 16832 16090 16896
rect 15770 16831 16090 16832
rect 7189 16690 7255 16693
rect 7414 16690 7420 16692
rect 7189 16688 7420 16690
rect 7189 16632 7194 16688
rect 7250 16632 7420 16688
rect 7189 16630 7420 16632
rect 7189 16627 7255 16630
rect 7414 16628 7420 16630
rect 7484 16628 7490 16692
rect 0 16328 800 16448
rect 6874 16352 7194 16353
rect 6874 16288 6882 16352
rect 6946 16288 6962 16352
rect 7026 16288 7042 16352
rect 7106 16288 7122 16352
rect 7186 16288 7194 16352
rect 6874 16287 7194 16288
rect 12805 16352 13125 16353
rect 12805 16288 12813 16352
rect 12877 16288 12893 16352
rect 12957 16288 12973 16352
rect 13037 16288 13053 16352
rect 13117 16288 13125 16352
rect 12805 16287 13125 16288
rect 10777 16146 10843 16149
rect 12617 16146 12683 16149
rect 12985 16146 13051 16149
rect 10777 16144 13051 16146
rect 10777 16088 10782 16144
rect 10838 16088 12622 16144
rect 12678 16088 12990 16144
rect 13046 16088 13051 16144
rect 10777 16086 13051 16088
rect 10777 16083 10843 16086
rect 12617 16083 12683 16086
rect 12985 16083 13051 16086
rect 7649 16010 7715 16013
rect 9213 16010 9279 16013
rect 18045 16010 18111 16013
rect 7649 16008 18111 16010
rect 7649 15952 7654 16008
rect 7710 15952 9218 16008
rect 9274 15952 18050 16008
rect 18106 15952 18111 16008
rect 7649 15950 18111 15952
rect 7649 15947 7715 15950
rect 9213 15947 9279 15950
rect 18045 15947 18111 15950
rect 3909 15808 4229 15809
rect 3909 15744 3917 15808
rect 3981 15744 3997 15808
rect 4061 15744 4077 15808
rect 4141 15744 4157 15808
rect 4221 15744 4229 15808
rect 3909 15743 4229 15744
rect 9840 15808 10160 15809
rect 9840 15744 9848 15808
rect 9912 15744 9928 15808
rect 9992 15744 10008 15808
rect 10072 15744 10088 15808
rect 10152 15744 10160 15808
rect 9840 15743 10160 15744
rect 15770 15808 16090 15809
rect 15770 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15938 15808
rect 16002 15744 16018 15808
rect 16082 15744 16090 15808
rect 15770 15743 16090 15744
rect 18321 15738 18387 15741
rect 19200 15738 20000 15768
rect 18321 15736 20000 15738
rect 18321 15680 18326 15736
rect 18382 15680 20000 15736
rect 18321 15678 20000 15680
rect 18321 15675 18387 15678
rect 19200 15648 20000 15678
rect 6874 15264 7194 15265
rect 6874 15200 6882 15264
rect 6946 15200 6962 15264
rect 7026 15200 7042 15264
rect 7106 15200 7122 15264
rect 7186 15200 7194 15264
rect 6874 15199 7194 15200
rect 12805 15264 13125 15265
rect 12805 15200 12813 15264
rect 12877 15200 12893 15264
rect 12957 15200 12973 15264
rect 13037 15200 13053 15264
rect 13117 15200 13125 15264
rect 12805 15199 13125 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 17861 15058 17927 15061
rect 19200 15058 20000 15088
rect 17861 15056 20000 15058
rect 17861 15000 17866 15056
rect 17922 15000 20000 15056
rect 17861 14998 20000 15000
rect 17861 14995 17927 14998
rect 19200 14968 20000 14998
rect 7097 14786 7163 14789
rect 8477 14786 8543 14789
rect 7097 14784 8543 14786
rect 7097 14728 7102 14784
rect 7158 14728 8482 14784
rect 8538 14728 8543 14784
rect 7097 14726 8543 14728
rect 7097 14723 7163 14726
rect 8477 14723 8543 14726
rect 3909 14720 4229 14721
rect 3909 14656 3917 14720
rect 3981 14656 3997 14720
rect 4061 14656 4077 14720
rect 4141 14656 4157 14720
rect 4221 14656 4229 14720
rect 3909 14655 4229 14656
rect 9840 14720 10160 14721
rect 9840 14656 9848 14720
rect 9912 14656 9928 14720
rect 9992 14656 10008 14720
rect 10072 14656 10088 14720
rect 10152 14656 10160 14720
rect 9840 14655 10160 14656
rect 15770 14720 16090 14721
rect 15770 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15938 14720
rect 16002 14656 16018 14720
rect 16082 14656 16090 14720
rect 15770 14655 16090 14656
rect 6729 14650 6795 14653
rect 8937 14650 9003 14653
rect 6729 14648 9003 14650
rect 6729 14592 6734 14648
rect 6790 14592 8942 14648
rect 8998 14592 9003 14648
rect 6729 14590 9003 14592
rect 6729 14587 6795 14590
rect 8937 14587 9003 14590
rect 7281 14514 7347 14517
rect 10133 14514 10199 14517
rect 7281 14512 10199 14514
rect 7281 14456 7286 14512
rect 7342 14456 10138 14512
rect 10194 14456 10199 14512
rect 7281 14454 10199 14456
rect 7281 14451 7347 14454
rect 10133 14451 10199 14454
rect 0 14378 800 14408
rect 1393 14378 1459 14381
rect 0 14376 1459 14378
rect 0 14320 1398 14376
rect 1454 14320 1459 14376
rect 0 14318 1459 14320
rect 0 14288 800 14318
rect 1393 14315 1459 14318
rect 7005 14378 7071 14381
rect 7741 14378 7807 14381
rect 7005 14376 7807 14378
rect 7005 14320 7010 14376
rect 7066 14320 7746 14376
rect 7802 14320 7807 14376
rect 7005 14318 7807 14320
rect 7005 14315 7071 14318
rect 7741 14315 7807 14318
rect 18321 14378 18387 14381
rect 19200 14378 20000 14408
rect 18321 14376 20000 14378
rect 18321 14320 18326 14376
rect 18382 14320 20000 14376
rect 18321 14318 20000 14320
rect 18321 14315 18387 14318
rect 19200 14288 20000 14318
rect 6874 14176 7194 14177
rect 6874 14112 6882 14176
rect 6946 14112 6962 14176
rect 7026 14112 7042 14176
rect 7106 14112 7122 14176
rect 7186 14112 7194 14176
rect 6874 14111 7194 14112
rect 12805 14176 13125 14177
rect 12805 14112 12813 14176
rect 12877 14112 12893 14176
rect 12957 14112 12973 14176
rect 13037 14112 13053 14176
rect 13117 14112 13125 14176
rect 12805 14111 13125 14112
rect 0 13608 800 13728
rect 3909 13632 4229 13633
rect 3909 13568 3917 13632
rect 3981 13568 3997 13632
rect 4061 13568 4077 13632
rect 4141 13568 4157 13632
rect 4221 13568 4229 13632
rect 3909 13567 4229 13568
rect 9840 13632 10160 13633
rect 9840 13568 9848 13632
rect 9912 13568 9928 13632
rect 9992 13568 10008 13632
rect 10072 13568 10088 13632
rect 10152 13568 10160 13632
rect 9840 13567 10160 13568
rect 15770 13632 16090 13633
rect 15770 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15938 13632
rect 16002 13568 16018 13632
rect 16082 13568 16090 13632
rect 15770 13567 16090 13568
rect 6874 13088 7194 13089
rect 6874 13024 6882 13088
rect 6946 13024 6962 13088
rect 7026 13024 7042 13088
rect 7106 13024 7122 13088
rect 7186 13024 7194 13088
rect 6874 13023 7194 13024
rect 12805 13088 13125 13089
rect 12805 13024 12813 13088
rect 12877 13024 12893 13088
rect 12957 13024 12973 13088
rect 13037 13024 13053 13088
rect 13117 13024 13125 13088
rect 12805 13023 13125 13024
rect 18229 13018 18295 13021
rect 19200 13018 20000 13048
rect 18229 13016 20000 13018
rect 18229 12960 18234 13016
rect 18290 12960 20000 13016
rect 18229 12958 20000 12960
rect 18229 12955 18295 12958
rect 19200 12928 20000 12958
rect 10685 12882 10751 12885
rect 14917 12882 14983 12885
rect 10685 12880 14983 12882
rect 10685 12824 10690 12880
rect 10746 12824 14922 12880
rect 14978 12824 14983 12880
rect 10685 12822 14983 12824
rect 10685 12819 10751 12822
rect 14917 12819 14983 12822
rect 3909 12544 4229 12545
rect 3909 12480 3917 12544
rect 3981 12480 3997 12544
rect 4061 12480 4077 12544
rect 4141 12480 4157 12544
rect 4221 12480 4229 12544
rect 3909 12479 4229 12480
rect 9840 12544 10160 12545
rect 9840 12480 9848 12544
rect 9912 12480 9928 12544
rect 9992 12480 10008 12544
rect 10072 12480 10088 12544
rect 10152 12480 10160 12544
rect 9840 12479 10160 12480
rect 15770 12544 16090 12545
rect 15770 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15938 12544
rect 16002 12480 16018 12544
rect 16082 12480 16090 12544
rect 15770 12479 16090 12480
rect 0 12248 800 12368
rect 19200 12248 20000 12368
rect 6874 12000 7194 12001
rect 6874 11936 6882 12000
rect 6946 11936 6962 12000
rect 7026 11936 7042 12000
rect 7106 11936 7122 12000
rect 7186 11936 7194 12000
rect 6874 11935 7194 11936
rect 12805 12000 13125 12001
rect 12805 11936 12813 12000
rect 12877 11936 12893 12000
rect 12957 11936 12973 12000
rect 13037 11936 13053 12000
rect 13117 11936 13125 12000
rect 12805 11935 13125 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 18321 11658 18387 11661
rect 19200 11658 20000 11688
rect 18321 11656 20000 11658
rect 18321 11600 18326 11656
rect 18382 11600 20000 11656
rect 18321 11598 20000 11600
rect 18321 11595 18387 11598
rect 19200 11568 20000 11598
rect 3909 11456 4229 11457
rect 3909 11392 3917 11456
rect 3981 11392 3997 11456
rect 4061 11392 4077 11456
rect 4141 11392 4157 11456
rect 4221 11392 4229 11456
rect 3909 11391 4229 11392
rect 9840 11456 10160 11457
rect 9840 11392 9848 11456
rect 9912 11392 9928 11456
rect 9992 11392 10008 11456
rect 10072 11392 10088 11456
rect 10152 11392 10160 11456
rect 9840 11391 10160 11392
rect 15770 11456 16090 11457
rect 15770 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15938 11456
rect 16002 11392 16018 11456
rect 16082 11392 16090 11456
rect 15770 11391 16090 11392
rect 15142 11052 15148 11116
rect 15212 11114 15218 11116
rect 15653 11114 15719 11117
rect 15212 11112 15719 11114
rect 15212 11056 15658 11112
rect 15714 11056 15719 11112
rect 15212 11054 15719 11056
rect 15212 11052 15218 11054
rect 15653 11051 15719 11054
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 6874 10912 7194 10913
rect 6874 10848 6882 10912
rect 6946 10848 6962 10912
rect 7026 10848 7042 10912
rect 7106 10848 7122 10912
rect 7186 10848 7194 10912
rect 6874 10847 7194 10848
rect 12805 10912 13125 10913
rect 12805 10848 12813 10912
rect 12877 10848 12893 10912
rect 12957 10848 12973 10912
rect 13037 10848 13053 10912
rect 13117 10848 13125 10912
rect 12805 10847 13125 10848
rect 3909 10368 4229 10369
rect 3909 10304 3917 10368
rect 3981 10304 3997 10368
rect 4061 10304 4077 10368
rect 4141 10304 4157 10368
rect 4221 10304 4229 10368
rect 3909 10303 4229 10304
rect 9840 10368 10160 10369
rect 9840 10304 9848 10368
rect 9912 10304 9928 10368
rect 9992 10304 10008 10368
rect 10072 10304 10088 10368
rect 10152 10304 10160 10368
rect 9840 10303 10160 10304
rect 15770 10368 16090 10369
rect 15770 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15938 10368
rect 16002 10304 16018 10368
rect 16082 10304 16090 10368
rect 15770 10303 16090 10304
rect 19200 10208 20000 10328
rect 3049 10162 3115 10165
rect 7414 10162 7420 10164
rect 3049 10160 7420 10162
rect 3049 10104 3054 10160
rect 3110 10104 7420 10160
rect 3049 10102 7420 10104
rect 3049 10099 3115 10102
rect 7414 10100 7420 10102
rect 7484 10100 7490 10164
rect 6874 9824 7194 9825
rect 6874 9760 6882 9824
rect 6946 9760 6962 9824
rect 7026 9760 7042 9824
rect 7106 9760 7122 9824
rect 7186 9760 7194 9824
rect 6874 9759 7194 9760
rect 12805 9824 13125 9825
rect 12805 9760 12813 9824
rect 12877 9760 12893 9824
rect 12957 9760 12973 9824
rect 13037 9760 13053 9824
rect 13117 9760 13125 9824
rect 12805 9759 13125 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 12525 9618 12591 9621
rect 17953 9618 18019 9621
rect 12525 9616 18019 9618
rect 12525 9560 12530 9616
rect 12586 9560 17958 9616
rect 18014 9560 18019 9616
rect 12525 9558 18019 9560
rect 12525 9555 12591 9558
rect 17953 9555 18019 9558
rect 18229 9618 18295 9621
rect 19200 9618 20000 9648
rect 18229 9616 20000 9618
rect 18229 9560 18234 9616
rect 18290 9560 20000 9616
rect 18229 9558 20000 9560
rect 18229 9555 18295 9558
rect 19200 9528 20000 9558
rect 11881 9482 11947 9485
rect 15561 9482 15627 9485
rect 17953 9482 18019 9485
rect 11881 9480 18019 9482
rect 11881 9424 11886 9480
rect 11942 9424 15566 9480
rect 15622 9424 17958 9480
rect 18014 9424 18019 9480
rect 11881 9422 18019 9424
rect 11881 9419 11947 9422
rect 15561 9419 15627 9422
rect 17953 9419 18019 9422
rect 3909 9280 4229 9281
rect 3909 9216 3917 9280
rect 3981 9216 3997 9280
rect 4061 9216 4077 9280
rect 4141 9216 4157 9280
rect 4221 9216 4229 9280
rect 3909 9215 4229 9216
rect 9840 9280 10160 9281
rect 9840 9216 9848 9280
rect 9912 9216 9928 9280
rect 9992 9216 10008 9280
rect 10072 9216 10088 9280
rect 10152 9216 10160 9280
rect 9840 9215 10160 9216
rect 15770 9280 16090 9281
rect 15770 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15938 9280
rect 16002 9216 16018 9280
rect 16082 9216 16090 9280
rect 15770 9215 16090 9216
rect 10869 9074 10935 9077
rect 12985 9074 13051 9077
rect 10869 9072 13051 9074
rect 10869 9016 10874 9072
rect 10930 9016 12990 9072
rect 13046 9016 13051 9072
rect 10869 9014 13051 9016
rect 10869 9011 10935 9014
rect 12985 9011 13051 9014
rect 0 8938 800 8968
rect 1485 8938 1551 8941
rect 0 8936 1551 8938
rect 0 8880 1490 8936
rect 1546 8880 1551 8936
rect 0 8878 1551 8880
rect 0 8848 800 8878
rect 1485 8875 1551 8878
rect 4429 8938 4495 8941
rect 12617 8938 12683 8941
rect 4429 8936 12683 8938
rect 4429 8880 4434 8936
rect 4490 8880 12622 8936
rect 12678 8880 12683 8936
rect 4429 8878 12683 8880
rect 4429 8875 4495 8878
rect 12617 8875 12683 8878
rect 17493 8938 17559 8941
rect 19200 8938 20000 8968
rect 17493 8936 20000 8938
rect 17493 8880 17498 8936
rect 17554 8880 20000 8936
rect 17493 8878 20000 8880
rect 17493 8875 17559 8878
rect 19200 8848 20000 8878
rect 6874 8736 7194 8737
rect 6874 8672 6882 8736
rect 6946 8672 6962 8736
rect 7026 8672 7042 8736
rect 7106 8672 7122 8736
rect 7186 8672 7194 8736
rect 6874 8671 7194 8672
rect 12805 8736 13125 8737
rect 12805 8672 12813 8736
rect 12877 8672 12893 8736
rect 12957 8672 12973 8736
rect 13037 8672 13053 8736
rect 13117 8672 13125 8736
rect 12805 8671 13125 8672
rect 5165 8530 5231 8533
rect 13353 8530 13419 8533
rect 13997 8532 14063 8533
rect 13997 8530 14044 8532
rect 5165 8528 13419 8530
rect 5165 8472 5170 8528
rect 5226 8472 13358 8528
rect 13414 8472 13419 8528
rect 5165 8470 13419 8472
rect 13952 8528 14044 8530
rect 13952 8472 14002 8528
rect 13952 8470 14044 8472
rect 5165 8467 5231 8470
rect 13353 8467 13419 8470
rect 13997 8468 14044 8470
rect 14108 8468 14114 8532
rect 14181 8530 14247 8533
rect 17125 8530 17191 8533
rect 14181 8528 17191 8530
rect 14181 8472 14186 8528
rect 14242 8472 17130 8528
rect 17186 8472 17191 8528
rect 14181 8470 17191 8472
rect 13997 8467 14063 8468
rect 14181 8467 14247 8470
rect 17125 8467 17191 8470
rect 12065 8394 12131 8397
rect 12985 8394 13051 8397
rect 13997 8394 14063 8397
rect 14273 8394 14339 8397
rect 12065 8392 14339 8394
rect 12065 8336 12070 8392
rect 12126 8336 12990 8392
rect 13046 8336 14002 8392
rect 14058 8336 14278 8392
rect 14334 8336 14339 8392
rect 12065 8334 14339 8336
rect 12065 8331 12131 8334
rect 12985 8331 13051 8334
rect 13997 8331 14063 8334
rect 14273 8331 14339 8334
rect 0 8168 800 8288
rect 3909 8192 4229 8193
rect 3909 8128 3917 8192
rect 3981 8128 3997 8192
rect 4061 8128 4077 8192
rect 4141 8128 4157 8192
rect 4221 8128 4229 8192
rect 3909 8127 4229 8128
rect 9840 8192 10160 8193
rect 9840 8128 9848 8192
rect 9912 8128 9928 8192
rect 9992 8128 10008 8192
rect 10072 8128 10088 8192
rect 10152 8128 10160 8192
rect 9840 8127 10160 8128
rect 15770 8192 16090 8193
rect 15770 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15938 8192
rect 16002 8128 16018 8192
rect 16082 8128 16090 8192
rect 15770 8127 16090 8128
rect 7833 7986 7899 7989
rect 14181 7986 14247 7989
rect 7833 7984 14247 7986
rect 7833 7928 7838 7984
rect 7894 7928 14186 7984
rect 14242 7928 14247 7984
rect 7833 7926 14247 7928
rect 7833 7923 7899 7926
rect 14181 7923 14247 7926
rect 10961 7850 11027 7853
rect 10918 7848 11027 7850
rect 10918 7792 10966 7848
rect 11022 7792 11027 7848
rect 10918 7787 11027 7792
rect 11881 7850 11947 7853
rect 13813 7850 13879 7853
rect 11881 7848 13879 7850
rect 11881 7792 11886 7848
rect 11942 7792 13818 7848
rect 13874 7792 13879 7848
rect 11881 7790 13879 7792
rect 11881 7787 11947 7790
rect 13813 7787 13879 7790
rect 10685 7714 10751 7717
rect 10918 7714 10978 7787
rect 10685 7712 10978 7714
rect 10685 7656 10690 7712
rect 10746 7656 10978 7712
rect 10685 7654 10978 7656
rect 13813 7714 13879 7717
rect 14457 7714 14523 7717
rect 13813 7712 14523 7714
rect 13813 7656 13818 7712
rect 13874 7656 14462 7712
rect 14518 7656 14523 7712
rect 13813 7654 14523 7656
rect 10685 7651 10751 7654
rect 13813 7651 13879 7654
rect 14457 7651 14523 7654
rect 6874 7648 7194 7649
rect 6874 7584 6882 7648
rect 6946 7584 6962 7648
rect 7026 7584 7042 7648
rect 7106 7584 7122 7648
rect 7186 7584 7194 7648
rect 6874 7583 7194 7584
rect 12805 7648 13125 7649
rect 12805 7584 12813 7648
rect 12877 7584 12893 7648
rect 12957 7584 12973 7648
rect 13037 7584 13053 7648
rect 13117 7584 13125 7648
rect 12805 7583 13125 7584
rect 16481 7578 16547 7581
rect 19200 7578 20000 7608
rect 16481 7576 20000 7578
rect 16481 7520 16486 7576
rect 16542 7520 20000 7576
rect 16481 7518 20000 7520
rect 16481 7515 16547 7518
rect 19200 7488 20000 7518
rect 3909 7104 4229 7105
rect 3909 7040 3917 7104
rect 3981 7040 3997 7104
rect 4061 7040 4077 7104
rect 4141 7040 4157 7104
rect 4221 7040 4229 7104
rect 3909 7039 4229 7040
rect 9840 7104 10160 7105
rect 9840 7040 9848 7104
rect 9912 7040 9928 7104
rect 9992 7040 10008 7104
rect 10072 7040 10088 7104
rect 10152 7040 10160 7104
rect 9840 7039 10160 7040
rect 15770 7104 16090 7105
rect 15770 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15938 7104
rect 16002 7040 16018 7104
rect 16082 7040 16090 7104
rect 15770 7039 16090 7040
rect 12382 6972 12388 7036
rect 12452 7034 12458 7036
rect 12893 7034 12959 7037
rect 15101 7034 15167 7037
rect 12452 7032 15167 7034
rect 12452 6976 12898 7032
rect 12954 6976 15106 7032
rect 15162 6976 15167 7032
rect 12452 6974 15167 6976
rect 12452 6972 12458 6974
rect 12893 6971 12959 6974
rect 15101 6971 15167 6974
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 2497 6898 2563 6901
rect 12249 6898 12315 6901
rect 17769 6898 17835 6901
rect 19200 6898 20000 6928
rect 2497 6896 12315 6898
rect 2497 6840 2502 6896
rect 2558 6840 12254 6896
rect 12310 6840 12315 6896
rect 2497 6838 12315 6840
rect 2497 6835 2563 6838
rect 12249 6835 12315 6838
rect 12574 6896 17835 6898
rect 12574 6840 17774 6896
rect 17830 6840 17835 6896
rect 12574 6838 17835 6840
rect 8109 6762 8175 6765
rect 12574 6762 12634 6838
rect 17769 6835 17835 6838
rect 17910 6838 20000 6898
rect 8109 6760 12634 6762
rect 8109 6704 8114 6760
rect 8170 6704 12634 6760
rect 8109 6702 12634 6704
rect 12801 6762 12867 6765
rect 15193 6762 15259 6765
rect 12801 6760 15259 6762
rect 12801 6704 12806 6760
rect 12862 6704 15198 6760
rect 15254 6704 15259 6760
rect 12801 6702 15259 6704
rect 8109 6699 8175 6702
rect 12801 6699 12867 6702
rect 15193 6699 15259 6702
rect 16389 6762 16455 6765
rect 17910 6762 17970 6838
rect 19200 6808 20000 6838
rect 16389 6760 17970 6762
rect 16389 6704 16394 6760
rect 16450 6704 17970 6760
rect 16389 6702 17970 6704
rect 16389 6699 16455 6702
rect 10501 6626 10567 6629
rect 11329 6626 11395 6629
rect 12525 6626 12591 6629
rect 10501 6624 12591 6626
rect 10501 6568 10506 6624
rect 10562 6568 11334 6624
rect 11390 6568 12530 6624
rect 12586 6568 12591 6624
rect 10501 6566 12591 6568
rect 10501 6563 10567 6566
rect 11329 6563 11395 6566
rect 12525 6563 12591 6566
rect 15009 6626 15075 6629
rect 15142 6626 15148 6628
rect 15009 6624 15148 6626
rect 15009 6568 15014 6624
rect 15070 6568 15148 6624
rect 15009 6566 15148 6568
rect 15009 6563 15075 6566
rect 15142 6564 15148 6566
rect 15212 6626 15218 6628
rect 15377 6626 15443 6629
rect 15212 6624 15443 6626
rect 15212 6568 15382 6624
rect 15438 6568 15443 6624
rect 15212 6566 15443 6568
rect 15212 6564 15218 6566
rect 15377 6563 15443 6566
rect 6874 6560 7194 6561
rect 6874 6496 6882 6560
rect 6946 6496 6962 6560
rect 7026 6496 7042 6560
rect 7106 6496 7122 6560
rect 7186 6496 7194 6560
rect 6874 6495 7194 6496
rect 12805 6560 13125 6561
rect 12805 6496 12813 6560
rect 12877 6496 12893 6560
rect 12957 6496 12973 6560
rect 13037 6496 13053 6560
rect 13117 6496 13125 6560
rect 12805 6495 13125 6496
rect 12249 6490 12315 6493
rect 12382 6490 12388 6492
rect 12249 6488 12388 6490
rect 12249 6432 12254 6488
rect 12310 6432 12388 6488
rect 12249 6430 12388 6432
rect 12249 6427 12315 6430
rect 12382 6428 12388 6430
rect 12452 6428 12458 6492
rect 5165 6354 5231 6357
rect 14641 6354 14707 6357
rect 5165 6352 14707 6354
rect 5165 6296 5170 6352
rect 5226 6296 14646 6352
rect 14702 6296 14707 6352
rect 5165 6294 14707 6296
rect 5165 6291 5231 6294
rect 14641 6291 14707 6294
rect 0 6218 800 6248
rect 1393 6218 1459 6221
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 800 6158
rect 1393 6155 1459 6158
rect 10869 6218 10935 6221
rect 13905 6218 13971 6221
rect 15285 6218 15351 6221
rect 10869 6216 15351 6218
rect 10869 6160 10874 6216
rect 10930 6160 13910 6216
rect 13966 6160 15290 6216
rect 15346 6160 15351 6216
rect 10869 6158 15351 6160
rect 10869 6155 10935 6158
rect 13905 6155 13971 6158
rect 15285 6155 15351 6158
rect 16297 6218 16363 6221
rect 19200 6218 20000 6248
rect 16297 6216 20000 6218
rect 16297 6160 16302 6216
rect 16358 6160 20000 6216
rect 16297 6158 20000 6160
rect 16297 6155 16363 6158
rect 19200 6128 20000 6158
rect 3909 6016 4229 6017
rect 3909 5952 3917 6016
rect 3981 5952 3997 6016
rect 4061 5952 4077 6016
rect 4141 5952 4157 6016
rect 4221 5952 4229 6016
rect 3909 5951 4229 5952
rect 9840 6016 10160 6017
rect 9840 5952 9848 6016
rect 9912 5952 9928 6016
rect 9992 5952 10008 6016
rect 10072 5952 10088 6016
rect 10152 5952 10160 6016
rect 9840 5951 10160 5952
rect 15770 6016 16090 6017
rect 15770 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15938 6016
rect 16002 5952 16018 6016
rect 16082 5952 16090 6016
rect 15770 5951 16090 5952
rect 10685 5674 10751 5677
rect 11145 5674 11211 5677
rect 10685 5672 11211 5674
rect 10685 5616 10690 5672
rect 10746 5616 11150 5672
rect 11206 5616 11211 5672
rect 10685 5614 11211 5616
rect 10685 5611 10751 5614
rect 11145 5611 11211 5614
rect 0 5448 800 5568
rect 14038 5476 14044 5540
rect 14108 5538 14114 5540
rect 14365 5538 14431 5541
rect 14108 5536 14431 5538
rect 14108 5480 14370 5536
rect 14426 5480 14431 5536
rect 14108 5478 14431 5480
rect 14108 5476 14114 5478
rect 14365 5475 14431 5478
rect 6874 5472 7194 5473
rect 6874 5408 6882 5472
rect 6946 5408 6962 5472
rect 7026 5408 7042 5472
rect 7106 5408 7122 5472
rect 7186 5408 7194 5472
rect 6874 5407 7194 5408
rect 12805 5472 13125 5473
rect 12805 5408 12813 5472
rect 12877 5408 12893 5472
rect 12957 5408 12973 5472
rect 13037 5408 13053 5472
rect 13117 5408 13125 5472
rect 12805 5407 13125 5408
rect 10501 5402 10567 5405
rect 12341 5402 12407 5405
rect 10501 5400 12407 5402
rect 10501 5344 10506 5400
rect 10562 5344 12346 5400
rect 12402 5344 12407 5400
rect 10501 5342 12407 5344
rect 10501 5339 10567 5342
rect 12341 5339 12407 5342
rect 11329 5266 11395 5269
rect 14181 5266 14247 5269
rect 11329 5264 14247 5266
rect 11329 5208 11334 5264
rect 11390 5208 14186 5264
rect 14242 5208 14247 5264
rect 11329 5206 14247 5208
rect 11329 5203 11395 5206
rect 14181 5203 14247 5206
rect 9949 5130 10015 5133
rect 10869 5130 10935 5133
rect 16481 5130 16547 5133
rect 9949 5128 16547 5130
rect 9949 5072 9954 5128
rect 10010 5072 10874 5128
rect 10930 5072 16486 5128
rect 16542 5072 16547 5128
rect 9949 5070 16547 5072
rect 9949 5067 10015 5070
rect 10869 5067 10935 5070
rect 16481 5067 16547 5070
rect 3909 4928 4229 4929
rect 3909 4864 3917 4928
rect 3981 4864 3997 4928
rect 4061 4864 4077 4928
rect 4141 4864 4157 4928
rect 4221 4864 4229 4928
rect 3909 4863 4229 4864
rect 9840 4928 10160 4929
rect 9840 4864 9848 4928
rect 9912 4864 9928 4928
rect 9992 4864 10008 4928
rect 10072 4864 10088 4928
rect 10152 4864 10160 4928
rect 9840 4863 10160 4864
rect 15770 4928 16090 4929
rect 15770 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15938 4928
rect 16002 4864 16018 4928
rect 16082 4864 16090 4928
rect 15770 4863 16090 4864
rect 16205 4858 16271 4861
rect 17493 4858 17559 4861
rect 19200 4858 20000 4888
rect 16205 4856 20000 4858
rect 16205 4800 16210 4856
rect 16266 4800 17498 4856
rect 17554 4800 20000 4856
rect 16205 4798 20000 4800
rect 16205 4795 16271 4798
rect 17493 4795 17559 4798
rect 19200 4768 20000 4798
rect 6874 4384 7194 4385
rect 6874 4320 6882 4384
rect 6946 4320 6962 4384
rect 7026 4320 7042 4384
rect 7106 4320 7122 4384
rect 7186 4320 7194 4384
rect 6874 4319 7194 4320
rect 12805 4384 13125 4385
rect 12805 4320 12813 4384
rect 12877 4320 12893 4384
rect 12957 4320 12973 4384
rect 13037 4320 13053 4384
rect 13117 4320 13125 4384
rect 12805 4319 13125 4320
rect 0 4088 800 4208
rect 18229 4178 18295 4181
rect 19200 4178 20000 4208
rect 18229 4176 20000 4178
rect 18229 4120 18234 4176
rect 18290 4120 20000 4176
rect 18229 4118 20000 4120
rect 18229 4115 18295 4118
rect 19200 4088 20000 4118
rect 13445 4042 13511 4045
rect 17677 4042 17743 4045
rect 13445 4040 17743 4042
rect 13445 3984 13450 4040
rect 13506 3984 17682 4040
rect 17738 3984 17743 4040
rect 13445 3982 17743 3984
rect 13445 3979 13511 3982
rect 17677 3979 17743 3982
rect 3909 3840 4229 3841
rect 3909 3776 3917 3840
rect 3981 3776 3997 3840
rect 4061 3776 4077 3840
rect 4141 3776 4157 3840
rect 4221 3776 4229 3840
rect 3909 3775 4229 3776
rect 9840 3840 10160 3841
rect 9840 3776 9848 3840
rect 9912 3776 9928 3840
rect 9992 3776 10008 3840
rect 10072 3776 10088 3840
rect 10152 3776 10160 3840
rect 9840 3775 10160 3776
rect 15770 3840 16090 3841
rect 15770 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15938 3840
rect 16002 3776 16018 3840
rect 16082 3776 16090 3840
rect 15770 3775 16090 3776
rect 0 3408 800 3528
rect 11237 3498 11303 3501
rect 17033 3498 17099 3501
rect 19200 3498 20000 3528
rect 11237 3496 17099 3498
rect 11237 3440 11242 3496
rect 11298 3440 17038 3496
rect 17094 3440 17099 3496
rect 11237 3438 17099 3440
rect 11237 3435 11303 3438
rect 17033 3435 17099 3438
rect 17174 3438 20000 3498
rect 15193 3362 15259 3365
rect 17174 3362 17234 3438
rect 19200 3408 20000 3438
rect 15193 3360 17234 3362
rect 15193 3304 15198 3360
rect 15254 3304 17234 3360
rect 15193 3302 17234 3304
rect 15193 3299 15259 3302
rect 6874 3296 7194 3297
rect 6874 3232 6882 3296
rect 6946 3232 6962 3296
rect 7026 3232 7042 3296
rect 7106 3232 7122 3296
rect 7186 3232 7194 3296
rect 6874 3231 7194 3232
rect 12805 3296 13125 3297
rect 12805 3232 12813 3296
rect 12877 3232 12893 3296
rect 12957 3232 12973 3296
rect 13037 3232 13053 3296
rect 13117 3232 13125 3296
rect 12805 3231 13125 3232
rect 13629 3090 13695 3093
rect 15377 3090 15443 3093
rect 13629 3088 15443 3090
rect 13629 3032 13634 3088
rect 13690 3032 15382 3088
rect 15438 3032 15443 3088
rect 13629 3030 15443 3032
rect 13629 3027 13695 3030
rect 15377 3027 15443 3030
rect 0 2818 800 2848
rect 2221 2818 2287 2821
rect 0 2816 2287 2818
rect 0 2760 2226 2816
rect 2282 2760 2287 2816
rect 0 2758 2287 2760
rect 0 2728 800 2758
rect 2221 2755 2287 2758
rect 3909 2752 4229 2753
rect 3909 2688 3917 2752
rect 3981 2688 3997 2752
rect 4061 2688 4077 2752
rect 4141 2688 4157 2752
rect 4221 2688 4229 2752
rect 3909 2687 4229 2688
rect 9840 2752 10160 2753
rect 9840 2688 9848 2752
rect 9912 2688 9928 2752
rect 9992 2688 10008 2752
rect 10072 2688 10088 2752
rect 10152 2688 10160 2752
rect 9840 2687 10160 2688
rect 15770 2752 16090 2753
rect 15770 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15938 2752
rect 16002 2688 16018 2752
rect 16082 2688 16090 2752
rect 15770 2687 16090 2688
rect 6874 2208 7194 2209
rect 6874 2144 6882 2208
rect 6946 2144 6962 2208
rect 7026 2144 7042 2208
rect 7106 2144 7122 2208
rect 7186 2144 7194 2208
rect 6874 2143 7194 2144
rect 12805 2208 13125 2209
rect 12805 2144 12813 2208
rect 12877 2144 12893 2208
rect 12957 2144 12973 2208
rect 13037 2144 13053 2208
rect 13117 2144 13125 2208
rect 12805 2143 13125 2144
rect 16113 2138 16179 2141
rect 19200 2138 20000 2168
rect 16113 2136 20000 2138
rect 16113 2080 16118 2136
rect 16174 2080 20000 2136
rect 16113 2078 20000 2080
rect 16113 2075 16179 2078
rect 19200 2048 20000 2078
rect 0 1458 800 1488
rect 3417 1458 3483 1461
rect 0 1456 3483 1458
rect 0 1400 3422 1456
rect 3478 1400 3483 1456
rect 0 1398 3483 1400
rect 0 1368 800 1398
rect 3417 1395 3483 1398
rect 19200 1368 20000 1488
rect 0 778 800 808
rect 2773 778 2839 781
rect 0 776 2839 778
rect 0 720 2778 776
rect 2834 720 2839 776
rect 0 718 2839 720
rect 0 688 800 718
rect 2773 715 2839 718
rect 17677 778 17743 781
rect 19200 778 20000 808
rect 17677 776 20000 778
rect 17677 720 17682 776
rect 17738 720 20000 776
rect 17677 718 20000 720
rect 17677 715 17743 718
rect 19200 688 20000 718
<< via3 >>
rect 6882 17436 6946 17440
rect 6882 17380 6886 17436
rect 6886 17380 6942 17436
rect 6942 17380 6946 17436
rect 6882 17376 6946 17380
rect 6962 17436 7026 17440
rect 6962 17380 6966 17436
rect 6966 17380 7022 17436
rect 7022 17380 7026 17436
rect 6962 17376 7026 17380
rect 7042 17436 7106 17440
rect 7042 17380 7046 17436
rect 7046 17380 7102 17436
rect 7102 17380 7106 17436
rect 7042 17376 7106 17380
rect 7122 17436 7186 17440
rect 7122 17380 7126 17436
rect 7126 17380 7182 17436
rect 7182 17380 7186 17436
rect 7122 17376 7186 17380
rect 12813 17436 12877 17440
rect 12813 17380 12817 17436
rect 12817 17380 12873 17436
rect 12873 17380 12877 17436
rect 12813 17376 12877 17380
rect 12893 17436 12957 17440
rect 12893 17380 12897 17436
rect 12897 17380 12953 17436
rect 12953 17380 12957 17436
rect 12893 17376 12957 17380
rect 12973 17436 13037 17440
rect 12973 17380 12977 17436
rect 12977 17380 13033 17436
rect 13033 17380 13037 17436
rect 12973 17376 13037 17380
rect 13053 17436 13117 17440
rect 13053 17380 13057 17436
rect 13057 17380 13113 17436
rect 13113 17380 13117 17436
rect 13053 17376 13117 17380
rect 3917 16892 3981 16896
rect 3917 16836 3921 16892
rect 3921 16836 3977 16892
rect 3977 16836 3981 16892
rect 3917 16832 3981 16836
rect 3997 16892 4061 16896
rect 3997 16836 4001 16892
rect 4001 16836 4057 16892
rect 4057 16836 4061 16892
rect 3997 16832 4061 16836
rect 4077 16892 4141 16896
rect 4077 16836 4081 16892
rect 4081 16836 4137 16892
rect 4137 16836 4141 16892
rect 4077 16832 4141 16836
rect 4157 16892 4221 16896
rect 4157 16836 4161 16892
rect 4161 16836 4217 16892
rect 4217 16836 4221 16892
rect 4157 16832 4221 16836
rect 9848 16892 9912 16896
rect 9848 16836 9852 16892
rect 9852 16836 9908 16892
rect 9908 16836 9912 16892
rect 9848 16832 9912 16836
rect 9928 16892 9992 16896
rect 9928 16836 9932 16892
rect 9932 16836 9988 16892
rect 9988 16836 9992 16892
rect 9928 16832 9992 16836
rect 10008 16892 10072 16896
rect 10008 16836 10012 16892
rect 10012 16836 10068 16892
rect 10068 16836 10072 16892
rect 10008 16832 10072 16836
rect 10088 16892 10152 16896
rect 10088 16836 10092 16892
rect 10092 16836 10148 16892
rect 10148 16836 10152 16892
rect 10088 16832 10152 16836
rect 15778 16892 15842 16896
rect 15778 16836 15782 16892
rect 15782 16836 15838 16892
rect 15838 16836 15842 16892
rect 15778 16832 15842 16836
rect 15858 16892 15922 16896
rect 15858 16836 15862 16892
rect 15862 16836 15918 16892
rect 15918 16836 15922 16892
rect 15858 16832 15922 16836
rect 15938 16892 16002 16896
rect 15938 16836 15942 16892
rect 15942 16836 15998 16892
rect 15998 16836 16002 16892
rect 15938 16832 16002 16836
rect 16018 16892 16082 16896
rect 16018 16836 16022 16892
rect 16022 16836 16078 16892
rect 16078 16836 16082 16892
rect 16018 16832 16082 16836
rect 7420 16628 7484 16692
rect 6882 16348 6946 16352
rect 6882 16292 6886 16348
rect 6886 16292 6942 16348
rect 6942 16292 6946 16348
rect 6882 16288 6946 16292
rect 6962 16348 7026 16352
rect 6962 16292 6966 16348
rect 6966 16292 7022 16348
rect 7022 16292 7026 16348
rect 6962 16288 7026 16292
rect 7042 16348 7106 16352
rect 7042 16292 7046 16348
rect 7046 16292 7102 16348
rect 7102 16292 7106 16348
rect 7042 16288 7106 16292
rect 7122 16348 7186 16352
rect 7122 16292 7126 16348
rect 7126 16292 7182 16348
rect 7182 16292 7186 16348
rect 7122 16288 7186 16292
rect 12813 16348 12877 16352
rect 12813 16292 12817 16348
rect 12817 16292 12873 16348
rect 12873 16292 12877 16348
rect 12813 16288 12877 16292
rect 12893 16348 12957 16352
rect 12893 16292 12897 16348
rect 12897 16292 12953 16348
rect 12953 16292 12957 16348
rect 12893 16288 12957 16292
rect 12973 16348 13037 16352
rect 12973 16292 12977 16348
rect 12977 16292 13033 16348
rect 13033 16292 13037 16348
rect 12973 16288 13037 16292
rect 13053 16348 13117 16352
rect 13053 16292 13057 16348
rect 13057 16292 13113 16348
rect 13113 16292 13117 16348
rect 13053 16288 13117 16292
rect 3917 15804 3981 15808
rect 3917 15748 3921 15804
rect 3921 15748 3977 15804
rect 3977 15748 3981 15804
rect 3917 15744 3981 15748
rect 3997 15804 4061 15808
rect 3997 15748 4001 15804
rect 4001 15748 4057 15804
rect 4057 15748 4061 15804
rect 3997 15744 4061 15748
rect 4077 15804 4141 15808
rect 4077 15748 4081 15804
rect 4081 15748 4137 15804
rect 4137 15748 4141 15804
rect 4077 15744 4141 15748
rect 4157 15804 4221 15808
rect 4157 15748 4161 15804
rect 4161 15748 4217 15804
rect 4217 15748 4221 15804
rect 4157 15744 4221 15748
rect 9848 15804 9912 15808
rect 9848 15748 9852 15804
rect 9852 15748 9908 15804
rect 9908 15748 9912 15804
rect 9848 15744 9912 15748
rect 9928 15804 9992 15808
rect 9928 15748 9932 15804
rect 9932 15748 9988 15804
rect 9988 15748 9992 15804
rect 9928 15744 9992 15748
rect 10008 15804 10072 15808
rect 10008 15748 10012 15804
rect 10012 15748 10068 15804
rect 10068 15748 10072 15804
rect 10008 15744 10072 15748
rect 10088 15804 10152 15808
rect 10088 15748 10092 15804
rect 10092 15748 10148 15804
rect 10148 15748 10152 15804
rect 10088 15744 10152 15748
rect 15778 15804 15842 15808
rect 15778 15748 15782 15804
rect 15782 15748 15838 15804
rect 15838 15748 15842 15804
rect 15778 15744 15842 15748
rect 15858 15804 15922 15808
rect 15858 15748 15862 15804
rect 15862 15748 15918 15804
rect 15918 15748 15922 15804
rect 15858 15744 15922 15748
rect 15938 15804 16002 15808
rect 15938 15748 15942 15804
rect 15942 15748 15998 15804
rect 15998 15748 16002 15804
rect 15938 15744 16002 15748
rect 16018 15804 16082 15808
rect 16018 15748 16022 15804
rect 16022 15748 16078 15804
rect 16078 15748 16082 15804
rect 16018 15744 16082 15748
rect 6882 15260 6946 15264
rect 6882 15204 6886 15260
rect 6886 15204 6942 15260
rect 6942 15204 6946 15260
rect 6882 15200 6946 15204
rect 6962 15260 7026 15264
rect 6962 15204 6966 15260
rect 6966 15204 7022 15260
rect 7022 15204 7026 15260
rect 6962 15200 7026 15204
rect 7042 15260 7106 15264
rect 7042 15204 7046 15260
rect 7046 15204 7102 15260
rect 7102 15204 7106 15260
rect 7042 15200 7106 15204
rect 7122 15260 7186 15264
rect 7122 15204 7126 15260
rect 7126 15204 7182 15260
rect 7182 15204 7186 15260
rect 7122 15200 7186 15204
rect 12813 15260 12877 15264
rect 12813 15204 12817 15260
rect 12817 15204 12873 15260
rect 12873 15204 12877 15260
rect 12813 15200 12877 15204
rect 12893 15260 12957 15264
rect 12893 15204 12897 15260
rect 12897 15204 12953 15260
rect 12953 15204 12957 15260
rect 12893 15200 12957 15204
rect 12973 15260 13037 15264
rect 12973 15204 12977 15260
rect 12977 15204 13033 15260
rect 13033 15204 13037 15260
rect 12973 15200 13037 15204
rect 13053 15260 13117 15264
rect 13053 15204 13057 15260
rect 13057 15204 13113 15260
rect 13113 15204 13117 15260
rect 13053 15200 13117 15204
rect 3917 14716 3981 14720
rect 3917 14660 3921 14716
rect 3921 14660 3977 14716
rect 3977 14660 3981 14716
rect 3917 14656 3981 14660
rect 3997 14716 4061 14720
rect 3997 14660 4001 14716
rect 4001 14660 4057 14716
rect 4057 14660 4061 14716
rect 3997 14656 4061 14660
rect 4077 14716 4141 14720
rect 4077 14660 4081 14716
rect 4081 14660 4137 14716
rect 4137 14660 4141 14716
rect 4077 14656 4141 14660
rect 4157 14716 4221 14720
rect 4157 14660 4161 14716
rect 4161 14660 4217 14716
rect 4217 14660 4221 14716
rect 4157 14656 4221 14660
rect 9848 14716 9912 14720
rect 9848 14660 9852 14716
rect 9852 14660 9908 14716
rect 9908 14660 9912 14716
rect 9848 14656 9912 14660
rect 9928 14716 9992 14720
rect 9928 14660 9932 14716
rect 9932 14660 9988 14716
rect 9988 14660 9992 14716
rect 9928 14656 9992 14660
rect 10008 14716 10072 14720
rect 10008 14660 10012 14716
rect 10012 14660 10068 14716
rect 10068 14660 10072 14716
rect 10008 14656 10072 14660
rect 10088 14716 10152 14720
rect 10088 14660 10092 14716
rect 10092 14660 10148 14716
rect 10148 14660 10152 14716
rect 10088 14656 10152 14660
rect 15778 14716 15842 14720
rect 15778 14660 15782 14716
rect 15782 14660 15838 14716
rect 15838 14660 15842 14716
rect 15778 14656 15842 14660
rect 15858 14716 15922 14720
rect 15858 14660 15862 14716
rect 15862 14660 15918 14716
rect 15918 14660 15922 14716
rect 15858 14656 15922 14660
rect 15938 14716 16002 14720
rect 15938 14660 15942 14716
rect 15942 14660 15998 14716
rect 15998 14660 16002 14716
rect 15938 14656 16002 14660
rect 16018 14716 16082 14720
rect 16018 14660 16022 14716
rect 16022 14660 16078 14716
rect 16078 14660 16082 14716
rect 16018 14656 16082 14660
rect 6882 14172 6946 14176
rect 6882 14116 6886 14172
rect 6886 14116 6942 14172
rect 6942 14116 6946 14172
rect 6882 14112 6946 14116
rect 6962 14172 7026 14176
rect 6962 14116 6966 14172
rect 6966 14116 7022 14172
rect 7022 14116 7026 14172
rect 6962 14112 7026 14116
rect 7042 14172 7106 14176
rect 7042 14116 7046 14172
rect 7046 14116 7102 14172
rect 7102 14116 7106 14172
rect 7042 14112 7106 14116
rect 7122 14172 7186 14176
rect 7122 14116 7126 14172
rect 7126 14116 7182 14172
rect 7182 14116 7186 14172
rect 7122 14112 7186 14116
rect 12813 14172 12877 14176
rect 12813 14116 12817 14172
rect 12817 14116 12873 14172
rect 12873 14116 12877 14172
rect 12813 14112 12877 14116
rect 12893 14172 12957 14176
rect 12893 14116 12897 14172
rect 12897 14116 12953 14172
rect 12953 14116 12957 14172
rect 12893 14112 12957 14116
rect 12973 14172 13037 14176
rect 12973 14116 12977 14172
rect 12977 14116 13033 14172
rect 13033 14116 13037 14172
rect 12973 14112 13037 14116
rect 13053 14172 13117 14176
rect 13053 14116 13057 14172
rect 13057 14116 13113 14172
rect 13113 14116 13117 14172
rect 13053 14112 13117 14116
rect 3917 13628 3981 13632
rect 3917 13572 3921 13628
rect 3921 13572 3977 13628
rect 3977 13572 3981 13628
rect 3917 13568 3981 13572
rect 3997 13628 4061 13632
rect 3997 13572 4001 13628
rect 4001 13572 4057 13628
rect 4057 13572 4061 13628
rect 3997 13568 4061 13572
rect 4077 13628 4141 13632
rect 4077 13572 4081 13628
rect 4081 13572 4137 13628
rect 4137 13572 4141 13628
rect 4077 13568 4141 13572
rect 4157 13628 4221 13632
rect 4157 13572 4161 13628
rect 4161 13572 4217 13628
rect 4217 13572 4221 13628
rect 4157 13568 4221 13572
rect 9848 13628 9912 13632
rect 9848 13572 9852 13628
rect 9852 13572 9908 13628
rect 9908 13572 9912 13628
rect 9848 13568 9912 13572
rect 9928 13628 9992 13632
rect 9928 13572 9932 13628
rect 9932 13572 9988 13628
rect 9988 13572 9992 13628
rect 9928 13568 9992 13572
rect 10008 13628 10072 13632
rect 10008 13572 10012 13628
rect 10012 13572 10068 13628
rect 10068 13572 10072 13628
rect 10008 13568 10072 13572
rect 10088 13628 10152 13632
rect 10088 13572 10092 13628
rect 10092 13572 10148 13628
rect 10148 13572 10152 13628
rect 10088 13568 10152 13572
rect 15778 13628 15842 13632
rect 15778 13572 15782 13628
rect 15782 13572 15838 13628
rect 15838 13572 15842 13628
rect 15778 13568 15842 13572
rect 15858 13628 15922 13632
rect 15858 13572 15862 13628
rect 15862 13572 15918 13628
rect 15918 13572 15922 13628
rect 15858 13568 15922 13572
rect 15938 13628 16002 13632
rect 15938 13572 15942 13628
rect 15942 13572 15998 13628
rect 15998 13572 16002 13628
rect 15938 13568 16002 13572
rect 16018 13628 16082 13632
rect 16018 13572 16022 13628
rect 16022 13572 16078 13628
rect 16078 13572 16082 13628
rect 16018 13568 16082 13572
rect 6882 13084 6946 13088
rect 6882 13028 6886 13084
rect 6886 13028 6942 13084
rect 6942 13028 6946 13084
rect 6882 13024 6946 13028
rect 6962 13084 7026 13088
rect 6962 13028 6966 13084
rect 6966 13028 7022 13084
rect 7022 13028 7026 13084
rect 6962 13024 7026 13028
rect 7042 13084 7106 13088
rect 7042 13028 7046 13084
rect 7046 13028 7102 13084
rect 7102 13028 7106 13084
rect 7042 13024 7106 13028
rect 7122 13084 7186 13088
rect 7122 13028 7126 13084
rect 7126 13028 7182 13084
rect 7182 13028 7186 13084
rect 7122 13024 7186 13028
rect 12813 13084 12877 13088
rect 12813 13028 12817 13084
rect 12817 13028 12873 13084
rect 12873 13028 12877 13084
rect 12813 13024 12877 13028
rect 12893 13084 12957 13088
rect 12893 13028 12897 13084
rect 12897 13028 12953 13084
rect 12953 13028 12957 13084
rect 12893 13024 12957 13028
rect 12973 13084 13037 13088
rect 12973 13028 12977 13084
rect 12977 13028 13033 13084
rect 13033 13028 13037 13084
rect 12973 13024 13037 13028
rect 13053 13084 13117 13088
rect 13053 13028 13057 13084
rect 13057 13028 13113 13084
rect 13113 13028 13117 13084
rect 13053 13024 13117 13028
rect 3917 12540 3981 12544
rect 3917 12484 3921 12540
rect 3921 12484 3977 12540
rect 3977 12484 3981 12540
rect 3917 12480 3981 12484
rect 3997 12540 4061 12544
rect 3997 12484 4001 12540
rect 4001 12484 4057 12540
rect 4057 12484 4061 12540
rect 3997 12480 4061 12484
rect 4077 12540 4141 12544
rect 4077 12484 4081 12540
rect 4081 12484 4137 12540
rect 4137 12484 4141 12540
rect 4077 12480 4141 12484
rect 4157 12540 4221 12544
rect 4157 12484 4161 12540
rect 4161 12484 4217 12540
rect 4217 12484 4221 12540
rect 4157 12480 4221 12484
rect 9848 12540 9912 12544
rect 9848 12484 9852 12540
rect 9852 12484 9908 12540
rect 9908 12484 9912 12540
rect 9848 12480 9912 12484
rect 9928 12540 9992 12544
rect 9928 12484 9932 12540
rect 9932 12484 9988 12540
rect 9988 12484 9992 12540
rect 9928 12480 9992 12484
rect 10008 12540 10072 12544
rect 10008 12484 10012 12540
rect 10012 12484 10068 12540
rect 10068 12484 10072 12540
rect 10008 12480 10072 12484
rect 10088 12540 10152 12544
rect 10088 12484 10092 12540
rect 10092 12484 10148 12540
rect 10148 12484 10152 12540
rect 10088 12480 10152 12484
rect 15778 12540 15842 12544
rect 15778 12484 15782 12540
rect 15782 12484 15838 12540
rect 15838 12484 15842 12540
rect 15778 12480 15842 12484
rect 15858 12540 15922 12544
rect 15858 12484 15862 12540
rect 15862 12484 15918 12540
rect 15918 12484 15922 12540
rect 15858 12480 15922 12484
rect 15938 12540 16002 12544
rect 15938 12484 15942 12540
rect 15942 12484 15998 12540
rect 15998 12484 16002 12540
rect 15938 12480 16002 12484
rect 16018 12540 16082 12544
rect 16018 12484 16022 12540
rect 16022 12484 16078 12540
rect 16078 12484 16082 12540
rect 16018 12480 16082 12484
rect 6882 11996 6946 12000
rect 6882 11940 6886 11996
rect 6886 11940 6942 11996
rect 6942 11940 6946 11996
rect 6882 11936 6946 11940
rect 6962 11996 7026 12000
rect 6962 11940 6966 11996
rect 6966 11940 7022 11996
rect 7022 11940 7026 11996
rect 6962 11936 7026 11940
rect 7042 11996 7106 12000
rect 7042 11940 7046 11996
rect 7046 11940 7102 11996
rect 7102 11940 7106 11996
rect 7042 11936 7106 11940
rect 7122 11996 7186 12000
rect 7122 11940 7126 11996
rect 7126 11940 7182 11996
rect 7182 11940 7186 11996
rect 7122 11936 7186 11940
rect 12813 11996 12877 12000
rect 12813 11940 12817 11996
rect 12817 11940 12873 11996
rect 12873 11940 12877 11996
rect 12813 11936 12877 11940
rect 12893 11996 12957 12000
rect 12893 11940 12897 11996
rect 12897 11940 12953 11996
rect 12953 11940 12957 11996
rect 12893 11936 12957 11940
rect 12973 11996 13037 12000
rect 12973 11940 12977 11996
rect 12977 11940 13033 11996
rect 13033 11940 13037 11996
rect 12973 11936 13037 11940
rect 13053 11996 13117 12000
rect 13053 11940 13057 11996
rect 13057 11940 13113 11996
rect 13113 11940 13117 11996
rect 13053 11936 13117 11940
rect 3917 11452 3981 11456
rect 3917 11396 3921 11452
rect 3921 11396 3977 11452
rect 3977 11396 3981 11452
rect 3917 11392 3981 11396
rect 3997 11452 4061 11456
rect 3997 11396 4001 11452
rect 4001 11396 4057 11452
rect 4057 11396 4061 11452
rect 3997 11392 4061 11396
rect 4077 11452 4141 11456
rect 4077 11396 4081 11452
rect 4081 11396 4137 11452
rect 4137 11396 4141 11452
rect 4077 11392 4141 11396
rect 4157 11452 4221 11456
rect 4157 11396 4161 11452
rect 4161 11396 4217 11452
rect 4217 11396 4221 11452
rect 4157 11392 4221 11396
rect 9848 11452 9912 11456
rect 9848 11396 9852 11452
rect 9852 11396 9908 11452
rect 9908 11396 9912 11452
rect 9848 11392 9912 11396
rect 9928 11452 9992 11456
rect 9928 11396 9932 11452
rect 9932 11396 9988 11452
rect 9988 11396 9992 11452
rect 9928 11392 9992 11396
rect 10008 11452 10072 11456
rect 10008 11396 10012 11452
rect 10012 11396 10068 11452
rect 10068 11396 10072 11452
rect 10008 11392 10072 11396
rect 10088 11452 10152 11456
rect 10088 11396 10092 11452
rect 10092 11396 10148 11452
rect 10148 11396 10152 11452
rect 10088 11392 10152 11396
rect 15778 11452 15842 11456
rect 15778 11396 15782 11452
rect 15782 11396 15838 11452
rect 15838 11396 15842 11452
rect 15778 11392 15842 11396
rect 15858 11452 15922 11456
rect 15858 11396 15862 11452
rect 15862 11396 15918 11452
rect 15918 11396 15922 11452
rect 15858 11392 15922 11396
rect 15938 11452 16002 11456
rect 15938 11396 15942 11452
rect 15942 11396 15998 11452
rect 15998 11396 16002 11452
rect 15938 11392 16002 11396
rect 16018 11452 16082 11456
rect 16018 11396 16022 11452
rect 16022 11396 16078 11452
rect 16078 11396 16082 11452
rect 16018 11392 16082 11396
rect 15148 11052 15212 11116
rect 6882 10908 6946 10912
rect 6882 10852 6886 10908
rect 6886 10852 6942 10908
rect 6942 10852 6946 10908
rect 6882 10848 6946 10852
rect 6962 10908 7026 10912
rect 6962 10852 6966 10908
rect 6966 10852 7022 10908
rect 7022 10852 7026 10908
rect 6962 10848 7026 10852
rect 7042 10908 7106 10912
rect 7042 10852 7046 10908
rect 7046 10852 7102 10908
rect 7102 10852 7106 10908
rect 7042 10848 7106 10852
rect 7122 10908 7186 10912
rect 7122 10852 7126 10908
rect 7126 10852 7182 10908
rect 7182 10852 7186 10908
rect 7122 10848 7186 10852
rect 12813 10908 12877 10912
rect 12813 10852 12817 10908
rect 12817 10852 12873 10908
rect 12873 10852 12877 10908
rect 12813 10848 12877 10852
rect 12893 10908 12957 10912
rect 12893 10852 12897 10908
rect 12897 10852 12953 10908
rect 12953 10852 12957 10908
rect 12893 10848 12957 10852
rect 12973 10908 13037 10912
rect 12973 10852 12977 10908
rect 12977 10852 13033 10908
rect 13033 10852 13037 10908
rect 12973 10848 13037 10852
rect 13053 10908 13117 10912
rect 13053 10852 13057 10908
rect 13057 10852 13113 10908
rect 13113 10852 13117 10908
rect 13053 10848 13117 10852
rect 3917 10364 3981 10368
rect 3917 10308 3921 10364
rect 3921 10308 3977 10364
rect 3977 10308 3981 10364
rect 3917 10304 3981 10308
rect 3997 10364 4061 10368
rect 3997 10308 4001 10364
rect 4001 10308 4057 10364
rect 4057 10308 4061 10364
rect 3997 10304 4061 10308
rect 4077 10364 4141 10368
rect 4077 10308 4081 10364
rect 4081 10308 4137 10364
rect 4137 10308 4141 10364
rect 4077 10304 4141 10308
rect 4157 10364 4221 10368
rect 4157 10308 4161 10364
rect 4161 10308 4217 10364
rect 4217 10308 4221 10364
rect 4157 10304 4221 10308
rect 9848 10364 9912 10368
rect 9848 10308 9852 10364
rect 9852 10308 9908 10364
rect 9908 10308 9912 10364
rect 9848 10304 9912 10308
rect 9928 10364 9992 10368
rect 9928 10308 9932 10364
rect 9932 10308 9988 10364
rect 9988 10308 9992 10364
rect 9928 10304 9992 10308
rect 10008 10364 10072 10368
rect 10008 10308 10012 10364
rect 10012 10308 10068 10364
rect 10068 10308 10072 10364
rect 10008 10304 10072 10308
rect 10088 10364 10152 10368
rect 10088 10308 10092 10364
rect 10092 10308 10148 10364
rect 10148 10308 10152 10364
rect 10088 10304 10152 10308
rect 15778 10364 15842 10368
rect 15778 10308 15782 10364
rect 15782 10308 15838 10364
rect 15838 10308 15842 10364
rect 15778 10304 15842 10308
rect 15858 10364 15922 10368
rect 15858 10308 15862 10364
rect 15862 10308 15918 10364
rect 15918 10308 15922 10364
rect 15858 10304 15922 10308
rect 15938 10364 16002 10368
rect 15938 10308 15942 10364
rect 15942 10308 15998 10364
rect 15998 10308 16002 10364
rect 15938 10304 16002 10308
rect 16018 10364 16082 10368
rect 16018 10308 16022 10364
rect 16022 10308 16078 10364
rect 16078 10308 16082 10364
rect 16018 10304 16082 10308
rect 7420 10100 7484 10164
rect 6882 9820 6946 9824
rect 6882 9764 6886 9820
rect 6886 9764 6942 9820
rect 6942 9764 6946 9820
rect 6882 9760 6946 9764
rect 6962 9820 7026 9824
rect 6962 9764 6966 9820
rect 6966 9764 7022 9820
rect 7022 9764 7026 9820
rect 6962 9760 7026 9764
rect 7042 9820 7106 9824
rect 7042 9764 7046 9820
rect 7046 9764 7102 9820
rect 7102 9764 7106 9820
rect 7042 9760 7106 9764
rect 7122 9820 7186 9824
rect 7122 9764 7126 9820
rect 7126 9764 7182 9820
rect 7182 9764 7186 9820
rect 7122 9760 7186 9764
rect 12813 9820 12877 9824
rect 12813 9764 12817 9820
rect 12817 9764 12873 9820
rect 12873 9764 12877 9820
rect 12813 9760 12877 9764
rect 12893 9820 12957 9824
rect 12893 9764 12897 9820
rect 12897 9764 12953 9820
rect 12953 9764 12957 9820
rect 12893 9760 12957 9764
rect 12973 9820 13037 9824
rect 12973 9764 12977 9820
rect 12977 9764 13033 9820
rect 13033 9764 13037 9820
rect 12973 9760 13037 9764
rect 13053 9820 13117 9824
rect 13053 9764 13057 9820
rect 13057 9764 13113 9820
rect 13113 9764 13117 9820
rect 13053 9760 13117 9764
rect 3917 9276 3981 9280
rect 3917 9220 3921 9276
rect 3921 9220 3977 9276
rect 3977 9220 3981 9276
rect 3917 9216 3981 9220
rect 3997 9276 4061 9280
rect 3997 9220 4001 9276
rect 4001 9220 4057 9276
rect 4057 9220 4061 9276
rect 3997 9216 4061 9220
rect 4077 9276 4141 9280
rect 4077 9220 4081 9276
rect 4081 9220 4137 9276
rect 4137 9220 4141 9276
rect 4077 9216 4141 9220
rect 4157 9276 4221 9280
rect 4157 9220 4161 9276
rect 4161 9220 4217 9276
rect 4217 9220 4221 9276
rect 4157 9216 4221 9220
rect 9848 9276 9912 9280
rect 9848 9220 9852 9276
rect 9852 9220 9908 9276
rect 9908 9220 9912 9276
rect 9848 9216 9912 9220
rect 9928 9276 9992 9280
rect 9928 9220 9932 9276
rect 9932 9220 9988 9276
rect 9988 9220 9992 9276
rect 9928 9216 9992 9220
rect 10008 9276 10072 9280
rect 10008 9220 10012 9276
rect 10012 9220 10068 9276
rect 10068 9220 10072 9276
rect 10008 9216 10072 9220
rect 10088 9276 10152 9280
rect 10088 9220 10092 9276
rect 10092 9220 10148 9276
rect 10148 9220 10152 9276
rect 10088 9216 10152 9220
rect 15778 9276 15842 9280
rect 15778 9220 15782 9276
rect 15782 9220 15838 9276
rect 15838 9220 15842 9276
rect 15778 9216 15842 9220
rect 15858 9276 15922 9280
rect 15858 9220 15862 9276
rect 15862 9220 15918 9276
rect 15918 9220 15922 9276
rect 15858 9216 15922 9220
rect 15938 9276 16002 9280
rect 15938 9220 15942 9276
rect 15942 9220 15998 9276
rect 15998 9220 16002 9276
rect 15938 9216 16002 9220
rect 16018 9276 16082 9280
rect 16018 9220 16022 9276
rect 16022 9220 16078 9276
rect 16078 9220 16082 9276
rect 16018 9216 16082 9220
rect 6882 8732 6946 8736
rect 6882 8676 6886 8732
rect 6886 8676 6942 8732
rect 6942 8676 6946 8732
rect 6882 8672 6946 8676
rect 6962 8732 7026 8736
rect 6962 8676 6966 8732
rect 6966 8676 7022 8732
rect 7022 8676 7026 8732
rect 6962 8672 7026 8676
rect 7042 8732 7106 8736
rect 7042 8676 7046 8732
rect 7046 8676 7102 8732
rect 7102 8676 7106 8732
rect 7042 8672 7106 8676
rect 7122 8732 7186 8736
rect 7122 8676 7126 8732
rect 7126 8676 7182 8732
rect 7182 8676 7186 8732
rect 7122 8672 7186 8676
rect 12813 8732 12877 8736
rect 12813 8676 12817 8732
rect 12817 8676 12873 8732
rect 12873 8676 12877 8732
rect 12813 8672 12877 8676
rect 12893 8732 12957 8736
rect 12893 8676 12897 8732
rect 12897 8676 12953 8732
rect 12953 8676 12957 8732
rect 12893 8672 12957 8676
rect 12973 8732 13037 8736
rect 12973 8676 12977 8732
rect 12977 8676 13033 8732
rect 13033 8676 13037 8732
rect 12973 8672 13037 8676
rect 13053 8732 13117 8736
rect 13053 8676 13057 8732
rect 13057 8676 13113 8732
rect 13113 8676 13117 8732
rect 13053 8672 13117 8676
rect 14044 8528 14108 8532
rect 14044 8472 14058 8528
rect 14058 8472 14108 8528
rect 14044 8468 14108 8472
rect 3917 8188 3981 8192
rect 3917 8132 3921 8188
rect 3921 8132 3977 8188
rect 3977 8132 3981 8188
rect 3917 8128 3981 8132
rect 3997 8188 4061 8192
rect 3997 8132 4001 8188
rect 4001 8132 4057 8188
rect 4057 8132 4061 8188
rect 3997 8128 4061 8132
rect 4077 8188 4141 8192
rect 4077 8132 4081 8188
rect 4081 8132 4137 8188
rect 4137 8132 4141 8188
rect 4077 8128 4141 8132
rect 4157 8188 4221 8192
rect 4157 8132 4161 8188
rect 4161 8132 4217 8188
rect 4217 8132 4221 8188
rect 4157 8128 4221 8132
rect 9848 8188 9912 8192
rect 9848 8132 9852 8188
rect 9852 8132 9908 8188
rect 9908 8132 9912 8188
rect 9848 8128 9912 8132
rect 9928 8188 9992 8192
rect 9928 8132 9932 8188
rect 9932 8132 9988 8188
rect 9988 8132 9992 8188
rect 9928 8128 9992 8132
rect 10008 8188 10072 8192
rect 10008 8132 10012 8188
rect 10012 8132 10068 8188
rect 10068 8132 10072 8188
rect 10008 8128 10072 8132
rect 10088 8188 10152 8192
rect 10088 8132 10092 8188
rect 10092 8132 10148 8188
rect 10148 8132 10152 8188
rect 10088 8128 10152 8132
rect 15778 8188 15842 8192
rect 15778 8132 15782 8188
rect 15782 8132 15838 8188
rect 15838 8132 15842 8188
rect 15778 8128 15842 8132
rect 15858 8188 15922 8192
rect 15858 8132 15862 8188
rect 15862 8132 15918 8188
rect 15918 8132 15922 8188
rect 15858 8128 15922 8132
rect 15938 8188 16002 8192
rect 15938 8132 15942 8188
rect 15942 8132 15998 8188
rect 15998 8132 16002 8188
rect 15938 8128 16002 8132
rect 16018 8188 16082 8192
rect 16018 8132 16022 8188
rect 16022 8132 16078 8188
rect 16078 8132 16082 8188
rect 16018 8128 16082 8132
rect 6882 7644 6946 7648
rect 6882 7588 6886 7644
rect 6886 7588 6942 7644
rect 6942 7588 6946 7644
rect 6882 7584 6946 7588
rect 6962 7644 7026 7648
rect 6962 7588 6966 7644
rect 6966 7588 7022 7644
rect 7022 7588 7026 7644
rect 6962 7584 7026 7588
rect 7042 7644 7106 7648
rect 7042 7588 7046 7644
rect 7046 7588 7102 7644
rect 7102 7588 7106 7644
rect 7042 7584 7106 7588
rect 7122 7644 7186 7648
rect 7122 7588 7126 7644
rect 7126 7588 7182 7644
rect 7182 7588 7186 7644
rect 7122 7584 7186 7588
rect 12813 7644 12877 7648
rect 12813 7588 12817 7644
rect 12817 7588 12873 7644
rect 12873 7588 12877 7644
rect 12813 7584 12877 7588
rect 12893 7644 12957 7648
rect 12893 7588 12897 7644
rect 12897 7588 12953 7644
rect 12953 7588 12957 7644
rect 12893 7584 12957 7588
rect 12973 7644 13037 7648
rect 12973 7588 12977 7644
rect 12977 7588 13033 7644
rect 13033 7588 13037 7644
rect 12973 7584 13037 7588
rect 13053 7644 13117 7648
rect 13053 7588 13057 7644
rect 13057 7588 13113 7644
rect 13113 7588 13117 7644
rect 13053 7584 13117 7588
rect 3917 7100 3981 7104
rect 3917 7044 3921 7100
rect 3921 7044 3977 7100
rect 3977 7044 3981 7100
rect 3917 7040 3981 7044
rect 3997 7100 4061 7104
rect 3997 7044 4001 7100
rect 4001 7044 4057 7100
rect 4057 7044 4061 7100
rect 3997 7040 4061 7044
rect 4077 7100 4141 7104
rect 4077 7044 4081 7100
rect 4081 7044 4137 7100
rect 4137 7044 4141 7100
rect 4077 7040 4141 7044
rect 4157 7100 4221 7104
rect 4157 7044 4161 7100
rect 4161 7044 4217 7100
rect 4217 7044 4221 7100
rect 4157 7040 4221 7044
rect 9848 7100 9912 7104
rect 9848 7044 9852 7100
rect 9852 7044 9908 7100
rect 9908 7044 9912 7100
rect 9848 7040 9912 7044
rect 9928 7100 9992 7104
rect 9928 7044 9932 7100
rect 9932 7044 9988 7100
rect 9988 7044 9992 7100
rect 9928 7040 9992 7044
rect 10008 7100 10072 7104
rect 10008 7044 10012 7100
rect 10012 7044 10068 7100
rect 10068 7044 10072 7100
rect 10008 7040 10072 7044
rect 10088 7100 10152 7104
rect 10088 7044 10092 7100
rect 10092 7044 10148 7100
rect 10148 7044 10152 7100
rect 10088 7040 10152 7044
rect 15778 7100 15842 7104
rect 15778 7044 15782 7100
rect 15782 7044 15838 7100
rect 15838 7044 15842 7100
rect 15778 7040 15842 7044
rect 15858 7100 15922 7104
rect 15858 7044 15862 7100
rect 15862 7044 15918 7100
rect 15918 7044 15922 7100
rect 15858 7040 15922 7044
rect 15938 7100 16002 7104
rect 15938 7044 15942 7100
rect 15942 7044 15998 7100
rect 15998 7044 16002 7100
rect 15938 7040 16002 7044
rect 16018 7100 16082 7104
rect 16018 7044 16022 7100
rect 16022 7044 16078 7100
rect 16078 7044 16082 7100
rect 16018 7040 16082 7044
rect 12388 6972 12452 7036
rect 15148 6564 15212 6628
rect 6882 6556 6946 6560
rect 6882 6500 6886 6556
rect 6886 6500 6942 6556
rect 6942 6500 6946 6556
rect 6882 6496 6946 6500
rect 6962 6556 7026 6560
rect 6962 6500 6966 6556
rect 6966 6500 7022 6556
rect 7022 6500 7026 6556
rect 6962 6496 7026 6500
rect 7042 6556 7106 6560
rect 7042 6500 7046 6556
rect 7046 6500 7102 6556
rect 7102 6500 7106 6556
rect 7042 6496 7106 6500
rect 7122 6556 7186 6560
rect 7122 6500 7126 6556
rect 7126 6500 7182 6556
rect 7182 6500 7186 6556
rect 7122 6496 7186 6500
rect 12813 6556 12877 6560
rect 12813 6500 12817 6556
rect 12817 6500 12873 6556
rect 12873 6500 12877 6556
rect 12813 6496 12877 6500
rect 12893 6556 12957 6560
rect 12893 6500 12897 6556
rect 12897 6500 12953 6556
rect 12953 6500 12957 6556
rect 12893 6496 12957 6500
rect 12973 6556 13037 6560
rect 12973 6500 12977 6556
rect 12977 6500 13033 6556
rect 13033 6500 13037 6556
rect 12973 6496 13037 6500
rect 13053 6556 13117 6560
rect 13053 6500 13057 6556
rect 13057 6500 13113 6556
rect 13113 6500 13117 6556
rect 13053 6496 13117 6500
rect 12388 6428 12452 6492
rect 3917 6012 3981 6016
rect 3917 5956 3921 6012
rect 3921 5956 3977 6012
rect 3977 5956 3981 6012
rect 3917 5952 3981 5956
rect 3997 6012 4061 6016
rect 3997 5956 4001 6012
rect 4001 5956 4057 6012
rect 4057 5956 4061 6012
rect 3997 5952 4061 5956
rect 4077 6012 4141 6016
rect 4077 5956 4081 6012
rect 4081 5956 4137 6012
rect 4137 5956 4141 6012
rect 4077 5952 4141 5956
rect 4157 6012 4221 6016
rect 4157 5956 4161 6012
rect 4161 5956 4217 6012
rect 4217 5956 4221 6012
rect 4157 5952 4221 5956
rect 9848 6012 9912 6016
rect 9848 5956 9852 6012
rect 9852 5956 9908 6012
rect 9908 5956 9912 6012
rect 9848 5952 9912 5956
rect 9928 6012 9992 6016
rect 9928 5956 9932 6012
rect 9932 5956 9988 6012
rect 9988 5956 9992 6012
rect 9928 5952 9992 5956
rect 10008 6012 10072 6016
rect 10008 5956 10012 6012
rect 10012 5956 10068 6012
rect 10068 5956 10072 6012
rect 10008 5952 10072 5956
rect 10088 6012 10152 6016
rect 10088 5956 10092 6012
rect 10092 5956 10148 6012
rect 10148 5956 10152 6012
rect 10088 5952 10152 5956
rect 15778 6012 15842 6016
rect 15778 5956 15782 6012
rect 15782 5956 15838 6012
rect 15838 5956 15842 6012
rect 15778 5952 15842 5956
rect 15858 6012 15922 6016
rect 15858 5956 15862 6012
rect 15862 5956 15918 6012
rect 15918 5956 15922 6012
rect 15858 5952 15922 5956
rect 15938 6012 16002 6016
rect 15938 5956 15942 6012
rect 15942 5956 15998 6012
rect 15998 5956 16002 6012
rect 15938 5952 16002 5956
rect 16018 6012 16082 6016
rect 16018 5956 16022 6012
rect 16022 5956 16078 6012
rect 16078 5956 16082 6012
rect 16018 5952 16082 5956
rect 14044 5476 14108 5540
rect 6882 5468 6946 5472
rect 6882 5412 6886 5468
rect 6886 5412 6942 5468
rect 6942 5412 6946 5468
rect 6882 5408 6946 5412
rect 6962 5468 7026 5472
rect 6962 5412 6966 5468
rect 6966 5412 7022 5468
rect 7022 5412 7026 5468
rect 6962 5408 7026 5412
rect 7042 5468 7106 5472
rect 7042 5412 7046 5468
rect 7046 5412 7102 5468
rect 7102 5412 7106 5468
rect 7042 5408 7106 5412
rect 7122 5468 7186 5472
rect 7122 5412 7126 5468
rect 7126 5412 7182 5468
rect 7182 5412 7186 5468
rect 7122 5408 7186 5412
rect 12813 5468 12877 5472
rect 12813 5412 12817 5468
rect 12817 5412 12873 5468
rect 12873 5412 12877 5468
rect 12813 5408 12877 5412
rect 12893 5468 12957 5472
rect 12893 5412 12897 5468
rect 12897 5412 12953 5468
rect 12953 5412 12957 5468
rect 12893 5408 12957 5412
rect 12973 5468 13037 5472
rect 12973 5412 12977 5468
rect 12977 5412 13033 5468
rect 13033 5412 13037 5468
rect 12973 5408 13037 5412
rect 13053 5468 13117 5472
rect 13053 5412 13057 5468
rect 13057 5412 13113 5468
rect 13113 5412 13117 5468
rect 13053 5408 13117 5412
rect 3917 4924 3981 4928
rect 3917 4868 3921 4924
rect 3921 4868 3977 4924
rect 3977 4868 3981 4924
rect 3917 4864 3981 4868
rect 3997 4924 4061 4928
rect 3997 4868 4001 4924
rect 4001 4868 4057 4924
rect 4057 4868 4061 4924
rect 3997 4864 4061 4868
rect 4077 4924 4141 4928
rect 4077 4868 4081 4924
rect 4081 4868 4137 4924
rect 4137 4868 4141 4924
rect 4077 4864 4141 4868
rect 4157 4924 4221 4928
rect 4157 4868 4161 4924
rect 4161 4868 4217 4924
rect 4217 4868 4221 4924
rect 4157 4864 4221 4868
rect 9848 4924 9912 4928
rect 9848 4868 9852 4924
rect 9852 4868 9908 4924
rect 9908 4868 9912 4924
rect 9848 4864 9912 4868
rect 9928 4924 9992 4928
rect 9928 4868 9932 4924
rect 9932 4868 9988 4924
rect 9988 4868 9992 4924
rect 9928 4864 9992 4868
rect 10008 4924 10072 4928
rect 10008 4868 10012 4924
rect 10012 4868 10068 4924
rect 10068 4868 10072 4924
rect 10008 4864 10072 4868
rect 10088 4924 10152 4928
rect 10088 4868 10092 4924
rect 10092 4868 10148 4924
rect 10148 4868 10152 4924
rect 10088 4864 10152 4868
rect 15778 4924 15842 4928
rect 15778 4868 15782 4924
rect 15782 4868 15838 4924
rect 15838 4868 15842 4924
rect 15778 4864 15842 4868
rect 15858 4924 15922 4928
rect 15858 4868 15862 4924
rect 15862 4868 15918 4924
rect 15918 4868 15922 4924
rect 15858 4864 15922 4868
rect 15938 4924 16002 4928
rect 15938 4868 15942 4924
rect 15942 4868 15998 4924
rect 15998 4868 16002 4924
rect 15938 4864 16002 4868
rect 16018 4924 16082 4928
rect 16018 4868 16022 4924
rect 16022 4868 16078 4924
rect 16078 4868 16082 4924
rect 16018 4864 16082 4868
rect 6882 4380 6946 4384
rect 6882 4324 6886 4380
rect 6886 4324 6942 4380
rect 6942 4324 6946 4380
rect 6882 4320 6946 4324
rect 6962 4380 7026 4384
rect 6962 4324 6966 4380
rect 6966 4324 7022 4380
rect 7022 4324 7026 4380
rect 6962 4320 7026 4324
rect 7042 4380 7106 4384
rect 7042 4324 7046 4380
rect 7046 4324 7102 4380
rect 7102 4324 7106 4380
rect 7042 4320 7106 4324
rect 7122 4380 7186 4384
rect 7122 4324 7126 4380
rect 7126 4324 7182 4380
rect 7182 4324 7186 4380
rect 7122 4320 7186 4324
rect 12813 4380 12877 4384
rect 12813 4324 12817 4380
rect 12817 4324 12873 4380
rect 12873 4324 12877 4380
rect 12813 4320 12877 4324
rect 12893 4380 12957 4384
rect 12893 4324 12897 4380
rect 12897 4324 12953 4380
rect 12953 4324 12957 4380
rect 12893 4320 12957 4324
rect 12973 4380 13037 4384
rect 12973 4324 12977 4380
rect 12977 4324 13033 4380
rect 13033 4324 13037 4380
rect 12973 4320 13037 4324
rect 13053 4380 13117 4384
rect 13053 4324 13057 4380
rect 13057 4324 13113 4380
rect 13113 4324 13117 4380
rect 13053 4320 13117 4324
rect 3917 3836 3981 3840
rect 3917 3780 3921 3836
rect 3921 3780 3977 3836
rect 3977 3780 3981 3836
rect 3917 3776 3981 3780
rect 3997 3836 4061 3840
rect 3997 3780 4001 3836
rect 4001 3780 4057 3836
rect 4057 3780 4061 3836
rect 3997 3776 4061 3780
rect 4077 3836 4141 3840
rect 4077 3780 4081 3836
rect 4081 3780 4137 3836
rect 4137 3780 4141 3836
rect 4077 3776 4141 3780
rect 4157 3836 4221 3840
rect 4157 3780 4161 3836
rect 4161 3780 4217 3836
rect 4217 3780 4221 3836
rect 4157 3776 4221 3780
rect 9848 3836 9912 3840
rect 9848 3780 9852 3836
rect 9852 3780 9908 3836
rect 9908 3780 9912 3836
rect 9848 3776 9912 3780
rect 9928 3836 9992 3840
rect 9928 3780 9932 3836
rect 9932 3780 9988 3836
rect 9988 3780 9992 3836
rect 9928 3776 9992 3780
rect 10008 3836 10072 3840
rect 10008 3780 10012 3836
rect 10012 3780 10068 3836
rect 10068 3780 10072 3836
rect 10008 3776 10072 3780
rect 10088 3836 10152 3840
rect 10088 3780 10092 3836
rect 10092 3780 10148 3836
rect 10148 3780 10152 3836
rect 10088 3776 10152 3780
rect 15778 3836 15842 3840
rect 15778 3780 15782 3836
rect 15782 3780 15838 3836
rect 15838 3780 15842 3836
rect 15778 3776 15842 3780
rect 15858 3836 15922 3840
rect 15858 3780 15862 3836
rect 15862 3780 15918 3836
rect 15918 3780 15922 3836
rect 15858 3776 15922 3780
rect 15938 3836 16002 3840
rect 15938 3780 15942 3836
rect 15942 3780 15998 3836
rect 15998 3780 16002 3836
rect 15938 3776 16002 3780
rect 16018 3836 16082 3840
rect 16018 3780 16022 3836
rect 16022 3780 16078 3836
rect 16078 3780 16082 3836
rect 16018 3776 16082 3780
rect 6882 3292 6946 3296
rect 6882 3236 6886 3292
rect 6886 3236 6942 3292
rect 6942 3236 6946 3292
rect 6882 3232 6946 3236
rect 6962 3292 7026 3296
rect 6962 3236 6966 3292
rect 6966 3236 7022 3292
rect 7022 3236 7026 3292
rect 6962 3232 7026 3236
rect 7042 3292 7106 3296
rect 7042 3236 7046 3292
rect 7046 3236 7102 3292
rect 7102 3236 7106 3292
rect 7042 3232 7106 3236
rect 7122 3292 7186 3296
rect 7122 3236 7126 3292
rect 7126 3236 7182 3292
rect 7182 3236 7186 3292
rect 7122 3232 7186 3236
rect 12813 3292 12877 3296
rect 12813 3236 12817 3292
rect 12817 3236 12873 3292
rect 12873 3236 12877 3292
rect 12813 3232 12877 3236
rect 12893 3292 12957 3296
rect 12893 3236 12897 3292
rect 12897 3236 12953 3292
rect 12953 3236 12957 3292
rect 12893 3232 12957 3236
rect 12973 3292 13037 3296
rect 12973 3236 12977 3292
rect 12977 3236 13033 3292
rect 13033 3236 13037 3292
rect 12973 3232 13037 3236
rect 13053 3292 13117 3296
rect 13053 3236 13057 3292
rect 13057 3236 13113 3292
rect 13113 3236 13117 3292
rect 13053 3232 13117 3236
rect 3917 2748 3981 2752
rect 3917 2692 3921 2748
rect 3921 2692 3977 2748
rect 3977 2692 3981 2748
rect 3917 2688 3981 2692
rect 3997 2748 4061 2752
rect 3997 2692 4001 2748
rect 4001 2692 4057 2748
rect 4057 2692 4061 2748
rect 3997 2688 4061 2692
rect 4077 2748 4141 2752
rect 4077 2692 4081 2748
rect 4081 2692 4137 2748
rect 4137 2692 4141 2748
rect 4077 2688 4141 2692
rect 4157 2748 4221 2752
rect 4157 2692 4161 2748
rect 4161 2692 4217 2748
rect 4217 2692 4221 2748
rect 4157 2688 4221 2692
rect 9848 2748 9912 2752
rect 9848 2692 9852 2748
rect 9852 2692 9908 2748
rect 9908 2692 9912 2748
rect 9848 2688 9912 2692
rect 9928 2748 9992 2752
rect 9928 2692 9932 2748
rect 9932 2692 9988 2748
rect 9988 2692 9992 2748
rect 9928 2688 9992 2692
rect 10008 2748 10072 2752
rect 10008 2692 10012 2748
rect 10012 2692 10068 2748
rect 10068 2692 10072 2748
rect 10008 2688 10072 2692
rect 10088 2748 10152 2752
rect 10088 2692 10092 2748
rect 10092 2692 10148 2748
rect 10148 2692 10152 2748
rect 10088 2688 10152 2692
rect 15778 2748 15842 2752
rect 15778 2692 15782 2748
rect 15782 2692 15838 2748
rect 15838 2692 15842 2748
rect 15778 2688 15842 2692
rect 15858 2748 15922 2752
rect 15858 2692 15862 2748
rect 15862 2692 15918 2748
rect 15918 2692 15922 2748
rect 15858 2688 15922 2692
rect 15938 2748 16002 2752
rect 15938 2692 15942 2748
rect 15942 2692 15998 2748
rect 15998 2692 16002 2748
rect 15938 2688 16002 2692
rect 16018 2748 16082 2752
rect 16018 2692 16022 2748
rect 16022 2692 16078 2748
rect 16078 2692 16082 2748
rect 16018 2688 16082 2692
rect 6882 2204 6946 2208
rect 6882 2148 6886 2204
rect 6886 2148 6942 2204
rect 6942 2148 6946 2204
rect 6882 2144 6946 2148
rect 6962 2204 7026 2208
rect 6962 2148 6966 2204
rect 6966 2148 7022 2204
rect 7022 2148 7026 2204
rect 6962 2144 7026 2148
rect 7042 2204 7106 2208
rect 7042 2148 7046 2204
rect 7046 2148 7102 2204
rect 7102 2148 7106 2204
rect 7042 2144 7106 2148
rect 7122 2204 7186 2208
rect 7122 2148 7126 2204
rect 7126 2148 7182 2204
rect 7182 2148 7186 2204
rect 7122 2144 7186 2148
rect 12813 2204 12877 2208
rect 12813 2148 12817 2204
rect 12817 2148 12873 2204
rect 12873 2148 12877 2204
rect 12813 2144 12877 2148
rect 12893 2204 12957 2208
rect 12893 2148 12897 2204
rect 12897 2148 12953 2204
rect 12953 2148 12957 2204
rect 12893 2144 12957 2148
rect 12973 2204 13037 2208
rect 12973 2148 12977 2204
rect 12977 2148 13033 2204
rect 13033 2148 13037 2204
rect 12973 2144 13037 2148
rect 13053 2204 13117 2208
rect 13053 2148 13057 2204
rect 13057 2148 13113 2204
rect 13113 2148 13117 2204
rect 13053 2144 13117 2148
<< metal4 >>
rect 3909 16896 4230 17456
rect 3909 16832 3917 16896
rect 3981 16832 3997 16896
rect 4061 16832 4077 16896
rect 4141 16832 4157 16896
rect 4221 16832 4230 16896
rect 3909 15808 4230 16832
rect 3909 15744 3917 15808
rect 3981 15744 3997 15808
rect 4061 15744 4077 15808
rect 4141 15744 4157 15808
rect 4221 15744 4230 15808
rect 3909 14720 4230 15744
rect 3909 14656 3917 14720
rect 3981 14656 3997 14720
rect 4061 14656 4077 14720
rect 4141 14656 4157 14720
rect 4221 14656 4230 14720
rect 3909 13632 4230 14656
rect 3909 13568 3917 13632
rect 3981 13568 3997 13632
rect 4061 13568 4077 13632
rect 4141 13568 4157 13632
rect 4221 13568 4230 13632
rect 3909 12544 4230 13568
rect 3909 12480 3917 12544
rect 3981 12480 3997 12544
rect 4061 12480 4077 12544
rect 4141 12480 4157 12544
rect 4221 12480 4230 12544
rect 3909 11456 4230 12480
rect 3909 11392 3917 11456
rect 3981 11392 3997 11456
rect 4061 11392 4077 11456
rect 4141 11392 4157 11456
rect 4221 11392 4230 11456
rect 3909 10368 4230 11392
rect 3909 10304 3917 10368
rect 3981 10304 3997 10368
rect 4061 10304 4077 10368
rect 4141 10304 4157 10368
rect 4221 10304 4230 10368
rect 3909 9280 4230 10304
rect 3909 9216 3917 9280
rect 3981 9216 3997 9280
rect 4061 9216 4077 9280
rect 4141 9216 4157 9280
rect 4221 9216 4230 9280
rect 3909 8192 4230 9216
rect 3909 8128 3917 8192
rect 3981 8128 3997 8192
rect 4061 8128 4077 8192
rect 4141 8128 4157 8192
rect 4221 8128 4230 8192
rect 3909 7104 4230 8128
rect 3909 7040 3917 7104
rect 3981 7040 3997 7104
rect 4061 7040 4077 7104
rect 4141 7040 4157 7104
rect 4221 7040 4230 7104
rect 3909 6016 4230 7040
rect 3909 5952 3917 6016
rect 3981 5952 3997 6016
rect 4061 5952 4077 6016
rect 4141 5952 4157 6016
rect 4221 5952 4230 6016
rect 3909 4928 4230 5952
rect 3909 4864 3917 4928
rect 3981 4864 3997 4928
rect 4061 4864 4077 4928
rect 4141 4864 4157 4928
rect 4221 4864 4230 4928
rect 3909 3840 4230 4864
rect 3909 3776 3917 3840
rect 3981 3776 3997 3840
rect 4061 3776 4077 3840
rect 4141 3776 4157 3840
rect 4221 3776 4230 3840
rect 3909 2752 4230 3776
rect 3909 2688 3917 2752
rect 3981 2688 3997 2752
rect 4061 2688 4077 2752
rect 4141 2688 4157 2752
rect 4221 2688 4230 2752
rect 3909 2128 4230 2688
rect 6874 17440 7194 17456
rect 6874 17376 6882 17440
rect 6946 17376 6962 17440
rect 7026 17376 7042 17440
rect 7106 17376 7122 17440
rect 7186 17376 7194 17440
rect 6874 16352 7194 17376
rect 9840 16896 10160 17456
rect 9840 16832 9848 16896
rect 9912 16832 9928 16896
rect 9992 16832 10008 16896
rect 10072 16832 10088 16896
rect 10152 16832 10160 16896
rect 7419 16692 7485 16693
rect 7419 16628 7420 16692
rect 7484 16628 7485 16692
rect 7419 16627 7485 16628
rect 6874 16288 6882 16352
rect 6946 16288 6962 16352
rect 7026 16288 7042 16352
rect 7106 16288 7122 16352
rect 7186 16288 7194 16352
rect 6874 15264 7194 16288
rect 6874 15200 6882 15264
rect 6946 15200 6962 15264
rect 7026 15200 7042 15264
rect 7106 15200 7122 15264
rect 7186 15200 7194 15264
rect 6874 14176 7194 15200
rect 6874 14112 6882 14176
rect 6946 14112 6962 14176
rect 7026 14112 7042 14176
rect 7106 14112 7122 14176
rect 7186 14112 7194 14176
rect 6874 13088 7194 14112
rect 6874 13024 6882 13088
rect 6946 13024 6962 13088
rect 7026 13024 7042 13088
rect 7106 13024 7122 13088
rect 7186 13024 7194 13088
rect 6874 12000 7194 13024
rect 6874 11936 6882 12000
rect 6946 11936 6962 12000
rect 7026 11936 7042 12000
rect 7106 11936 7122 12000
rect 7186 11936 7194 12000
rect 6874 10912 7194 11936
rect 6874 10848 6882 10912
rect 6946 10848 6962 10912
rect 7026 10848 7042 10912
rect 7106 10848 7122 10912
rect 7186 10848 7194 10912
rect 6874 9824 7194 10848
rect 7422 10165 7482 16627
rect 9840 15808 10160 16832
rect 9840 15744 9848 15808
rect 9912 15744 9928 15808
rect 9992 15744 10008 15808
rect 10072 15744 10088 15808
rect 10152 15744 10160 15808
rect 9840 14720 10160 15744
rect 9840 14656 9848 14720
rect 9912 14656 9928 14720
rect 9992 14656 10008 14720
rect 10072 14656 10088 14720
rect 10152 14656 10160 14720
rect 9840 13632 10160 14656
rect 9840 13568 9848 13632
rect 9912 13568 9928 13632
rect 9992 13568 10008 13632
rect 10072 13568 10088 13632
rect 10152 13568 10160 13632
rect 9840 12544 10160 13568
rect 9840 12480 9848 12544
rect 9912 12480 9928 12544
rect 9992 12480 10008 12544
rect 10072 12480 10088 12544
rect 10152 12480 10160 12544
rect 9840 11456 10160 12480
rect 9840 11392 9848 11456
rect 9912 11392 9928 11456
rect 9992 11392 10008 11456
rect 10072 11392 10088 11456
rect 10152 11392 10160 11456
rect 9840 10368 10160 11392
rect 9840 10304 9848 10368
rect 9912 10304 9928 10368
rect 9992 10304 10008 10368
rect 10072 10304 10088 10368
rect 10152 10304 10160 10368
rect 7419 10164 7485 10165
rect 7419 10100 7420 10164
rect 7484 10100 7485 10164
rect 7419 10099 7485 10100
rect 6874 9760 6882 9824
rect 6946 9760 6962 9824
rect 7026 9760 7042 9824
rect 7106 9760 7122 9824
rect 7186 9760 7194 9824
rect 6874 8736 7194 9760
rect 6874 8672 6882 8736
rect 6946 8672 6962 8736
rect 7026 8672 7042 8736
rect 7106 8672 7122 8736
rect 7186 8672 7194 8736
rect 6874 7648 7194 8672
rect 6874 7584 6882 7648
rect 6946 7584 6962 7648
rect 7026 7584 7042 7648
rect 7106 7584 7122 7648
rect 7186 7584 7194 7648
rect 6874 6560 7194 7584
rect 6874 6496 6882 6560
rect 6946 6496 6962 6560
rect 7026 6496 7042 6560
rect 7106 6496 7122 6560
rect 7186 6496 7194 6560
rect 6874 5472 7194 6496
rect 6874 5408 6882 5472
rect 6946 5408 6962 5472
rect 7026 5408 7042 5472
rect 7106 5408 7122 5472
rect 7186 5408 7194 5472
rect 6874 4384 7194 5408
rect 6874 4320 6882 4384
rect 6946 4320 6962 4384
rect 7026 4320 7042 4384
rect 7106 4320 7122 4384
rect 7186 4320 7194 4384
rect 6874 3296 7194 4320
rect 6874 3232 6882 3296
rect 6946 3232 6962 3296
rect 7026 3232 7042 3296
rect 7106 3232 7122 3296
rect 7186 3232 7194 3296
rect 6874 2208 7194 3232
rect 6874 2144 6882 2208
rect 6946 2144 6962 2208
rect 7026 2144 7042 2208
rect 7106 2144 7122 2208
rect 7186 2144 7194 2208
rect 6874 2128 7194 2144
rect 9840 9280 10160 10304
rect 9840 9216 9848 9280
rect 9912 9216 9928 9280
rect 9992 9216 10008 9280
rect 10072 9216 10088 9280
rect 10152 9216 10160 9280
rect 9840 8192 10160 9216
rect 9840 8128 9848 8192
rect 9912 8128 9928 8192
rect 9992 8128 10008 8192
rect 10072 8128 10088 8192
rect 10152 8128 10160 8192
rect 9840 7104 10160 8128
rect 9840 7040 9848 7104
rect 9912 7040 9928 7104
rect 9992 7040 10008 7104
rect 10072 7040 10088 7104
rect 10152 7040 10160 7104
rect 9840 6016 10160 7040
rect 12805 17440 13125 17456
rect 12805 17376 12813 17440
rect 12877 17376 12893 17440
rect 12957 17376 12973 17440
rect 13037 17376 13053 17440
rect 13117 17376 13125 17440
rect 12805 16352 13125 17376
rect 12805 16288 12813 16352
rect 12877 16288 12893 16352
rect 12957 16288 12973 16352
rect 13037 16288 13053 16352
rect 13117 16288 13125 16352
rect 12805 15264 13125 16288
rect 12805 15200 12813 15264
rect 12877 15200 12893 15264
rect 12957 15200 12973 15264
rect 13037 15200 13053 15264
rect 13117 15200 13125 15264
rect 12805 14176 13125 15200
rect 12805 14112 12813 14176
rect 12877 14112 12893 14176
rect 12957 14112 12973 14176
rect 13037 14112 13053 14176
rect 13117 14112 13125 14176
rect 12805 13088 13125 14112
rect 12805 13024 12813 13088
rect 12877 13024 12893 13088
rect 12957 13024 12973 13088
rect 13037 13024 13053 13088
rect 13117 13024 13125 13088
rect 12805 12000 13125 13024
rect 12805 11936 12813 12000
rect 12877 11936 12893 12000
rect 12957 11936 12973 12000
rect 13037 11936 13053 12000
rect 13117 11936 13125 12000
rect 12805 10912 13125 11936
rect 15770 16896 16091 17456
rect 15770 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15938 16896
rect 16002 16832 16018 16896
rect 16082 16832 16091 16896
rect 15770 15808 16091 16832
rect 15770 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15938 15808
rect 16002 15744 16018 15808
rect 16082 15744 16091 15808
rect 15770 14720 16091 15744
rect 15770 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15938 14720
rect 16002 14656 16018 14720
rect 16082 14656 16091 14720
rect 15770 13632 16091 14656
rect 15770 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15938 13632
rect 16002 13568 16018 13632
rect 16082 13568 16091 13632
rect 15770 12544 16091 13568
rect 15770 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15938 12544
rect 16002 12480 16018 12544
rect 16082 12480 16091 12544
rect 15770 11456 16091 12480
rect 15770 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15938 11456
rect 16002 11392 16018 11456
rect 16082 11392 16091 11456
rect 15147 11116 15213 11117
rect 15147 11052 15148 11116
rect 15212 11052 15213 11116
rect 15147 11051 15213 11052
rect 12805 10848 12813 10912
rect 12877 10848 12893 10912
rect 12957 10848 12973 10912
rect 13037 10848 13053 10912
rect 13117 10848 13125 10912
rect 12805 9824 13125 10848
rect 12805 9760 12813 9824
rect 12877 9760 12893 9824
rect 12957 9760 12973 9824
rect 13037 9760 13053 9824
rect 13117 9760 13125 9824
rect 12805 8736 13125 9760
rect 12805 8672 12813 8736
rect 12877 8672 12893 8736
rect 12957 8672 12973 8736
rect 13037 8672 13053 8736
rect 13117 8672 13125 8736
rect 12805 7648 13125 8672
rect 14043 8532 14109 8533
rect 14043 8468 14044 8532
rect 14108 8468 14109 8532
rect 14043 8467 14109 8468
rect 12805 7584 12813 7648
rect 12877 7584 12893 7648
rect 12957 7584 12973 7648
rect 13037 7584 13053 7648
rect 13117 7584 13125 7648
rect 12387 7036 12453 7037
rect 12387 6972 12388 7036
rect 12452 6972 12453 7036
rect 12387 6971 12453 6972
rect 12390 6493 12450 6971
rect 12805 6560 13125 7584
rect 12805 6496 12813 6560
rect 12877 6496 12893 6560
rect 12957 6496 12973 6560
rect 13037 6496 13053 6560
rect 13117 6496 13125 6560
rect 12387 6492 12453 6493
rect 12387 6428 12388 6492
rect 12452 6428 12453 6492
rect 12387 6427 12453 6428
rect 9840 5952 9848 6016
rect 9912 5952 9928 6016
rect 9992 5952 10008 6016
rect 10072 5952 10088 6016
rect 10152 5952 10160 6016
rect 9840 4928 10160 5952
rect 9840 4864 9848 4928
rect 9912 4864 9928 4928
rect 9992 4864 10008 4928
rect 10072 4864 10088 4928
rect 10152 4864 10160 4928
rect 9840 3840 10160 4864
rect 9840 3776 9848 3840
rect 9912 3776 9928 3840
rect 9992 3776 10008 3840
rect 10072 3776 10088 3840
rect 10152 3776 10160 3840
rect 9840 2752 10160 3776
rect 9840 2688 9848 2752
rect 9912 2688 9928 2752
rect 9992 2688 10008 2752
rect 10072 2688 10088 2752
rect 10152 2688 10160 2752
rect 9840 2128 10160 2688
rect 12805 5472 13125 6496
rect 14046 5541 14106 8467
rect 15150 6629 15210 11051
rect 15770 10368 16091 11392
rect 15770 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15938 10368
rect 16002 10304 16018 10368
rect 16082 10304 16091 10368
rect 15770 9280 16091 10304
rect 15770 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15938 9280
rect 16002 9216 16018 9280
rect 16082 9216 16091 9280
rect 15770 8192 16091 9216
rect 15770 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15938 8192
rect 16002 8128 16018 8192
rect 16082 8128 16091 8192
rect 15770 7104 16091 8128
rect 15770 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15938 7104
rect 16002 7040 16018 7104
rect 16082 7040 16091 7104
rect 15147 6628 15213 6629
rect 15147 6564 15148 6628
rect 15212 6564 15213 6628
rect 15147 6563 15213 6564
rect 15770 6016 16091 7040
rect 15770 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15938 6016
rect 16002 5952 16018 6016
rect 16082 5952 16091 6016
rect 14043 5540 14109 5541
rect 14043 5476 14044 5540
rect 14108 5476 14109 5540
rect 14043 5475 14109 5476
rect 12805 5408 12813 5472
rect 12877 5408 12893 5472
rect 12957 5408 12973 5472
rect 13037 5408 13053 5472
rect 13117 5408 13125 5472
rect 12805 4384 13125 5408
rect 12805 4320 12813 4384
rect 12877 4320 12893 4384
rect 12957 4320 12973 4384
rect 13037 4320 13053 4384
rect 13117 4320 13125 4384
rect 12805 3296 13125 4320
rect 12805 3232 12813 3296
rect 12877 3232 12893 3296
rect 12957 3232 12973 3296
rect 13037 3232 13053 3296
rect 13117 3232 13125 3296
rect 12805 2208 13125 3232
rect 12805 2144 12813 2208
rect 12877 2144 12893 2208
rect 12957 2144 12973 2208
rect 13037 2144 13053 2208
rect 13117 2144 13125 2208
rect 12805 2128 13125 2144
rect 15770 4928 16091 5952
rect 15770 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15938 4928
rect 16002 4864 16018 4928
rect 16082 4864 16091 4928
rect 15770 3840 16091 4864
rect 15770 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15938 3840
rect 16002 3776 16018 3840
rect 16082 3776 16091 3840
rect 15770 2752 16091 3776
rect 15770 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15938 2752
rect 16002 2688 16018 2752
rect 16082 2688 16091 2752
rect 15770 2128 16091 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__329__B pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13064 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1644511149
transform -1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1644511149
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A
timestamp 1644511149
transform 1 0 15824 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__A
timestamp 1644511149
transform 1 0 14260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clock_A
timestamp 1644511149
transform -1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 6256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 12972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 14076 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 14536 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 10120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 2024 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 16008 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 15456 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 2760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 17940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 16744 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 3956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 2392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 17572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1644511149
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1644511149
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1644511149
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1644511149
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72
timestamp 1644511149
transform 1 0 7728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1644511149
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_93
timestamp 1644511149
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_104
timestamp 1644511149
transform 1 0 10672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1644511149
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_123
timestamp 1644511149
transform 1 0 12420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1644511149
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132
timestamp 1644511149
transform 1 0 13248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1644511149
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_159
timestamp 1644511149
transform 1 0 15732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1644511149
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_188
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_20
timestamp 1644511149
transform 1 0 2944 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_25
timestamp 1644511149
transform 1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_47
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1644511149
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp 1644511149
transform 1 0 7820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_78
timestamp 1644511149
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_97
timestamp 1644511149
transform 1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_102
timestamp 1644511149
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1644511149
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_130
timestamp 1644511149
transform 1 0 13064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1644511149
transform 1 0 14168 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1644511149
transform 1 0 14536 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_185
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1644511149
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_8
timestamp 1644511149
transform 1 0 1840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1644511149
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1644511149
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1644511149
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1644511149
transform 1 0 6256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_60
timestamp 1644511149
transform 1 0 6624 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1644511149
transform 1 0 7176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_70 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1644511149
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1644511149
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_98
timestamp 1644511149
transform 1 0 10120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_116
timestamp 1644511149
transform 1 0 11776 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1644511149
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_127
timestamp 1644511149
transform 1 0 12788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_131
timestamp 1644511149
transform 1 0 13156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1644511149
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_150
timestamp 1644511149
transform 1 0 14904 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_155
timestamp 1644511149
transform 1 0 15364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_162
timestamp 1644511149
transform 1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_169
timestamp 1644511149
transform 1 0 16652 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_176
timestamp 1644511149
transform 1 0 17296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_180
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_14
timestamp 1644511149
transform 1 0 2392 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp 1644511149
transform 1 0 2760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_29
timestamp 1644511149
transform 1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 1644511149
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1644511149
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1644511149
transform 1 0 7544 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_88
timestamp 1644511149
transform 1 0 9200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_96
timestamp 1644511149
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1644511149
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_119
timestamp 1644511149
transform 1 0 12052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_124
timestamp 1644511149
transform 1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_129
timestamp 1644511149
transform 1 0 12972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_134
timestamp 1644511149
transform 1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_141
timestamp 1644511149
transform 1 0 14076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_146
timestamp 1644511149
transform 1 0 14536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1644511149
transform 1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 1644511149
transform 1 0 15640 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1644511149
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_182
timestamp 1644511149
transform 1 0 17848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1644511149
transform 1 0 18400 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1644511149
transform 1 0 3128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1644511149
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_33
timestamp 1644511149
transform 1 0 4140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_39
timestamp 1644511149
transform 1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_46
timestamp 1644511149
transform 1 0 5336 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_55
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_59 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1644511149
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9660 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_115
timestamp 1644511149
transform 1 0 11684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_125
timestamp 1644511149
transform 1 0 12604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1644511149
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1644511149
transform 1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_162
timestamp 1644511149
transform 1 0 16008 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_169
timestamp 1644511149
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1644511149
transform 1 0 18400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_5
timestamp 1644511149
transform 1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_12
timestamp 1644511149
transform 1 0 2208 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1644511149
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_43
timestamp 1644511149
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_47
timestamp 1644511149
transform 1 0 5428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1644511149
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1644511149
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_71
timestamp 1644511149
transform 1 0 7636 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_95
timestamp 1644511149
transform 1 0 9844 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1644511149
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1644511149
transform 1 0 11960 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_136
timestamp 1644511149
transform 1 0 13616 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_142
timestamp 1644511149
transform 1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_153
timestamp 1644511149
transform 1 0 15180 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1644511149
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_185
timestamp 1644511149
transform 1 0 18124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1644511149
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1644511149
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_39
timestamp 1644511149
transform 1 0 4692 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_61
timestamp 1644511149
transform 1 0 6716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1644511149
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_92
timestamp 1644511149
transform 1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp 1644511149
transform 1 0 10396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1644511149
transform 1 0 11224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_119
timestamp 1644511149
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_126
timestamp 1644511149
transform 1 0 12696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_130
timestamp 1644511149
transform 1 0 13064 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1644511149
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_145
timestamp 1644511149
transform 1 0 14444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_164
timestamp 1644511149
transform 1 0 16192 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_175
timestamp 1644511149
transform 1 0 17204 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_188
timestamp 1644511149
transform 1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_13
timestamp 1644511149
transform 1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp 1644511149
transform 1 0 3312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1644511149
transform 1 0 3956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_42
timestamp 1644511149
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_48
timestamp 1644511149
transform 1 0 5520 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1644511149
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_64
timestamp 1644511149
transform 1 0 6992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1644511149
transform 1 0 7636 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_83
timestamp 1644511149
transform 1 0 8740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_94
timestamp 1644511149
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_103
timestamp 1644511149
transform 1 0 10580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1644511149
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1644511149
transform 1 0 12144 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_126
timestamp 1644511149
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1644511149
transform 1 0 13524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_144
timestamp 1644511149
transform 1 0 14352 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_153
timestamp 1644511149
transform 1 0 15180 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_159
timestamp 1644511149
transform 1 0 15732 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1644511149
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_187
timestamp 1644511149
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_6
timestamp 1644511149
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_14
timestamp 1644511149
transform 1 0 2392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1644511149
transform 1 0 2852 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1644511149
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1644511149
transform 1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_60
timestamp 1644511149
transform 1 0 6624 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 1644511149
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1644511149
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1644511149
transform 1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_108
timestamp 1644511149
transform 1 0 11040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_119
timestamp 1644511149
transform 1 0 12052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1644511149
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1644511149
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_148
timestamp 1644511149
transform 1 0 14720 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_157
timestamp 1644511149
transform 1 0 15548 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1644511149
transform 1 0 16100 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_174
timestamp 1644511149
transform 1 0 17112 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_185
timestamp 1644511149
transform 1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_22
timestamp 1644511149
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_26
timestamp 1644511149
transform 1 0 3496 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1644511149
transform 1 0 4508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_44
timestamp 1644511149
transform 1 0 5152 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1644511149
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_64
timestamp 1644511149
transform 1 0 6992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1644511149
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1644511149
transform 1 0 8280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_90
timestamp 1644511149
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_95
timestamp 1644511149
transform 1 0 9844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_101
timestamp 1644511149
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1644511149
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1644511149
transform 1 0 12420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 1644511149
transform 1 0 12972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_140
timestamp 1644511149
transform 1 0 13984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_150
timestamp 1644511149
transform 1 0 14904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_159
timestamp 1644511149
transform 1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1644511149
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1644511149
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_12
timestamp 1644511149
transform 1 0 2208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1644511149
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1644511149
transform 1 0 4692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_51
timestamp 1644511149
transform 1 0 5796 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_56
timestamp 1644511149
transform 1 0 6256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_63
timestamp 1644511149
transform 1 0 6900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_67
timestamp 1644511149
transform 1 0 7268 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_95
timestamp 1644511149
transform 1 0 9844 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_108
timestamp 1644511149
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_114
timestamp 1644511149
transform 1 0 11592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_123
timestamp 1644511149
transform 1 0 12420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_132
timestamp 1644511149
transform 1 0 13248 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1644511149
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1644511149
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_155
timestamp 1644511149
transform 1 0 15364 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_159
timestamp 1644511149
transform 1 0 15732 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_163
timestamp 1644511149
transform 1 0 16100 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_174
timestamp 1644511149
transform 1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1644511149
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_12
timestamp 1644511149
transform 1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1644511149
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_28
timestamp 1644511149
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_45
timestamp 1644511149
transform 1 0 5244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_73
timestamp 1644511149
transform 1 0 7820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp 1644511149
transform 1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_91
timestamp 1644511149
transform 1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1644511149
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_117
timestamp 1644511149
transform 1 0 11868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_127
timestamp 1644511149
transform 1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_148
timestamp 1644511149
transform 1 0 14720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1644511149
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_186
timestamp 1644511149
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_21
timestamp 1644511149
transform 1 0 3036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1644511149
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_47
timestamp 1644511149
transform 1 0 5428 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_57
timestamp 1644511149
transform 1 0 6348 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp 1644511149
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_67
timestamp 1644511149
transform 1 0 7268 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1644511149
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1644511149
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_117
timestamp 1644511149
transform 1 0 11868 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_122
timestamp 1644511149
transform 1 0 12328 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_126
timestamp 1644511149
transform 1 0 12696 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_134
timestamp 1644511149
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1644511149
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_150
timestamp 1644511149
transform 1 0 14904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_154
timestamp 1644511149
transform 1 0 15272 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_158
timestamp 1644511149
transform 1 0 15640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_162
timestamp 1644511149
transform 1 0 16008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_169
timestamp 1644511149
transform 1 0 16652 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_174
timestamp 1644511149
transform 1 0 17112 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_179
timestamp 1644511149
transform 1 0 17572 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1644511149
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1644511149
transform 1 0 2576 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_21
timestamp 1644511149
transform 1 0 3036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1644511149
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_36
timestamp 1644511149
transform 1 0 4416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1644511149
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_61
timestamp 1644511149
transform 1 0 6716 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_87
timestamp 1644511149
transform 1 0 9108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1644511149
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1644511149
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_134
timestamp 1644511149
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_141
timestamp 1644511149
transform 1 0 14076 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_145
timestamp 1644511149
transform 1 0 14444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1644511149
transform 1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_160
timestamp 1644511149
transform 1 0 15824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1644511149
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_174
timestamp 1644511149
transform 1 0 17112 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_182
timestamp 1644511149
transform 1 0 17848 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1644511149
transform 1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_6
timestamp 1644511149
transform 1 0 1656 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_10
timestamp 1644511149
transform 1 0 2024 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_14
timestamp 1644511149
transform 1 0 2392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1644511149
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_35
timestamp 1644511149
transform 1 0 4324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_40
timestamp 1644511149
transform 1 0 4784 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_44
timestamp 1644511149
transform 1 0 5152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_49
timestamp 1644511149
transform 1 0 5612 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_54
timestamp 1644511149
transform 1 0 6072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1644511149
transform 1 0 7728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1644511149
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1644511149
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_103
timestamp 1644511149
transform 1 0 10580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_119
timestamp 1644511149
transform 1 0 12052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1644511149
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_157
timestamp 1644511149
transform 1 0 15548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1644511149
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1644511149
transform 1 0 18400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_23
timestamp 1644511149
transform 1 0 3220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_29
timestamp 1644511149
transform 1 0 3772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_46
timestamp 1644511149
transform 1 0 5336 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1644511149
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_65
timestamp 1644511149
transform 1 0 7084 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1644511149
transform 1 0 7636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_76
timestamp 1644511149
transform 1 0 8096 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_88
timestamp 1644511149
transform 1 0 9200 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_98
timestamp 1644511149
transform 1 0 10120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_104
timestamp 1644511149
transform 1 0 10672 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1644511149
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_121
timestamp 1644511149
transform 1 0 12236 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1644511149
transform 1 0 13524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1644511149
transform 1 0 14076 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1644511149
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1644511149
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_185
timestamp 1644511149
transform 1 0 18124 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1644511149
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_6
timestamp 1644511149
transform 1 0 1656 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_17
timestamp 1644511149
transform 1 0 2668 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1644511149
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_34
timestamp 1644511149
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_40
timestamp 1644511149
transform 1 0 4784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1644511149
transform 1 0 5336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_51
timestamp 1644511149
transform 1 0 5796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1644511149
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_74
timestamp 1644511149
transform 1 0 7912 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_78
timestamp 1644511149
transform 1 0 8280 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1644511149
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1644511149
transform 1 0 9384 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_101
timestamp 1644511149
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_108
timestamp 1644511149
transform 1 0 11040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_114
timestamp 1644511149
transform 1 0 11592 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1644511149
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1644511149
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1644511149
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_155
timestamp 1644511149
transform 1 0 15364 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_161
timestamp 1644511149
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_172
timestamp 1644511149
transform 1 0 16928 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_176
timestamp 1644511149
transform 1 0 17296 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_179
timestamp 1644511149
transform 1 0 17572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_183
timestamp 1644511149
transform 1 0 17940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp 1644511149
transform 1 0 18400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_6
timestamp 1644511149
transform 1 0 1656 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_24
timestamp 1644511149
transform 1 0 3312 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_28
timestamp 1644511149
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_45
timestamp 1644511149
transform 1 0 5244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1644511149
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_65
timestamp 1644511149
transform 1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1644511149
transform 1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_102
timestamp 1644511149
transform 1 0 10488 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1644511149
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_129
timestamp 1644511149
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1644511149
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_156
timestamp 1644511149
transform 1 0 15456 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1644511149
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_186
timestamp 1644511149
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1644511149
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_38
timestamp 1644511149
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_45
timestamp 1644511149
transform 1 0 5244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_54
timestamp 1644511149
transform 1 0 6072 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_59
timestamp 1644511149
transform 1 0 6532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_67
timestamp 1644511149
transform 1 0 7268 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_73
timestamp 1644511149
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1644511149
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_95
timestamp 1644511149
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_104
timestamp 1644511149
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_111
timestamp 1644511149
transform 1 0 11316 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_118
timestamp 1644511149
transform 1 0 11960 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1644511149
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1644511149
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1644511149
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_156
timestamp 1644511149
transform 1 0 15456 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1644511149
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1644511149
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1644511149
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_13
timestamp 1644511149
transform 1 0 2300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_24
timestamp 1644511149
transform 1 0 3312 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1644511149
transform 1 0 4048 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_38
timestamp 1644511149
transform 1 0 4600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_45
timestamp 1644511149
transform 1 0 5244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1644511149
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_60
timestamp 1644511149
transform 1 0 6624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1644511149
transform 1 0 8280 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_90
timestamp 1644511149
transform 1 0 9384 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1644511149
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1644511149
transform 1 0 10304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1644511149
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1644511149
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_135
timestamp 1644511149
transform 1 0 13524 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_143
timestamp 1644511149
transform 1 0 14260 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_154
timestamp 1644511149
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1644511149
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_178
timestamp 1644511149
transform 1 0 17480 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_188
timestamp 1644511149
transform 1 0 18400 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1644511149
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1644511149
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1644511149
transform 1 0 4048 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_37
timestamp 1644511149
transform 1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_42
timestamp 1644511149
transform 1 0 4968 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1644511149
transform 1 0 5520 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_55
timestamp 1644511149
transform 1 0 6164 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1644511149
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_67
timestamp 1644511149
transform 1 0 7268 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_88
timestamp 1644511149
transform 1 0 9200 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_94
timestamp 1644511149
transform 1 0 9752 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_111
timestamp 1644511149
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1644511149
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1644511149
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_147
timestamp 1644511149
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_158
timestamp 1644511149
transform 1 0 15640 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_170
timestamp 1644511149
transform 1 0 16744 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_188
timestamp 1644511149
transform 1 0 18400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_23
timestamp 1644511149
transform 1 0 3220 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_40
timestamp 1644511149
transform 1 0 4784 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_44
timestamp 1644511149
transform 1 0 5152 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1644511149
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_63
timestamp 1644511149
transform 1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_74
timestamp 1644511149
transform 1 0 7912 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_87
timestamp 1644511149
transform 1 0 9108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_94
timestamp 1644511149
transform 1 0 9752 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1644511149
transform 1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_103
timestamp 1644511149
transform 1 0 10580 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1644511149
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_124
timestamp 1644511149
transform 1 0 12512 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_142
timestamp 1644511149
transform 1 0 14168 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1644511149
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1644511149
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_6
timestamp 1644511149
transform 1 0 1656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp 1644511149
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1644511149
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_35
timestamp 1644511149
transform 1 0 4324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_50
timestamp 1644511149
transform 1 0 5704 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1644511149
transform 1 0 6532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_74
timestamp 1644511149
transform 1 0 7912 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1644511149
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1644511149
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_100
timestamp 1644511149
transform 1 0 10304 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_106
timestamp 1644511149
transform 1 0 10856 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1644511149
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_117
timestamp 1644511149
transform 1 0 11868 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_125
timestamp 1644511149
transform 1 0 12604 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1644511149
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_150
timestamp 1644511149
transform 1 0 14904 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_155
timestamp 1644511149
transform 1 0 15364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_160
timestamp 1644511149
transform 1 0 15824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_166
timestamp 1644511149
transform 1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_170
timestamp 1644511149
transform 1 0 16744 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_178
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1644511149
transform 1 0 17940 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_6
timestamp 1644511149
transform 1 0 1656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_24
timestamp 1644511149
transform 1 0 3312 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_35
timestamp 1644511149
transform 1 0 4324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_43
timestamp 1644511149
transform 1 0 5060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_64
timestamp 1644511149
transform 1 0 6992 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_75
timestamp 1644511149
transform 1 0 8004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_79
timestamp 1644511149
transform 1 0 8372 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_88
timestamp 1644511149
transform 1 0 9200 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_100
timestamp 1644511149
transform 1 0 10304 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1644511149
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1644511149
transform 1 0 12144 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1644511149
transform 1 0 12788 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_147
timestamp 1644511149
transform 1 0 14628 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1644511149
transform 1 0 15456 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1644511149
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_174
timestamp 1644511149
transform 1 0 17112 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_179
timestamp 1644511149
transform 1 0 17572 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_188
timestamp 1644511149
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_20
timestamp 1644511149
transform 1 0 2944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1644511149
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_39
timestamp 1644511149
transform 1 0 4692 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_61
timestamp 1644511149
transform 1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_69
timestamp 1644511149
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1644511149
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_95
timestamp 1644511149
transform 1 0 9844 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1644511149
transform 1 0 10488 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_111
timestamp 1644511149
transform 1 0 11316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1644511149
transform 1 0 12420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_132
timestamp 1644511149
transform 1 0 13248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1644511149
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1644511149
transform 1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1644511149
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1644511149
transform 1 0 16560 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_188
timestamp 1644511149
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_6
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_10
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_14
timestamp 1644511149
transform 1 0 2392 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_22
timestamp 1644511149
transform 1 0 3128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_31
timestamp 1644511149
transform 1 0 3956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_43
timestamp 1644511149
transform 1 0 5060 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1644511149
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_64
timestamp 1644511149
transform 1 0 6992 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_88
timestamp 1644511149
transform 1 0 9200 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1644511149
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1644511149
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1644511149
transform 1 0 12420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1644511149
transform 1 0 13248 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_139
timestamp 1644511149
transform 1 0 13892 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_150
timestamp 1644511149
transform 1 0 14904 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1644511149
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_174
timestamp 1644511149
transform 1 0 17112 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1644511149
transform 1 0 17572 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_184
timestamp 1644511149
transform 1 0 18032 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_9
timestamp 1644511149
transform 1 0 1932 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_19
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1644511149
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_45
timestamp 1644511149
transform 1 0 5244 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_50
timestamp 1644511149
transform 1 0 5704 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_69
timestamp 1644511149
transform 1 0 7452 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1644511149
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_103
timestamp 1644511149
transform 1 0 10580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_107
timestamp 1644511149
transform 1 0 10948 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1644511149
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1644511149
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1644511149
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_159
timestamp 1644511149
transform 1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_166
timestamp 1644511149
transform 1 0 16376 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_184
timestamp 1644511149
transform 1 0 18032 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_13
timestamp 1644511149
transform 1 0 2300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_18
timestamp 1644511149
transform 1 0 2760 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_23
timestamp 1644511149
transform 1 0 3220 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_31
timestamp 1644511149
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_43
timestamp 1644511149
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_63
timestamp 1644511149
transform 1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_77
timestamp 1644511149
transform 1 0 8188 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1644511149
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_97
timestamp 1644511149
transform 1 0 10028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_103
timestamp 1644511149
transform 1 0 10580 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1644511149
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_124
timestamp 1644511149
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_129
timestamp 1644511149
transform 1 0 12972 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_134
timestamp 1644511149
transform 1 0 13432 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1644511149
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_147
timestamp 1644511149
transform 1 0 14628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_152
timestamp 1644511149
transform 1 0 15088 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_156
timestamp 1644511149
transform 1 0 15456 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1644511149
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_172
timestamp 1644511149
transform 1 0 16928 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_182
timestamp 1644511149
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_188
timestamp 1644511149
transform 1 0 18400 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _315_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1644511149
transform -1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _317_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _318_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9568 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _319_
timestamp 1644511149
transform 1 0 14628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _320_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13984 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _321_
timestamp 1644511149
transform 1 0 12880 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _322_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13800 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _323_
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _324_
timestamp 1644511149
transform 1 0 8464 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _325_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _326_
timestamp 1644511149
transform 1 0 10856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _327_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18216 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _328_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16192 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _329_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _330_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9936 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_2  _331_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7820 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _332_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _333_
timestamp 1644511149
transform 1 0 12328 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _334_
timestamp 1644511149
transform 1 0 7728 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _335_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9752 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _336_
timestamp 1644511149
transform 1 0 12788 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _337_
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _338_
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _339_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9844 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _340_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7176 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _341_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _342_
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _343_
timestamp 1644511149
transform -1 0 12420 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _344_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 13248 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _345_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9108 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _346_
timestamp 1644511149
transform 1 0 13800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _347_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12788 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _348_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17296 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _349_
timestamp 1644511149
transform -1 0 18216 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _350_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _351_
timestamp 1644511149
transform -1 0 13708 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _352_
timestamp 1644511149
transform 1 0 17296 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _353_
timestamp 1644511149
transform 1 0 9752 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _354_
timestamp 1644511149
transform 1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _355_
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _356_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 11224 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _357_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14352 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _358_
timestamp 1644511149
transform -1 0 15824 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _359_
timestamp 1644511149
transform 1 0 15088 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _360_
timestamp 1644511149
transform 1 0 14904 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _361_
timestamp 1644511149
transform -1 0 14904 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _362_
timestamp 1644511149
transform 1 0 14628 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _363_
timestamp 1644511149
transform -1 0 17296 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _364_
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _365_
timestamp 1644511149
transform -1 0 15180 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _366_
timestamp 1644511149
transform -1 0 16100 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _367_
timestamp 1644511149
transform -1 0 16376 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _368_
timestamp 1644511149
transform -1 0 11960 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _369_
timestamp 1644511149
transform 1 0 11408 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _370_
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _371_
timestamp 1644511149
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _372_
timestamp 1644511149
transform -1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _373_
timestamp 1644511149
transform 1 0 5520 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _374_
timestamp 1644511149
transform 1 0 11224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _375_
timestamp 1644511149
transform 1 0 10120 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _376_
timestamp 1644511149
transform 1 0 12788 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _377_
timestamp 1644511149
transform -1 0 12052 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _378_
timestamp 1644511149
transform 1 0 13892 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _379_
timestamp 1644511149
transform -1 0 12420 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _380_
timestamp 1644511149
transform 1 0 10396 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _381_
timestamp 1644511149
transform 1 0 10488 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _382_
timestamp 1644511149
transform -1 0 11132 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _383_
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _384_
timestamp 1644511149
transform -1 0 8280 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_2  _385_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4968 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _386_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _387_
timestamp 1644511149
transform 1 0 3680 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _388_
timestamp 1644511149
transform -1 0 10488 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _389_
timestamp 1644511149
transform -1 0 9844 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _390_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _391_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7636 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _392_
timestamp 1644511149
transform -1 0 8004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _393_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 5796 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _394_
timestamp 1644511149
transform 1 0 9384 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _395_
timestamp 1644511149
transform -1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _396_
timestamp 1644511149
transform 1 0 15088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _397_
timestamp 1644511149
transform 1 0 14260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _398_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _399_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _400_
timestamp 1644511149
transform -1 0 4968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _401_
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _402_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 6072 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _403_
timestamp 1644511149
transform -1 0 9384 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _404_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10212 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _405_
timestamp 1644511149
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _406_
timestamp 1644511149
transform -1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _407_
timestamp 1644511149
transform 1 0 10212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _408_
timestamp 1644511149
transform 1 0 9108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1644511149
transform -1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _410_
timestamp 1644511149
transform -1 0 5428 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1644511149
transform 1 0 4048 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _412_
timestamp 1644511149
transform 1 0 3956 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _413_
timestamp 1644511149
transform 1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1644511149
transform -1 0 4692 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _415_
timestamp 1644511149
transform -1 0 5888 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _416_
timestamp 1644511149
transform -1 0 3496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp 1644511149
transform -1 0 4968 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _418_
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _419_
timestamp 1644511149
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _420_
timestamp 1644511149
transform 1 0 4140 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _421_
timestamp 1644511149
transform 1 0 3036 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _422_
timestamp 1644511149
transform -1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _423_
timestamp 1644511149
transform 1 0 3864 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _424_
timestamp 1644511149
transform 1 0 3496 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _425_
timestamp 1644511149
transform 1 0 3864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _426_
timestamp 1644511149
transform -1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _427_
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _428_
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _429_
timestamp 1644511149
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _430_
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _431_
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _432_
timestamp 1644511149
transform -1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _433_
timestamp 1644511149
transform 1 0 6716 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _434_
timestamp 1644511149
transform 1 0 6716 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _435_
timestamp 1644511149
transform 1 0 7360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _436_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _437_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _438_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8188 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _439_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 11868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _440_
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _441_
timestamp 1644511149
transform -1 0 14076 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _442_
timestamp 1644511149
transform -1 0 13432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _444_
timestamp 1644511149
transform 1 0 16192 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _445_
timestamp 1644511149
transform -1 0 17112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _446_
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _447_
timestamp 1644511149
transform 1 0 13340 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _448_
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _449_
timestamp 1644511149
transform -1 0 16744 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _450_
timestamp 1644511149
transform -1 0 17112 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _451_
timestamp 1644511149
transform -1 0 16376 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _452_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _453_
timestamp 1644511149
transform -1 0 13800 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _454_
timestamp 1644511149
transform -1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _455_
timestamp 1644511149
transform 1 0 11592 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _456_
timestamp 1644511149
transform -1 0 11224 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _457_
timestamp 1644511149
transform -1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _458_
timestamp 1644511149
transform 1 0 4416 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _459_
timestamp 1644511149
transform 1 0 12144 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _460_
timestamp 1644511149
transform 1 0 10672 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _461_
timestamp 1644511149
transform -1 0 11040 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1644511149
transform 1 0 9568 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _463_
timestamp 1644511149
transform -1 0 9384 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _464_
timestamp 1644511149
transform -1 0 8648 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _465_
timestamp 1644511149
transform -1 0 9384 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _466_
timestamp 1644511149
transform 1 0 7360 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _467_
timestamp 1644511149
transform -1 0 6900 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _468_
timestamp 1644511149
transform -1 0 6348 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1644511149
transform -1 0 7452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _470_
timestamp 1644511149
transform 1 0 6716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _471_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7912 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _472_
timestamp 1644511149
transform -1 0 4324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _473_
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _474_
timestamp 1644511149
transform -1 0 2668 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _475_
timestamp 1644511149
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _476_
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _477_
timestamp 1644511149
transform 1 0 2116 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _478_
timestamp 1644511149
transform 1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _479_
timestamp 1644511149
transform -1 0 4508 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _480_
timestamp 1644511149
transform 1 0 2392 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _481_
timestamp 1644511149
transform -1 0 2392 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _482_
timestamp 1644511149
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _483_
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _484_
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _485_
timestamp 1644511149
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _486_
timestamp 1644511149
transform 1 0 2392 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _487_
timestamp 1644511149
transform -1 0 2392 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _488_
timestamp 1644511149
transform -1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _489_
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _490_
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _491_
timestamp 1644511149
transform 1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _492_
timestamp 1644511149
transform 1 0 3864 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _493_
timestamp 1644511149
transform 1 0 3956 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _494_
timestamp 1644511149
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _495_
timestamp 1644511149
transform -1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _496_
timestamp 1644511149
transform 1 0 6532 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _497_
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _498_
timestamp 1644511149
transform 1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _499_
timestamp 1644511149
transform 1 0 13248 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _500_
timestamp 1644511149
transform -1 0 13524 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _501_
timestamp 1644511149
transform 1 0 16100 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _502_
timestamp 1644511149
transform 1 0 14996 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _503_
timestamp 1644511149
transform 1 0 12144 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _504_
timestamp 1644511149
transform -1 0 16376 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _505_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _506_
timestamp 1644511149
transform 1 0 15456 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _507_
timestamp 1644511149
transform -1 0 16744 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _508_
timestamp 1644511149
transform 1 0 15916 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _509_
timestamp 1644511149
transform 1 0 14996 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _510_
timestamp 1644511149
transform -1 0 16376 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _511_
timestamp 1644511149
transform 1 0 14812 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _512_
timestamp 1644511149
transform 1 0 14352 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _513_
timestamp 1644511149
transform -1 0 15272 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _514_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _515_
timestamp 1644511149
transform 1 0 11500 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _516_
timestamp 1644511149
transform -1 0 13432 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _517_
timestamp 1644511149
transform 1 0 12696 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _518_
timestamp 1644511149
transform 1 0 10856 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _519_
timestamp 1644511149
transform 1 0 11776 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _520_
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _521_
timestamp 1644511149
transform 1 0 7820 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _522_
timestamp 1644511149
transform 1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _523_
timestamp 1644511149
transform 1 0 16376 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _524_
timestamp 1644511149
transform 1 0 16192 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1644511149
transform -1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _526_
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _527_
timestamp 1644511149
transform -1 0 16376 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _528_
timestamp 1644511149
transform -1 0 16100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _529_
timestamp 1644511149
transform 1 0 17296 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _530_
timestamp 1644511149
transform -1 0 16376 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _531_
timestamp 1644511149
transform -1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _532_
timestamp 1644511149
transform -1 0 13800 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _533_
timestamp 1644511149
transform 1 0 13616 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _534_
timestamp 1644511149
transform -1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _535_
timestamp 1644511149
transform -1 0 12604 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _536_
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _537_
timestamp 1644511149
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _538_
timestamp 1644511149
transform 1 0 9292 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _539_
timestamp 1644511149
transform 1 0 9568 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _540_
timestamp 1644511149
transform 1 0 10396 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _541_
timestamp 1644511149
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _542_
timestamp 1644511149
transform 1 0 8832 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _543_
timestamp 1644511149
transform 1 0 7912 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _544_
timestamp 1644511149
transform 1 0 7820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _545_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5244 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _546_
timestamp 1644511149
transform -1 0 9200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _547_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 11868 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _548_
timestamp 1644511149
transform -1 0 12236 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _549_
timestamp 1644511149
transform -1 0 12328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _550_
timestamp 1644511149
transform 1 0 6808 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _551_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12052 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _552_
timestamp 1644511149
transform -1 0 5336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _553_
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1644511149
transform -1 0 3496 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _555_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5704 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _556_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _557_
timestamp 1644511149
transform 1 0 10580 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _558_
timestamp 1644511149
transform 1 0 5888 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _559_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _560_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14996 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _561_
timestamp 1644511149
transform -1 0 11868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _562_
timestamp 1644511149
transform -1 0 12144 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _563_
timestamp 1644511149
transform -1 0 11316 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _564_
timestamp 1644511149
transform 1 0 9844 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _565_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 10948 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _566_
timestamp 1644511149
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _567_
timestamp 1644511149
transform 1 0 15640 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _568_
timestamp 1644511149
transform -1 0 13248 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _569_
timestamp 1644511149
transform -1 0 10212 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _570_
timestamp 1644511149
transform 1 0 9292 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _571_
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _572_
timestamp 1644511149
transform -1 0 9200 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _573_
timestamp 1644511149
transform -1 0 11408 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _574_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11040 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _575_
timestamp 1644511149
transform -1 0 12512 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _576_
timestamp 1644511149
transform -1 0 12144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _577_
timestamp 1644511149
transform -1 0 13892 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _578_
timestamp 1644511149
transform 1 0 9844 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _579_
timestamp 1644511149
transform -1 0 11224 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _580_
timestamp 1644511149
transform 1 0 9384 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _581_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 12420 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _582_
timestamp 1644511149
transform 1 0 12328 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _583_
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _584_
timestamp 1644511149
transform 1 0 13432 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _585_
timestamp 1644511149
transform 1 0 16100 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _586_
timestamp 1644511149
transform 1 0 16100 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _587_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _588_
timestamp 1644511149
transform 1 0 17296 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _589_
timestamp 1644511149
transform 1 0 15456 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _590_
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _591_
timestamp 1644511149
transform 1 0 14260 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _592_
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _593_
timestamp 1644511149
transform 1 0 15916 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _594_
timestamp 1644511149
transform 1 0 17296 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _595_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _596_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _597_
timestamp 1644511149
transform 1 0 5428 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _598_
timestamp 1644511149
transform 1 0 5520 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _599_
timestamp 1644511149
transform -1 0 7636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _600_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _601_
timestamp 1644511149
transform 1 0 6716 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _602_
timestamp 1644511149
transform -1 0 5520 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _603_
timestamp 1644511149
transform 1 0 8464 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _604_
timestamp 1644511149
transform -1 0 8556 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _605_
timestamp 1644511149
transform 1 0 7820 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _606_
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _607_
timestamp 1644511149
transform 1 0 7268 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _608_
timestamp 1644511149
transform 1 0 6808 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _609_
timestamp 1644511149
transform -1 0 7268 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _610_
timestamp 1644511149
transform 1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _611_
timestamp 1644511149
transform 1 0 4140 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _612_
timestamp 1644511149
transform -1 0 6900 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _613_
timestamp 1644511149
transform -1 0 3496 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _614_
timestamp 1644511149
transform -1 0 2760 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _615_
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _616_
timestamp 1644511149
transform -1 0 3496 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _617_
timestamp 1644511149
transform 1 0 2760 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _618_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _619_
timestamp 1644511149
transform 1 0 4508 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _620_
timestamp 1644511149
transform 1 0 3312 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _621_
timestamp 1644511149
transform -1 0 5888 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _622_
timestamp 1644511149
transform -1 0 6992 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _623_
timestamp 1644511149
transform 1 0 5428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _624_
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _625_
timestamp 1644511149
transform -1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _626_
timestamp 1644511149
transform -1 0 5244 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _627_
timestamp 1644511149
transform 1 0 2024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _628_
timestamp 1644511149
transform -1 0 5244 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _629_
timestamp 1644511149
transform 1 0 3036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _630_
timestamp 1644511149
transform 1 0 4140 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _631_
timestamp 1644511149
transform 1 0 6256 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _632_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16928 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _633_
timestamp 1644511149
transform 1 0 16928 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _634_
timestamp 1644511149
transform 1 0 14720 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _635_
timestamp 1644511149
transform 1 0 14260 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _636_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _637_
timestamp 1644511149
transform 1 0 8372 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _638_
timestamp 1644511149
transform 1 0 14904 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _639_
timestamp 1644511149
transform -1 0 11776 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _640_
timestamp 1644511149
transform 1 0 7728 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _641_
timestamp 1644511149
transform 1 0 9844 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _642_
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _643_
timestamp 1644511149
transform -1 0 6072 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _644_
timestamp 1644511149
transform 1 0 3772 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _645_
timestamp 1644511149
transform 1 0 5244 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _646_
timestamp 1644511149
transform -1 0 6624 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _647_
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _648_
timestamp 1644511149
transform 1 0 4600 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _649_
timestamp 1644511149
transform 1 0 6900 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _650_
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _651_
timestamp 1644511149
transform -1 0 15548 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _652_
timestamp 1644511149
transform 1 0 16744 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _653_
timestamp 1644511149
transform 1 0 14720 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _654_
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _655_
timestamp 1644511149
transform 1 0 14260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _656_
timestamp 1644511149
transform -1 0 13064 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _657_
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _658_
timestamp 1644511149
transform 1 0 9016 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _659_
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _660_
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _661_
timestamp 1644511149
transform 1 0 1564 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _662_
timestamp 1644511149
transform 1 0 1656 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _663_
timestamp 1644511149
transform 1 0 1472 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _664_
timestamp 1644511149
transform 1 0 1656 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _665_
timestamp 1644511149
transform 1 0 2024 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _666_
timestamp 1644511149
transform 1 0 3956 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _667_
timestamp 1644511149
transform -1 0 7820 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _668_
timestamp 1644511149
transform 1 0 13156 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _669_
timestamp 1644511149
transform 1 0 16744 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _670_
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _671_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _672_
timestamp 1644511149
transform -1 0 16192 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _673_
timestamp 1644511149
transform 1 0 12696 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _674_
timestamp 1644511149
transform 1 0 11500 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _675_
timestamp 1644511149
transform 1 0 7728 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _676_
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _677_
timestamp 1644511149
transform 1 0 16928 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _678_
timestamp 1644511149
transform 1 0 16836 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _679_
timestamp 1644511149
transform -1 0 15640 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _680_
timestamp 1644511149
transform 1 0 12144 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _681_
timestamp 1644511149
transform -1 0 10580 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _682_
timestamp 1644511149
transform 1 0 7636 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _683_
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _684_
timestamp 1644511149
transform 1 0 6256 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _685_
timestamp 1644511149
transform -1 0 12972 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _686_
timestamp 1644511149
transform 1 0 3864 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _687_
timestamp 1644511149
transform 1 0 7360 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _688_
timestamp 1644511149
transform -1 0 11132 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _689_
timestamp 1644511149
transform 1 0 12328 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _690_
timestamp 1644511149
transform 1 0 9108 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _691_
timestamp 1644511149
transform 1 0 13156 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _692_
timestamp 1644511149
transform 1 0 16928 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _693_
timestamp 1644511149
transform 1 0 14260 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _694_
timestamp 1644511149
transform 1 0 16560 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _695_
timestamp 1644511149
transform -1 0 7452 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _696_
timestamp 1644511149
transform 1 0 3312 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _697_
timestamp 1644511149
transform -1 0 8280 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _698_
timestamp 1644511149
transform 1 0 2024 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _699_
timestamp 1644511149
transform -1 0 5244 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _700_
timestamp 1644511149
transform 1 0 1472 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _701_
timestamp 1644511149
transform 1 0 1840 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _702_
timestamp 1644511149
transform 1 0 5244 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _703_
timestamp 1644511149
transform -1 0 7452 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _704_
timestamp 1644511149
transform 1 0 16928 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _705_
timestamp 1644511149
transform 1 0 1656 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _706_
timestamp 1644511149
transform 1 0 1840 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _707_
timestamp 1644511149
transform 1 0 3772 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _708__35 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _709__36
timestamp 1644511149
transform 1 0 17572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _710__37
timestamp 1644511149
transform -1 0 18032 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _711__38
timestamp 1644511149
transform -1 0 11040 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _712__39
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _713__40
timestamp 1644511149
transform 1 0 15824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _714__41
timestamp 1644511149
transform 1 0 17296 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _715__42
timestamp 1644511149
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _716__43
timestamp 1644511149
transform 1 0 18124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _717__44
timestamp 1644511149
transform 1 0 15732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _718__45
timestamp 1644511149
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _719__46
timestamp 1644511149
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _720__47
timestamp 1644511149
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _721__48
timestamp 1644511149
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _722__49
timestamp 1644511149
transform 1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _723__50
timestamp 1644511149
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _724__51
timestamp 1644511149
transform -1 0 12972 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _725__52
timestamp 1644511149
transform -1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _726__53
timestamp 1644511149
transform 1 0 17664 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _727__54
timestamp 1644511149
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _728__55
timestamp 1644511149
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _729__56
timestamp 1644511149
transform -1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _730__57
timestamp 1644511149
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _731__58
timestamp 1644511149
transform -1 0 13432 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clock pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clock
timestamp 1644511149
transform -1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clock
timestamp 1644511149
transform 1 0 10856 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_clock
timestamp 1644511149
transform -1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_clock
timestamp 1644511149
transform -1 0 5980 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_clock
timestamp 1644511149
transform 1 0 13432 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_clock
timestamp 1644511149
transform 1 0 13156 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clock
timestamp 1644511149
transform -1 0 5520 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clock
timestamp 1644511149
transform 1 0 6624 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clock
timestamp 1644511149
transform -1 0 4600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clock
timestamp 1644511149
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clock
timestamp 1644511149
transform -1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clock
timestamp 1644511149
transform 1 0 14996 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clock
timestamp 1644511149
transform -1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clock
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform 1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1644511149
transform 1 0 9108 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1644511149
transform 1 0 17480 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1644511149
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1644511149
transform -1 0 6072 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform -1 0 13156 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 15364 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform -1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1644511149
transform 1 0 1564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 17480 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform -1 0 15916 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 18124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform -1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 15548 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1644511149
transform -1 0 2300 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform -1 0 18400 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1644511149
transform 1 0 18032 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1644511149
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1644511149
transform -1 0 8188 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1644511149
transform -1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1644511149
transform 1 0 18032 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1644511149
transform 1 0 18032 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1644511149
transform -1 0 16284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1644511149
transform -1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1644511149
transform -1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1644511149
transform -1 0 10580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1644511149
transform 1 0 17480 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1644511149
transform -1 0 11224 0 1 2176
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 1368 800 1488 6 clock
port 0 nsew signal input
rlabel metal2 s 18050 19200 18106 20000 6 io_spi_clk
port 1 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 io_spi_cs
port 2 nsew signal tristate
rlabel metal2 s 18050 0 18106 800 6 io_spi_intr
port 3 nsew signal tristate
rlabel metal2 s 7102 19200 7158 20000 6 io_spi_miso
port 4 nsew signal input
rlabel metal2 s 7746 19200 7802 20000 6 io_spi_mosi
port 5 nsew signal tristate
rlabel metal2 s 9034 19200 9090 20000 6 io_spi_select
port 6 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 io_wbs_ack_o
port 7 nsew signal tristate
rlabel metal3 s 19200 4088 20000 4208 6 io_wbs_data_o[0]
port 8 nsew signal tristate
rlabel metal2 s 17406 19200 17462 20000 6 io_wbs_data_o[10]
port 9 nsew signal tristate
rlabel metal2 s 10322 19200 10378 20000 6 io_wbs_data_o[11]
port 10 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 io_wbs_data_o[12]
port 11 nsew signal tristate
rlabel metal3 s 19200 6128 20000 6248 6 io_wbs_data_o[13]
port 12 nsew signal tristate
rlabel metal3 s 19200 8848 20000 8968 6 io_wbs_data_o[14]
port 13 nsew signal tristate
rlabel metal3 s 19200 17688 20000 17808 6 io_wbs_data_o[15]
port 14 nsew signal tristate
rlabel metal3 s 19200 15648 20000 15768 6 io_wbs_data_o[16]
port 15 nsew signal tristate
rlabel metal3 s 19200 2048 20000 2168 6 io_wbs_data_o[17]
port 16 nsew signal tristate
rlabel metal3 s 0 14288 800 14408 6 io_wbs_data_o[18]
port 17 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 io_wbs_data_o[19]
port 18 nsew signal tristate
rlabel metal3 s 19200 12928 20000 13048 6 io_wbs_data_o[1]
port 19 nsew signal tristate
rlabel metal3 s 0 14968 800 15088 6 io_wbs_data_o[20]
port 20 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 io_wbs_data_o[21]
port 21 nsew signal tristate
rlabel metal3 s 19200 14288 20000 14408 6 io_wbs_data_o[22]
port 22 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 io_wbs_data_o[23]
port 23 nsew signal tristate
rlabel metal2 s 12254 19200 12310 20000 6 io_wbs_data_o[24]
port 24 nsew signal tristate
rlabel metal2 s 18 19200 74 20000 6 io_wbs_data_o[25]
port 25 nsew signal tristate
rlabel metal3 s 19200 14968 20000 15088 6 io_wbs_data_o[26]
port 26 nsew signal tristate
rlabel metal3 s 0 9528 800 9648 6 io_wbs_data_o[27]
port 27 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 io_wbs_data_o[28]
port 28 nsew signal tristate
rlabel metal3 s 0 688 800 808 6 io_wbs_data_o[29]
port 29 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 io_wbs_data_o[2]
port 30 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 io_wbs_data_o[30]
port 31 nsew signal tristate
rlabel metal2 s 12898 19200 12954 20000 6 io_wbs_data_o[31]
port 32 nsew signal tristate
rlabel metal2 s 14186 19200 14242 20000 6 io_wbs_data_o[3]
port 33 nsew signal tristate
rlabel metal2 s 16762 0 16818 800 6 io_wbs_data_o[4]
port 34 nsew signal tristate
rlabel metal2 s 9678 19200 9734 20000 6 io_wbs_data_o[5]
port 35 nsew signal tristate
rlabel metal3 s 19200 17008 20000 17128 6 io_wbs_data_o[6]
port 36 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 io_wbs_data_o[7]
port 37 nsew signal tristate
rlabel metal3 s 0 10888 800 11008 6 io_wbs_data_o[8]
port 38 nsew signal tristate
rlabel metal3 s 19200 688 20000 808 6 io_wbs_data_o[9]
port 39 nsew signal tristate
rlabel metal3 s 19200 7488 20000 7608 6 io_wbs_m2s_addr[0]
port 40 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 io_wbs_m2s_addr[10]
port 41 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 io_wbs_m2s_addr[11]
port 42 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 io_wbs_m2s_addr[12]
port 43 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 io_wbs_m2s_addr[13]
port 44 nsew signal input
rlabel metal3 s 19200 18368 20000 18488 6 io_wbs_m2s_addr[14]
port 45 nsew signal input
rlabel metal2 s 3882 19200 3938 20000 6 io_wbs_m2s_addr[15]
port 46 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 io_wbs_m2s_addr[1]
port 47 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 io_wbs_m2s_addr[2]
port 48 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 io_wbs_m2s_addr[3]
port 49 nsew signal input
rlabel metal3 s 19200 6808 20000 6928 6 io_wbs_m2s_addr[4]
port 50 nsew signal input
rlabel metal3 s 19200 3408 20000 3528 6 io_wbs_m2s_addr[5]
port 51 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 io_wbs_m2s_addr[6]
port 52 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_wbs_m2s_addr[7]
port 53 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_wbs_m2s_addr[8]
port 54 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 io_wbs_m2s_addr[9]
port 55 nsew signal input
rlabel metal3 s 19200 4768 20000 4888 6 io_wbs_m2s_data[0]
port 56 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 io_wbs_m2s_data[10]
port 57 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_wbs_m2s_data[11]
port 58 nsew signal input
rlabel metal3 s 19200 12248 20000 12368 6 io_wbs_m2s_data[12]
port 59 nsew signal input
rlabel metal2 s 5170 19200 5226 20000 6 io_wbs_m2s_data[13]
port 60 nsew signal input
rlabel metal2 s 2594 19200 2650 20000 6 io_wbs_m2s_data[14]
port 61 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 io_wbs_m2s_data[15]
port 62 nsew signal input
rlabel metal2 s 18 0 74 800 6 io_wbs_m2s_data[16]
port 63 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 io_wbs_m2s_data[17]
port 64 nsew signal input
rlabel metal2 s 6458 19200 6514 20000 6 io_wbs_m2s_data[18]
port 65 nsew signal input
rlabel metal2 s 11610 19200 11666 20000 6 io_wbs_m2s_data[19]
port 66 nsew signal input
rlabel metal2 s 16762 19200 16818 20000 6 io_wbs_m2s_data[1]
port 67 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 io_wbs_m2s_data[20]
port 68 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 io_wbs_m2s_data[21]
port 69 nsew signal input
rlabel metal2 s 662 0 718 800 6 io_wbs_m2s_data[22]
port 70 nsew signal input
rlabel metal2 s 19338 19200 19394 20000 6 io_wbs_m2s_data[23]
port 71 nsew signal input
rlabel metal2 s 14830 19200 14886 20000 6 io_wbs_m2s_data[24]
port 72 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_wbs_m2s_data[25]
port 73 nsew signal input
rlabel metal3 s 19200 19728 20000 19848 6 io_wbs_m2s_data[26]
port 74 nsew signal input
rlabel metal3 s 19200 1368 20000 1488 6 io_wbs_m2s_data[27]
port 75 nsew signal input
rlabel metal2 s 1950 19200 2006 20000 6 io_wbs_m2s_data[28]
port 76 nsew signal input
rlabel metal3 s 19200 10208 20000 10328 6 io_wbs_m2s_data[29]
port 77 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 io_wbs_m2s_data[2]
port 78 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 io_wbs_m2s_data[30]
port 79 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 io_wbs_m2s_data[31]
port 80 nsew signal input
rlabel metal3 s 19200 11568 20000 11688 6 io_wbs_m2s_data[3]
port 81 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 io_wbs_m2s_data[4]
port 82 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 io_wbs_m2s_data[5]
port 83 nsew signal input
rlabel metal2 s 15474 19200 15530 20000 6 io_wbs_m2s_data[6]
port 84 nsew signal input
rlabel metal2 s 1306 19200 1362 20000 6 io_wbs_m2s_data[7]
port 85 nsew signal input
rlabel metal2 s 4526 19200 4582 20000 6 io_wbs_m2s_data[8]
port 86 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 io_wbs_m2s_data[9]
port 87 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 io_wbs_m2s_stb
port 88 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 io_wbs_m2s_we
port 89 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 reset
port 90 nsew signal input
rlabel metal4 s 3910 2128 4230 17456 6 vccd1
port 91 nsew power input
rlabel metal4 s 9840 2128 10160 17456 6 vccd1
port 91 nsew power input
rlabel metal4 s 15771 2128 16091 17456 6 vccd1
port 91 nsew power input
rlabel metal4 s 6874 2128 7194 17456 6 vssd1
port 92 nsew ground input
rlabel metal4 s 12805 2128 13125 17456 6 vssd1
port 92 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
