magic
tech sky130A
magscale 1 2
timestamp 1647766204
<< nwell >>
rect 1066 97093 98846 97414
rect 1066 96005 98846 96571
rect 1066 94917 98846 95483
rect 1066 93829 98846 94395
rect 1066 92741 98846 93307
rect 1066 91653 98846 92219
rect 1066 90565 98846 91131
rect 1066 89477 98846 90043
rect 1066 88389 98846 88955
rect 1066 87301 98846 87867
rect 1066 86213 98846 86779
rect 1066 85125 98846 85691
rect 1066 84037 98846 84603
rect 1066 82949 98846 83515
rect 1066 81861 98846 82427
rect 1066 80773 98846 81339
rect 1066 79685 98846 80251
rect 1066 78597 98846 79163
rect 1066 77509 98846 78075
rect 1066 76421 98846 76987
rect 1066 75333 98846 75899
rect 1066 74245 98846 74811
rect 1066 73157 98846 73723
rect 1066 72069 98846 72635
rect 1066 70981 98846 71547
rect 1066 69893 98846 70459
rect 1066 68805 98846 69371
rect 1066 67717 98846 68283
rect 1066 66629 98846 67195
rect 1066 65541 98846 66107
rect 1066 64453 98846 65019
rect 1066 63365 98846 63931
rect 1066 62277 98846 62843
rect 1066 61189 98846 61755
rect 1066 60101 98846 60667
rect 1066 59013 98846 59579
rect 1066 57925 98846 58491
rect 1066 56837 98846 57403
rect 1066 55749 98846 56315
rect 1066 54661 98846 55227
rect 1066 53573 98846 54139
rect 1066 52485 98846 53051
rect 1066 51397 98846 51963
rect 1066 50309 98846 50875
rect 1066 49221 98846 49787
rect 1066 48133 98846 48699
rect 1066 47045 98846 47611
rect 1066 45957 98846 46523
rect 1066 44869 98846 45435
rect 1066 43781 98846 44347
rect 1066 42693 98846 43259
rect 1066 41605 98846 42171
rect 1066 40517 98846 41083
rect 1066 39429 98846 39995
rect 1066 38341 98846 38907
rect 1066 37253 98846 37819
rect 1066 36165 98846 36731
rect 1066 35077 98846 35643
rect 1066 33989 98846 34555
rect 1066 32901 98846 33467
rect 1066 31813 98846 32379
rect 1066 30725 98846 31291
rect 1066 29637 98846 30203
rect 1066 28549 98846 29115
rect 1066 27461 98846 28027
rect 1066 26373 98846 26939
rect 1066 25285 98846 25851
rect 1066 24197 98846 24763
rect 1066 23109 98846 23675
rect 1066 22021 98846 22587
rect 1066 20933 98846 21499
rect 1066 19845 98846 20411
rect 1066 18757 98846 19323
rect 1066 17669 98846 18235
rect 1066 16581 98846 17147
rect 1066 15493 98846 16059
rect 1066 14405 98846 14971
rect 1066 13317 98846 13883
rect 1066 12229 98846 12795
rect 1066 11141 98846 11707
rect 1066 10053 98846 10619
rect 1066 8965 98846 9531
rect 1066 7877 98846 8443
rect 1066 6789 98846 7355
rect 1066 5701 98846 6267
rect 1066 4613 98846 5179
rect 1066 3525 98846 4091
rect 1066 2437 98846 3003
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2048 99990 97708
<< metal2 >>
rect 49974 99200 50030 100000
rect 24950 0 25006 800
rect 74906 0 74962 800
<< obsm2 >>
rect 1400 99144 49918 99657
rect 50086 99144 99986 99657
rect 1400 856 99986 99144
rect 1400 303 24894 856
rect 25062 303 74850 856
rect 75018 303 99986 856
<< metal3 >>
rect 99200 99560 100000 99680
rect 99200 99016 100000 99136
rect 99200 98472 100000 98592
rect 99200 97792 100000 97912
rect 99200 97248 100000 97368
rect 99200 96704 100000 96824
rect 99200 96024 100000 96144
rect 99200 95480 100000 95600
rect 99200 94936 100000 95056
rect 99200 94392 100000 94512
rect 99200 93712 100000 93832
rect 99200 93168 100000 93288
rect 99200 92624 100000 92744
rect 99200 91944 100000 92064
rect 99200 91400 100000 91520
rect 99200 90856 100000 90976
rect 99200 90176 100000 90296
rect 99200 89632 100000 89752
rect 99200 89088 100000 89208
rect 99200 88544 100000 88664
rect 99200 87864 100000 87984
rect 99200 87320 100000 87440
rect 99200 86776 100000 86896
rect 99200 86096 100000 86216
rect 99200 85552 100000 85672
rect 99200 85008 100000 85128
rect 99200 84328 100000 84448
rect 99200 83784 100000 83904
rect 99200 83240 100000 83360
rect 99200 82696 100000 82816
rect 99200 82016 100000 82136
rect 99200 81472 100000 81592
rect 99200 80928 100000 81048
rect 99200 80248 100000 80368
rect 99200 79704 100000 79824
rect 99200 79160 100000 79280
rect 99200 78480 100000 78600
rect 99200 77936 100000 78056
rect 99200 77392 100000 77512
rect 99200 76848 100000 76968
rect 99200 76168 100000 76288
rect 99200 75624 100000 75744
rect 99200 75080 100000 75200
rect 99200 74400 100000 74520
rect 99200 73856 100000 73976
rect 99200 73312 100000 73432
rect 99200 72632 100000 72752
rect 99200 72088 100000 72208
rect 99200 71544 100000 71664
rect 99200 71000 100000 71120
rect 99200 70320 100000 70440
rect 99200 69776 100000 69896
rect 99200 69232 100000 69352
rect 99200 68552 100000 68672
rect 99200 68008 100000 68128
rect 99200 67464 100000 67584
rect 99200 66920 100000 67040
rect 99200 66240 100000 66360
rect 99200 65696 100000 65816
rect 99200 65152 100000 65272
rect 99200 64472 100000 64592
rect 99200 63928 100000 64048
rect 99200 63384 100000 63504
rect 99200 62704 100000 62824
rect 99200 62160 100000 62280
rect 99200 61616 100000 61736
rect 99200 61072 100000 61192
rect 99200 60392 100000 60512
rect 99200 59848 100000 59968
rect 99200 59304 100000 59424
rect 99200 58624 100000 58744
rect 99200 58080 100000 58200
rect 99200 57536 100000 57656
rect 99200 56856 100000 56976
rect 99200 56312 100000 56432
rect 99200 55768 100000 55888
rect 99200 55224 100000 55344
rect 99200 54544 100000 54664
rect 99200 54000 100000 54120
rect 99200 53456 100000 53576
rect 99200 52776 100000 52896
rect 99200 52232 100000 52352
rect 99200 51688 100000 51808
rect 99200 51008 100000 51128
rect 99200 50464 100000 50584
rect 99200 49920 100000 50040
rect 99200 49376 100000 49496
rect 99200 48696 100000 48816
rect 99200 48152 100000 48272
rect 99200 47608 100000 47728
rect 99200 46928 100000 47048
rect 99200 46384 100000 46504
rect 99200 45840 100000 45960
rect 99200 45160 100000 45280
rect 99200 44616 100000 44736
rect 99200 44072 100000 44192
rect 99200 43528 100000 43648
rect 99200 42848 100000 42968
rect 99200 42304 100000 42424
rect 99200 41760 100000 41880
rect 99200 41080 100000 41200
rect 99200 40536 100000 40656
rect 99200 39992 100000 40112
rect 99200 39312 100000 39432
rect 99200 38768 100000 38888
rect 99200 38224 100000 38344
rect 99200 37680 100000 37800
rect 99200 37000 100000 37120
rect 99200 36456 100000 36576
rect 99200 35912 100000 36032
rect 99200 35232 100000 35352
rect 99200 34688 100000 34808
rect 99200 34144 100000 34264
rect 99200 33600 100000 33720
rect 99200 32920 100000 33040
rect 99200 32376 100000 32496
rect 99200 31832 100000 31952
rect 99200 31152 100000 31272
rect 99200 30608 100000 30728
rect 99200 30064 100000 30184
rect 99200 29384 100000 29504
rect 99200 28840 100000 28960
rect 99200 28296 100000 28416
rect 99200 27752 100000 27872
rect 99200 27072 100000 27192
rect 99200 26528 100000 26648
rect 99200 25984 100000 26104
rect 99200 25304 100000 25424
rect 99200 24760 100000 24880
rect 99200 24216 100000 24336
rect 99200 23536 100000 23656
rect 99200 22992 100000 23112
rect 99200 22448 100000 22568
rect 99200 21904 100000 22024
rect 99200 21224 100000 21344
rect 99200 20680 100000 20800
rect 99200 20136 100000 20256
rect 99200 19456 100000 19576
rect 99200 18912 100000 19032
rect 99200 18368 100000 18488
rect 99200 17688 100000 17808
rect 99200 17144 100000 17264
rect 99200 16600 100000 16720
rect 99200 16056 100000 16176
rect 99200 15376 100000 15496
rect 99200 14832 100000 14952
rect 99200 14288 100000 14408
rect 99200 13608 100000 13728
rect 99200 13064 100000 13184
rect 99200 12520 100000 12640
rect 99200 11840 100000 11960
rect 99200 11296 100000 11416
rect 99200 10752 100000 10872
rect 99200 10208 100000 10328
rect 99200 9528 100000 9648
rect 99200 8984 100000 9104
rect 99200 8440 100000 8560
rect 99200 7760 100000 7880
rect 99200 7216 100000 7336
rect 99200 6672 100000 6792
rect 99200 5992 100000 6112
rect 99200 5448 100000 5568
rect 99200 4904 100000 5024
rect 99200 4360 100000 4480
rect 99200 3680 100000 3800
rect 99200 3136 100000 3256
rect 99200 2592 100000 2712
rect 99200 1912 100000 2032
rect 99200 1368 100000 1488
rect 99200 824 100000 944
rect 99200 280 100000 400
<< obsm3 >>
rect 3141 99480 99120 99653
rect 3141 99216 99991 99480
rect 3141 98936 99120 99216
rect 3141 98672 99991 98936
rect 3141 98392 99120 98672
rect 3141 97992 99991 98392
rect 3141 97712 99120 97992
rect 3141 97448 99991 97712
rect 3141 97168 99120 97448
rect 3141 96904 99991 97168
rect 3141 96624 99120 96904
rect 3141 96224 99991 96624
rect 3141 95944 99120 96224
rect 3141 95680 99991 95944
rect 3141 95400 99120 95680
rect 3141 95136 99991 95400
rect 3141 94856 99120 95136
rect 3141 94592 99991 94856
rect 3141 94312 99120 94592
rect 3141 93912 99991 94312
rect 3141 93632 99120 93912
rect 3141 93368 99991 93632
rect 3141 93088 99120 93368
rect 3141 92824 99991 93088
rect 3141 92544 99120 92824
rect 3141 92144 99991 92544
rect 3141 91864 99120 92144
rect 3141 91600 99991 91864
rect 3141 91320 99120 91600
rect 3141 91056 99991 91320
rect 3141 90776 99120 91056
rect 3141 90376 99991 90776
rect 3141 90096 99120 90376
rect 3141 89832 99991 90096
rect 3141 89552 99120 89832
rect 3141 89288 99991 89552
rect 3141 89008 99120 89288
rect 3141 88744 99991 89008
rect 3141 88464 99120 88744
rect 3141 88064 99991 88464
rect 3141 87784 99120 88064
rect 3141 87520 99991 87784
rect 3141 87240 99120 87520
rect 3141 86976 99991 87240
rect 3141 86696 99120 86976
rect 3141 86296 99991 86696
rect 3141 86016 99120 86296
rect 3141 85752 99991 86016
rect 3141 85472 99120 85752
rect 3141 85208 99991 85472
rect 3141 84928 99120 85208
rect 3141 84528 99991 84928
rect 3141 84248 99120 84528
rect 3141 83984 99991 84248
rect 3141 83704 99120 83984
rect 3141 83440 99991 83704
rect 3141 83160 99120 83440
rect 3141 82896 99991 83160
rect 3141 82616 99120 82896
rect 3141 82216 99991 82616
rect 3141 81936 99120 82216
rect 3141 81672 99991 81936
rect 3141 81392 99120 81672
rect 3141 81128 99991 81392
rect 3141 80848 99120 81128
rect 3141 80448 99991 80848
rect 3141 80168 99120 80448
rect 3141 79904 99991 80168
rect 3141 79624 99120 79904
rect 3141 79360 99991 79624
rect 3141 79080 99120 79360
rect 3141 78680 99991 79080
rect 3141 78400 99120 78680
rect 3141 78136 99991 78400
rect 3141 77856 99120 78136
rect 3141 77592 99991 77856
rect 3141 77312 99120 77592
rect 3141 77048 99991 77312
rect 3141 76768 99120 77048
rect 3141 76368 99991 76768
rect 3141 76088 99120 76368
rect 3141 75824 99991 76088
rect 3141 75544 99120 75824
rect 3141 75280 99991 75544
rect 3141 75000 99120 75280
rect 3141 74600 99991 75000
rect 3141 74320 99120 74600
rect 3141 74056 99991 74320
rect 3141 73776 99120 74056
rect 3141 73512 99991 73776
rect 3141 73232 99120 73512
rect 3141 72832 99991 73232
rect 3141 72552 99120 72832
rect 3141 72288 99991 72552
rect 3141 72008 99120 72288
rect 3141 71744 99991 72008
rect 3141 71464 99120 71744
rect 3141 71200 99991 71464
rect 3141 70920 99120 71200
rect 3141 70520 99991 70920
rect 3141 70240 99120 70520
rect 3141 69976 99991 70240
rect 3141 69696 99120 69976
rect 3141 69432 99991 69696
rect 3141 69152 99120 69432
rect 3141 68752 99991 69152
rect 3141 68472 99120 68752
rect 3141 68208 99991 68472
rect 3141 67928 99120 68208
rect 3141 67664 99991 67928
rect 3141 67384 99120 67664
rect 3141 67120 99991 67384
rect 3141 66840 99120 67120
rect 3141 66440 99991 66840
rect 3141 66160 99120 66440
rect 3141 65896 99991 66160
rect 3141 65616 99120 65896
rect 3141 65352 99991 65616
rect 3141 65072 99120 65352
rect 3141 64672 99991 65072
rect 3141 64392 99120 64672
rect 3141 64128 99991 64392
rect 3141 63848 99120 64128
rect 3141 63584 99991 63848
rect 3141 63304 99120 63584
rect 3141 62904 99991 63304
rect 3141 62624 99120 62904
rect 3141 62360 99991 62624
rect 3141 62080 99120 62360
rect 3141 61816 99991 62080
rect 3141 61536 99120 61816
rect 3141 61272 99991 61536
rect 3141 60992 99120 61272
rect 3141 60592 99991 60992
rect 3141 60312 99120 60592
rect 3141 60048 99991 60312
rect 3141 59768 99120 60048
rect 3141 59504 99991 59768
rect 3141 59224 99120 59504
rect 3141 58824 99991 59224
rect 3141 58544 99120 58824
rect 3141 58280 99991 58544
rect 3141 58000 99120 58280
rect 3141 57736 99991 58000
rect 3141 57456 99120 57736
rect 3141 57056 99991 57456
rect 3141 56776 99120 57056
rect 3141 56512 99991 56776
rect 3141 56232 99120 56512
rect 3141 55968 99991 56232
rect 3141 55688 99120 55968
rect 3141 55424 99991 55688
rect 3141 55144 99120 55424
rect 3141 54744 99991 55144
rect 3141 54464 99120 54744
rect 3141 54200 99991 54464
rect 3141 53920 99120 54200
rect 3141 53656 99991 53920
rect 3141 53376 99120 53656
rect 3141 52976 99991 53376
rect 3141 52696 99120 52976
rect 3141 52432 99991 52696
rect 3141 52152 99120 52432
rect 3141 51888 99991 52152
rect 3141 51608 99120 51888
rect 3141 51208 99991 51608
rect 3141 50928 99120 51208
rect 3141 50664 99991 50928
rect 3141 50384 99120 50664
rect 3141 50120 99991 50384
rect 3141 49840 99120 50120
rect 3141 49576 99991 49840
rect 3141 49296 99120 49576
rect 3141 48896 99991 49296
rect 3141 48616 99120 48896
rect 3141 48352 99991 48616
rect 3141 48072 99120 48352
rect 3141 47808 99991 48072
rect 3141 47528 99120 47808
rect 3141 47128 99991 47528
rect 3141 46848 99120 47128
rect 3141 46584 99991 46848
rect 3141 46304 99120 46584
rect 3141 46040 99991 46304
rect 3141 45760 99120 46040
rect 3141 45360 99991 45760
rect 3141 45080 99120 45360
rect 3141 44816 99991 45080
rect 3141 44536 99120 44816
rect 3141 44272 99991 44536
rect 3141 43992 99120 44272
rect 3141 43728 99991 43992
rect 3141 43448 99120 43728
rect 3141 43048 99991 43448
rect 3141 42768 99120 43048
rect 3141 42504 99991 42768
rect 3141 42224 99120 42504
rect 3141 41960 99991 42224
rect 3141 41680 99120 41960
rect 3141 41280 99991 41680
rect 3141 41000 99120 41280
rect 3141 40736 99991 41000
rect 3141 40456 99120 40736
rect 3141 40192 99991 40456
rect 3141 39912 99120 40192
rect 3141 39512 99991 39912
rect 3141 39232 99120 39512
rect 3141 38968 99991 39232
rect 3141 38688 99120 38968
rect 3141 38424 99991 38688
rect 3141 38144 99120 38424
rect 3141 37880 99991 38144
rect 3141 37600 99120 37880
rect 3141 37200 99991 37600
rect 3141 36920 99120 37200
rect 3141 36656 99991 36920
rect 3141 36376 99120 36656
rect 3141 36112 99991 36376
rect 3141 35832 99120 36112
rect 3141 35432 99991 35832
rect 3141 35152 99120 35432
rect 3141 34888 99991 35152
rect 3141 34608 99120 34888
rect 3141 34344 99991 34608
rect 3141 34064 99120 34344
rect 3141 33800 99991 34064
rect 3141 33520 99120 33800
rect 3141 33120 99991 33520
rect 3141 32840 99120 33120
rect 3141 32576 99991 32840
rect 3141 32296 99120 32576
rect 3141 32032 99991 32296
rect 3141 31752 99120 32032
rect 3141 31352 99991 31752
rect 3141 31072 99120 31352
rect 3141 30808 99991 31072
rect 3141 30528 99120 30808
rect 3141 30264 99991 30528
rect 3141 29984 99120 30264
rect 3141 29584 99991 29984
rect 3141 29304 99120 29584
rect 3141 29040 99991 29304
rect 3141 28760 99120 29040
rect 3141 28496 99991 28760
rect 3141 28216 99120 28496
rect 3141 27952 99991 28216
rect 3141 27672 99120 27952
rect 3141 27272 99991 27672
rect 3141 26992 99120 27272
rect 3141 26728 99991 26992
rect 3141 26448 99120 26728
rect 3141 26184 99991 26448
rect 3141 25904 99120 26184
rect 3141 25504 99991 25904
rect 3141 25224 99120 25504
rect 3141 24960 99991 25224
rect 3141 24680 99120 24960
rect 3141 24416 99991 24680
rect 3141 24136 99120 24416
rect 3141 23736 99991 24136
rect 3141 23456 99120 23736
rect 3141 23192 99991 23456
rect 3141 22912 99120 23192
rect 3141 22648 99991 22912
rect 3141 22368 99120 22648
rect 3141 22104 99991 22368
rect 3141 21824 99120 22104
rect 3141 21424 99991 21824
rect 3141 21144 99120 21424
rect 3141 20880 99991 21144
rect 3141 20600 99120 20880
rect 3141 20336 99991 20600
rect 3141 20056 99120 20336
rect 3141 19656 99991 20056
rect 3141 19376 99120 19656
rect 3141 19112 99991 19376
rect 3141 18832 99120 19112
rect 3141 18568 99991 18832
rect 3141 18288 99120 18568
rect 3141 17888 99991 18288
rect 3141 17608 99120 17888
rect 3141 17344 99991 17608
rect 3141 17064 99120 17344
rect 3141 16800 99991 17064
rect 3141 16520 99120 16800
rect 3141 16256 99991 16520
rect 3141 15976 99120 16256
rect 3141 15576 99991 15976
rect 3141 15296 99120 15576
rect 3141 15032 99991 15296
rect 3141 14752 99120 15032
rect 3141 14488 99991 14752
rect 3141 14208 99120 14488
rect 3141 13808 99991 14208
rect 3141 13528 99120 13808
rect 3141 13264 99991 13528
rect 3141 12984 99120 13264
rect 3141 12720 99991 12984
rect 3141 12440 99120 12720
rect 3141 12040 99991 12440
rect 3141 11760 99120 12040
rect 3141 11496 99991 11760
rect 3141 11216 99120 11496
rect 3141 10952 99991 11216
rect 3141 10672 99120 10952
rect 3141 10408 99991 10672
rect 3141 10128 99120 10408
rect 3141 9728 99991 10128
rect 3141 9448 99120 9728
rect 3141 9184 99991 9448
rect 3141 8904 99120 9184
rect 3141 8640 99991 8904
rect 3141 8360 99120 8640
rect 3141 7960 99991 8360
rect 3141 7680 99120 7960
rect 3141 7416 99991 7680
rect 3141 7136 99120 7416
rect 3141 6872 99991 7136
rect 3141 6592 99120 6872
rect 3141 6192 99991 6592
rect 3141 5912 99120 6192
rect 3141 5648 99991 5912
rect 3141 5368 99120 5648
rect 3141 5104 99991 5368
rect 3141 4824 99120 5104
rect 3141 4560 99991 4824
rect 3141 4280 99120 4560
rect 3141 3880 99991 4280
rect 3141 3600 99120 3880
rect 3141 3336 99991 3600
rect 3141 3056 99120 3336
rect 3141 2792 99991 3056
rect 3141 2512 99120 2792
rect 3141 2112 99991 2512
rect 3141 1832 99120 2112
rect 3141 1568 99991 1832
rect 3141 1288 99120 1568
rect 3141 1024 99991 1288
rect 3141 744 99120 1024
rect 3141 480 99991 744
rect 3141 307 99120 480
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 8339 2619 19488 97205
rect 19968 2619 34848 97205
rect 35328 2619 50208 97205
rect 50688 2619 65568 97205
rect 66048 2619 80928 97205
rect 81408 2619 96288 97205
rect 96768 2619 98197 97205
<< labels >>
rlabel metal2 s 24950 0 25006 800 6 clock
port 1 nsew signal input
rlabel metal3 s 99200 1912 100000 2032 6 io_dbus_addr[0]
port 2 nsew signal output
rlabel metal3 s 99200 22448 100000 22568 6 io_dbus_addr[10]
port 3 nsew signal output
rlabel metal3 s 99200 24216 100000 24336 6 io_dbus_addr[11]
port 4 nsew signal output
rlabel metal3 s 99200 25984 100000 26104 6 io_dbus_addr[12]
port 5 nsew signal output
rlabel metal3 s 99200 27752 100000 27872 6 io_dbus_addr[13]
port 6 nsew signal output
rlabel metal3 s 99200 29384 100000 29504 6 io_dbus_addr[14]
port 7 nsew signal output
rlabel metal3 s 99200 31152 100000 31272 6 io_dbus_addr[15]
port 8 nsew signal output
rlabel metal3 s 99200 32920 100000 33040 6 io_dbus_addr[16]
port 9 nsew signal output
rlabel metal3 s 99200 34688 100000 34808 6 io_dbus_addr[17]
port 10 nsew signal output
rlabel metal3 s 99200 36456 100000 36576 6 io_dbus_addr[18]
port 11 nsew signal output
rlabel metal3 s 99200 38224 100000 38344 6 io_dbus_addr[19]
port 12 nsew signal output
rlabel metal3 s 99200 4904 100000 5024 6 io_dbus_addr[1]
port 13 nsew signal output
rlabel metal3 s 99200 39992 100000 40112 6 io_dbus_addr[20]
port 14 nsew signal output
rlabel metal3 s 99200 41760 100000 41880 6 io_dbus_addr[21]
port 15 nsew signal output
rlabel metal3 s 99200 43528 100000 43648 6 io_dbus_addr[22]
port 16 nsew signal output
rlabel metal3 s 99200 45160 100000 45280 6 io_dbus_addr[23]
port 17 nsew signal output
rlabel metal3 s 99200 46928 100000 47048 6 io_dbus_addr[24]
port 18 nsew signal output
rlabel metal3 s 99200 48696 100000 48816 6 io_dbus_addr[25]
port 19 nsew signal output
rlabel metal3 s 99200 50464 100000 50584 6 io_dbus_addr[26]
port 20 nsew signal output
rlabel metal3 s 99200 52232 100000 52352 6 io_dbus_addr[27]
port 21 nsew signal output
rlabel metal3 s 99200 54000 100000 54120 6 io_dbus_addr[28]
port 22 nsew signal output
rlabel metal3 s 99200 55768 100000 55888 6 io_dbus_addr[29]
port 23 nsew signal output
rlabel metal3 s 99200 7760 100000 7880 6 io_dbus_addr[2]
port 24 nsew signal output
rlabel metal3 s 99200 57536 100000 57656 6 io_dbus_addr[30]
port 25 nsew signal output
rlabel metal3 s 99200 59304 100000 59424 6 io_dbus_addr[31]
port 26 nsew signal output
rlabel metal3 s 99200 10208 100000 10328 6 io_dbus_addr[3]
port 27 nsew signal output
rlabel metal3 s 99200 11840 100000 11960 6 io_dbus_addr[4]
port 28 nsew signal output
rlabel metal3 s 99200 13608 100000 13728 6 io_dbus_addr[5]
port 29 nsew signal output
rlabel metal3 s 99200 15376 100000 15496 6 io_dbus_addr[6]
port 30 nsew signal output
rlabel metal3 s 99200 17144 100000 17264 6 io_dbus_addr[7]
port 31 nsew signal output
rlabel metal3 s 99200 18912 100000 19032 6 io_dbus_addr[8]
port 32 nsew signal output
rlabel metal3 s 99200 20680 100000 20800 6 io_dbus_addr[9]
port 33 nsew signal output
rlabel metal3 s 99200 2592 100000 2712 6 io_dbus_ld_type[0]
port 34 nsew signal output
rlabel metal3 s 99200 5448 100000 5568 6 io_dbus_ld_type[1]
port 35 nsew signal output
rlabel metal3 s 99200 8440 100000 8560 6 io_dbus_ld_type[2]
port 36 nsew signal output
rlabel metal3 s 99200 280 100000 400 6 io_dbus_rd_en
port 37 nsew signal output
rlabel metal3 s 99200 3136 100000 3256 6 io_dbus_rdata[0]
port 38 nsew signal input
rlabel metal3 s 99200 22992 100000 23112 6 io_dbus_rdata[10]
port 39 nsew signal input
rlabel metal3 s 99200 24760 100000 24880 6 io_dbus_rdata[11]
port 40 nsew signal input
rlabel metal3 s 99200 26528 100000 26648 6 io_dbus_rdata[12]
port 41 nsew signal input
rlabel metal3 s 99200 28296 100000 28416 6 io_dbus_rdata[13]
port 42 nsew signal input
rlabel metal3 s 99200 30064 100000 30184 6 io_dbus_rdata[14]
port 43 nsew signal input
rlabel metal3 s 99200 31832 100000 31952 6 io_dbus_rdata[15]
port 44 nsew signal input
rlabel metal3 s 99200 33600 100000 33720 6 io_dbus_rdata[16]
port 45 nsew signal input
rlabel metal3 s 99200 35232 100000 35352 6 io_dbus_rdata[17]
port 46 nsew signal input
rlabel metal3 s 99200 37000 100000 37120 6 io_dbus_rdata[18]
port 47 nsew signal input
rlabel metal3 s 99200 38768 100000 38888 6 io_dbus_rdata[19]
port 48 nsew signal input
rlabel metal3 s 99200 5992 100000 6112 6 io_dbus_rdata[1]
port 49 nsew signal input
rlabel metal3 s 99200 40536 100000 40656 6 io_dbus_rdata[20]
port 50 nsew signal input
rlabel metal3 s 99200 42304 100000 42424 6 io_dbus_rdata[21]
port 51 nsew signal input
rlabel metal3 s 99200 44072 100000 44192 6 io_dbus_rdata[22]
port 52 nsew signal input
rlabel metal3 s 99200 45840 100000 45960 6 io_dbus_rdata[23]
port 53 nsew signal input
rlabel metal3 s 99200 47608 100000 47728 6 io_dbus_rdata[24]
port 54 nsew signal input
rlabel metal3 s 99200 49376 100000 49496 6 io_dbus_rdata[25]
port 55 nsew signal input
rlabel metal3 s 99200 51008 100000 51128 6 io_dbus_rdata[26]
port 56 nsew signal input
rlabel metal3 s 99200 52776 100000 52896 6 io_dbus_rdata[27]
port 57 nsew signal input
rlabel metal3 s 99200 54544 100000 54664 6 io_dbus_rdata[28]
port 58 nsew signal input
rlabel metal3 s 99200 56312 100000 56432 6 io_dbus_rdata[29]
port 59 nsew signal input
rlabel metal3 s 99200 8984 100000 9104 6 io_dbus_rdata[2]
port 60 nsew signal input
rlabel metal3 s 99200 58080 100000 58200 6 io_dbus_rdata[30]
port 61 nsew signal input
rlabel metal3 s 99200 59848 100000 59968 6 io_dbus_rdata[31]
port 62 nsew signal input
rlabel metal3 s 99200 10752 100000 10872 6 io_dbus_rdata[3]
port 63 nsew signal input
rlabel metal3 s 99200 12520 100000 12640 6 io_dbus_rdata[4]
port 64 nsew signal input
rlabel metal3 s 99200 14288 100000 14408 6 io_dbus_rdata[5]
port 65 nsew signal input
rlabel metal3 s 99200 16056 100000 16176 6 io_dbus_rdata[6]
port 66 nsew signal input
rlabel metal3 s 99200 17688 100000 17808 6 io_dbus_rdata[7]
port 67 nsew signal input
rlabel metal3 s 99200 19456 100000 19576 6 io_dbus_rdata[8]
port 68 nsew signal input
rlabel metal3 s 99200 21224 100000 21344 6 io_dbus_rdata[9]
port 69 nsew signal input
rlabel metal3 s 99200 3680 100000 3800 6 io_dbus_st_type[0]
port 70 nsew signal output
rlabel metal3 s 99200 6672 100000 6792 6 io_dbus_st_type[1]
port 71 nsew signal output
rlabel metal3 s 99200 824 100000 944 6 io_dbus_valid
port 72 nsew signal input
rlabel metal3 s 99200 4360 100000 4480 6 io_dbus_wdata[0]
port 73 nsew signal output
rlabel metal3 s 99200 23536 100000 23656 6 io_dbus_wdata[10]
port 74 nsew signal output
rlabel metal3 s 99200 25304 100000 25424 6 io_dbus_wdata[11]
port 75 nsew signal output
rlabel metal3 s 99200 27072 100000 27192 6 io_dbus_wdata[12]
port 76 nsew signal output
rlabel metal3 s 99200 28840 100000 28960 6 io_dbus_wdata[13]
port 77 nsew signal output
rlabel metal3 s 99200 30608 100000 30728 6 io_dbus_wdata[14]
port 78 nsew signal output
rlabel metal3 s 99200 32376 100000 32496 6 io_dbus_wdata[15]
port 79 nsew signal output
rlabel metal3 s 99200 34144 100000 34264 6 io_dbus_wdata[16]
port 80 nsew signal output
rlabel metal3 s 99200 35912 100000 36032 6 io_dbus_wdata[17]
port 81 nsew signal output
rlabel metal3 s 99200 37680 100000 37800 6 io_dbus_wdata[18]
port 82 nsew signal output
rlabel metal3 s 99200 39312 100000 39432 6 io_dbus_wdata[19]
port 83 nsew signal output
rlabel metal3 s 99200 7216 100000 7336 6 io_dbus_wdata[1]
port 84 nsew signal output
rlabel metal3 s 99200 41080 100000 41200 6 io_dbus_wdata[20]
port 85 nsew signal output
rlabel metal3 s 99200 42848 100000 42968 6 io_dbus_wdata[21]
port 86 nsew signal output
rlabel metal3 s 99200 44616 100000 44736 6 io_dbus_wdata[22]
port 87 nsew signal output
rlabel metal3 s 99200 46384 100000 46504 6 io_dbus_wdata[23]
port 88 nsew signal output
rlabel metal3 s 99200 48152 100000 48272 6 io_dbus_wdata[24]
port 89 nsew signal output
rlabel metal3 s 99200 49920 100000 50040 6 io_dbus_wdata[25]
port 90 nsew signal output
rlabel metal3 s 99200 51688 100000 51808 6 io_dbus_wdata[26]
port 91 nsew signal output
rlabel metal3 s 99200 53456 100000 53576 6 io_dbus_wdata[27]
port 92 nsew signal output
rlabel metal3 s 99200 55224 100000 55344 6 io_dbus_wdata[28]
port 93 nsew signal output
rlabel metal3 s 99200 56856 100000 56976 6 io_dbus_wdata[29]
port 94 nsew signal output
rlabel metal3 s 99200 9528 100000 9648 6 io_dbus_wdata[2]
port 95 nsew signal output
rlabel metal3 s 99200 58624 100000 58744 6 io_dbus_wdata[30]
port 96 nsew signal output
rlabel metal3 s 99200 60392 100000 60512 6 io_dbus_wdata[31]
port 97 nsew signal output
rlabel metal3 s 99200 11296 100000 11416 6 io_dbus_wdata[3]
port 98 nsew signal output
rlabel metal3 s 99200 13064 100000 13184 6 io_dbus_wdata[4]
port 99 nsew signal output
rlabel metal3 s 99200 14832 100000 14952 6 io_dbus_wdata[5]
port 100 nsew signal output
rlabel metal3 s 99200 16600 100000 16720 6 io_dbus_wdata[6]
port 101 nsew signal output
rlabel metal3 s 99200 18368 100000 18488 6 io_dbus_wdata[7]
port 102 nsew signal output
rlabel metal3 s 99200 20136 100000 20256 6 io_dbus_wdata[8]
port 103 nsew signal output
rlabel metal3 s 99200 21904 100000 22024 6 io_dbus_wdata[9]
port 104 nsew signal output
rlabel metal3 s 99200 1368 100000 1488 6 io_dbus_wr_en
port 105 nsew signal output
rlabel metal3 s 99200 61616 100000 61736 6 io_ibus_addr[0]
port 106 nsew signal output
rlabel metal3 s 99200 73312 100000 73432 6 io_ibus_addr[10]
port 107 nsew signal output
rlabel metal3 s 99200 74400 100000 74520 6 io_ibus_addr[11]
port 108 nsew signal output
rlabel metal3 s 99200 75624 100000 75744 6 io_ibus_addr[12]
port 109 nsew signal output
rlabel metal3 s 99200 76848 100000 76968 6 io_ibus_addr[13]
port 110 nsew signal output
rlabel metal3 s 99200 77936 100000 78056 6 io_ibus_addr[14]
port 111 nsew signal output
rlabel metal3 s 99200 79160 100000 79280 6 io_ibus_addr[15]
port 112 nsew signal output
rlabel metal3 s 99200 80248 100000 80368 6 io_ibus_addr[16]
port 113 nsew signal output
rlabel metal3 s 99200 81472 100000 81592 6 io_ibus_addr[17]
port 114 nsew signal output
rlabel metal3 s 99200 82696 100000 82816 6 io_ibus_addr[18]
port 115 nsew signal output
rlabel metal3 s 99200 83784 100000 83904 6 io_ibus_addr[19]
port 116 nsew signal output
rlabel metal3 s 99200 62704 100000 62824 6 io_ibus_addr[1]
port 117 nsew signal output
rlabel metal3 s 99200 85008 100000 85128 6 io_ibus_addr[20]
port 118 nsew signal output
rlabel metal3 s 99200 86096 100000 86216 6 io_ibus_addr[21]
port 119 nsew signal output
rlabel metal3 s 99200 87320 100000 87440 6 io_ibus_addr[22]
port 120 nsew signal output
rlabel metal3 s 99200 88544 100000 88664 6 io_ibus_addr[23]
port 121 nsew signal output
rlabel metal3 s 99200 89632 100000 89752 6 io_ibus_addr[24]
port 122 nsew signal output
rlabel metal3 s 99200 90856 100000 90976 6 io_ibus_addr[25]
port 123 nsew signal output
rlabel metal3 s 99200 91944 100000 92064 6 io_ibus_addr[26]
port 124 nsew signal output
rlabel metal3 s 99200 93168 100000 93288 6 io_ibus_addr[27]
port 125 nsew signal output
rlabel metal3 s 99200 94392 100000 94512 6 io_ibus_addr[28]
port 126 nsew signal output
rlabel metal3 s 99200 95480 100000 95600 6 io_ibus_addr[29]
port 127 nsew signal output
rlabel metal3 s 99200 63928 100000 64048 6 io_ibus_addr[2]
port 128 nsew signal output
rlabel metal3 s 99200 96704 100000 96824 6 io_ibus_addr[30]
port 129 nsew signal output
rlabel metal3 s 99200 97792 100000 97912 6 io_ibus_addr[31]
port 130 nsew signal output
rlabel metal3 s 99200 65152 100000 65272 6 io_ibus_addr[3]
port 131 nsew signal output
rlabel metal3 s 99200 66240 100000 66360 6 io_ibus_addr[4]
port 132 nsew signal output
rlabel metal3 s 99200 67464 100000 67584 6 io_ibus_addr[5]
port 133 nsew signal output
rlabel metal3 s 99200 68552 100000 68672 6 io_ibus_addr[6]
port 134 nsew signal output
rlabel metal3 s 99200 69776 100000 69896 6 io_ibus_addr[7]
port 135 nsew signal output
rlabel metal3 s 99200 71000 100000 71120 6 io_ibus_addr[8]
port 136 nsew signal output
rlabel metal3 s 99200 72088 100000 72208 6 io_ibus_addr[9]
port 137 nsew signal output
rlabel metal3 s 99200 62160 100000 62280 6 io_ibus_inst[0]
port 138 nsew signal input
rlabel metal3 s 99200 73856 100000 73976 6 io_ibus_inst[10]
port 139 nsew signal input
rlabel metal3 s 99200 75080 100000 75200 6 io_ibus_inst[11]
port 140 nsew signal input
rlabel metal3 s 99200 76168 100000 76288 6 io_ibus_inst[12]
port 141 nsew signal input
rlabel metal3 s 99200 77392 100000 77512 6 io_ibus_inst[13]
port 142 nsew signal input
rlabel metal3 s 99200 78480 100000 78600 6 io_ibus_inst[14]
port 143 nsew signal input
rlabel metal3 s 99200 79704 100000 79824 6 io_ibus_inst[15]
port 144 nsew signal input
rlabel metal3 s 99200 80928 100000 81048 6 io_ibus_inst[16]
port 145 nsew signal input
rlabel metal3 s 99200 82016 100000 82136 6 io_ibus_inst[17]
port 146 nsew signal input
rlabel metal3 s 99200 83240 100000 83360 6 io_ibus_inst[18]
port 147 nsew signal input
rlabel metal3 s 99200 84328 100000 84448 6 io_ibus_inst[19]
port 148 nsew signal input
rlabel metal3 s 99200 63384 100000 63504 6 io_ibus_inst[1]
port 149 nsew signal input
rlabel metal3 s 99200 85552 100000 85672 6 io_ibus_inst[20]
port 150 nsew signal input
rlabel metal3 s 99200 86776 100000 86896 6 io_ibus_inst[21]
port 151 nsew signal input
rlabel metal3 s 99200 87864 100000 87984 6 io_ibus_inst[22]
port 152 nsew signal input
rlabel metal3 s 99200 89088 100000 89208 6 io_ibus_inst[23]
port 153 nsew signal input
rlabel metal3 s 99200 90176 100000 90296 6 io_ibus_inst[24]
port 154 nsew signal input
rlabel metal3 s 99200 91400 100000 91520 6 io_ibus_inst[25]
port 155 nsew signal input
rlabel metal3 s 99200 92624 100000 92744 6 io_ibus_inst[26]
port 156 nsew signal input
rlabel metal3 s 99200 93712 100000 93832 6 io_ibus_inst[27]
port 157 nsew signal input
rlabel metal3 s 99200 94936 100000 95056 6 io_ibus_inst[28]
port 158 nsew signal input
rlabel metal3 s 99200 96024 100000 96144 6 io_ibus_inst[29]
port 159 nsew signal input
rlabel metal3 s 99200 64472 100000 64592 6 io_ibus_inst[2]
port 160 nsew signal input
rlabel metal3 s 99200 97248 100000 97368 6 io_ibus_inst[30]
port 161 nsew signal input
rlabel metal3 s 99200 98472 100000 98592 6 io_ibus_inst[31]
port 162 nsew signal input
rlabel metal3 s 99200 65696 100000 65816 6 io_ibus_inst[3]
port 163 nsew signal input
rlabel metal3 s 99200 66920 100000 67040 6 io_ibus_inst[4]
port 164 nsew signal input
rlabel metal3 s 99200 68008 100000 68128 6 io_ibus_inst[5]
port 165 nsew signal input
rlabel metal3 s 99200 69232 100000 69352 6 io_ibus_inst[6]
port 166 nsew signal input
rlabel metal3 s 99200 70320 100000 70440 6 io_ibus_inst[7]
port 167 nsew signal input
rlabel metal3 s 99200 71544 100000 71664 6 io_ibus_inst[8]
port 168 nsew signal input
rlabel metal3 s 99200 72632 100000 72752 6 io_ibus_inst[9]
port 169 nsew signal input
rlabel metal3 s 99200 61072 100000 61192 6 io_ibus_valid
port 170 nsew signal input
rlabel metal2 s 49974 99200 50030 100000 6 io_irq_motor_irq
port 171 nsew signal input
rlabel metal3 s 99200 99016 100000 99136 6 io_irq_spi_irq
port 172 nsew signal input
rlabel metal3 s 99200 99560 100000 99680 6 io_irq_uart_irq
port 173 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 reset
port 174 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 175 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 175 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 175 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 175 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 176 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 176 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 176 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35273096
string GDS_FILE /home/ali11-2000/FYP/mpw/UETRV-ECORE/openlane/Core/runs/Core/results/finishing/Core.magic.gds
string GDS_START 1362456
<< end >>

