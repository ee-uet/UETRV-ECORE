magic
tech sky130A
magscale 1 2
timestamp 1647604492
<< viali >>
rect 2053 27557 2087 27591
rect 3341 27557 3375 27591
rect 6377 27557 6411 27591
rect 12357 27557 12391 27591
rect 14289 27557 14323 27591
rect 15117 27557 15151 27591
rect 16865 27557 16899 27591
rect 19257 27557 19291 27591
rect 20361 27557 20395 27591
rect 21833 27557 21867 27591
rect 24961 27557 24995 27591
rect 26525 27557 26559 27591
rect 28089 27557 28123 27591
rect 19809 27489 19843 27523
rect 1409 27421 1443 27455
rect 4077 27421 4111 27455
rect 14105 27421 14139 27455
rect 14933 27421 14967 27455
rect 16681 27421 16715 27455
rect 18153 27421 18187 27455
rect 19993 27421 20027 27455
rect 20085 27421 20119 27455
rect 25329 27421 25363 27455
rect 27261 27421 27295 27455
rect 27905 27421 27939 27455
rect 4445 27353 4479 27387
rect 25697 27353 25731 27387
rect 1593 27285 1627 27319
rect 17969 27285 18003 27319
rect 19809 27285 19843 27319
rect 27353 27285 27387 27319
rect 1869 27081 1903 27115
rect 14657 27081 14691 27115
rect 16313 27081 16347 27115
rect 20821 27081 20855 27115
rect 21465 27081 21499 27115
rect 24041 27081 24075 27115
rect 26617 27081 26651 27115
rect 15200 27013 15234 27047
rect 17776 27013 17810 27047
rect 20300 27013 20334 27047
rect 22946 27013 22980 27047
rect 24501 27013 24535 27047
rect 1409 26945 1443 26979
rect 13277 26945 13311 26979
rect 13544 26945 13578 26979
rect 14933 26945 14967 26979
rect 21005 26945 21039 26979
rect 21281 26945 21315 26979
rect 25504 26945 25538 26979
rect 26985 26945 27019 26979
rect 27241 26945 27275 26979
rect 17509 26877 17543 26911
rect 20545 26877 20579 26911
rect 23213 26877 23247 26911
rect 25237 26877 25271 26911
rect 19165 26809 19199 26843
rect 24685 26809 24719 26843
rect 18889 26741 18923 26775
rect 21833 26741 21867 26775
rect 28365 26741 28399 26775
rect 18061 26537 18095 26571
rect 18245 26537 18279 26571
rect 19349 26537 19383 26571
rect 20269 26537 20303 26571
rect 20453 26537 20487 26571
rect 21465 26537 21499 26571
rect 21925 26537 21959 26571
rect 28181 26537 28215 26571
rect 21741 26469 21775 26503
rect 1685 26333 1719 26367
rect 2145 26333 2179 26367
rect 16129 26333 16163 26367
rect 19533 26333 19567 26367
rect 19809 26333 19843 26367
rect 21005 26333 21039 26367
rect 21281 26333 21315 26367
rect 28365 26333 28399 26367
rect 1869 26265 1903 26299
rect 16396 26265 16430 26299
rect 18229 26265 18263 26299
rect 18429 26265 18463 26299
rect 20085 26265 20119 26299
rect 20285 26265 20319 26299
rect 22109 26265 22143 26299
rect 25145 26265 25179 26299
rect 26801 26265 26835 26299
rect 17509 26197 17543 26231
rect 19717 26197 19751 26231
rect 21097 26197 21131 26231
rect 21909 26197 21943 26231
rect 16681 25993 16715 26027
rect 18337 25993 18371 26027
rect 22569 25993 22603 26027
rect 16313 25925 16347 25959
rect 19257 25925 19291 25959
rect 19457 25925 19491 25959
rect 22293 25925 22327 25959
rect 25697 25925 25731 25959
rect 15485 25857 15519 25891
rect 16957 25857 16991 25891
rect 17049 25857 17083 25891
rect 17141 25857 17175 25891
rect 17325 25857 17359 25891
rect 17601 25857 17635 25891
rect 17785 25857 17819 25891
rect 18602 25857 18636 25891
rect 18706 25857 18740 25891
rect 20085 25857 20119 25891
rect 21833 25857 21867 25891
rect 21925 25857 21959 25891
rect 22109 25857 22143 25891
rect 22569 25857 22603 25891
rect 22753 25857 22787 25891
rect 23756 25857 23790 25891
rect 25421 25857 25455 25891
rect 25605 25857 25639 25891
rect 25789 25857 25823 25891
rect 18521 25789 18555 25823
rect 18797 25789 18831 25823
rect 19901 25789 19935 25823
rect 20453 25789 20487 25823
rect 20729 25789 20763 25823
rect 23489 25789 23523 25823
rect 19625 25721 19659 25755
rect 15301 25653 15335 25687
rect 17601 25653 17635 25687
rect 19441 25653 19475 25687
rect 24869 25653 24903 25687
rect 25973 25653 26007 25687
rect 17141 25449 17175 25483
rect 17233 25449 17267 25483
rect 23857 25449 23891 25483
rect 25789 25449 25823 25483
rect 16589 25381 16623 25415
rect 22017 25381 22051 25415
rect 14841 25313 14875 25347
rect 16497 25313 16531 25347
rect 17785 25313 17819 25347
rect 20361 25313 20395 25347
rect 20453 25313 20487 25347
rect 20821 25313 20855 25347
rect 24961 25313 24995 25347
rect 16681 25245 16715 25279
rect 16773 25245 16807 25279
rect 17049 25245 17083 25279
rect 17371 25245 17405 25279
rect 17509 25245 17543 25279
rect 19441 25245 19475 25279
rect 19717 25245 19751 25279
rect 20545 25245 20579 25279
rect 20637 25245 20671 25279
rect 21097 25245 21131 25279
rect 21281 25245 21315 25279
rect 21373 25245 21407 25279
rect 21465 25245 21499 25279
rect 23397 25245 23431 25279
rect 24041 25245 24075 25279
rect 24869 25245 24903 25279
rect 27169 25245 27203 25279
rect 15108 25177 15142 25211
rect 19625 25177 19659 25211
rect 21741 25177 21775 25211
rect 23130 25177 23164 25211
rect 24777 25177 24811 25211
rect 26902 25177 26936 25211
rect 16221 25109 16255 25143
rect 18015 25109 18049 25143
rect 19257 25109 19291 25143
rect 24409 25109 24443 25143
rect 15853 24905 15887 24939
rect 19073 24905 19107 24939
rect 19717 24905 19751 24939
rect 20085 24905 20119 24939
rect 21281 24905 21315 24939
rect 22569 24905 22603 24939
rect 25513 24905 25547 24939
rect 16021 24837 16055 24871
rect 16221 24837 16255 24871
rect 18889 24837 18923 24871
rect 23029 24837 23063 24871
rect 28089 24837 28123 24871
rect 15025 24769 15059 24803
rect 17141 24769 17175 24803
rect 19165 24769 19199 24803
rect 19809 24769 19843 24803
rect 19901 24769 19935 24803
rect 20545 24769 20579 24803
rect 20637 24769 20671 24803
rect 21373 24769 21407 24803
rect 22201 24769 22235 24803
rect 22477 24769 22511 24803
rect 22661 24769 22695 24803
rect 23581 24769 23615 24803
rect 23765 24769 23799 24803
rect 25145 24769 25179 24803
rect 27813 24769 27847 24803
rect 28273 24769 28307 24803
rect 15301 24701 15335 24735
rect 16865 24701 16899 24735
rect 16957 24701 16991 24735
rect 17049 24701 17083 24735
rect 18337 24701 18371 24735
rect 18613 24701 18647 24735
rect 20361 24701 20395 24735
rect 22109 24701 22143 24735
rect 25053 24701 25087 24735
rect 19533 24633 19567 24667
rect 15117 24565 15151 24599
rect 15209 24565 15243 24599
rect 16037 24565 16071 24599
rect 16681 24565 16715 24599
rect 18889 24565 18923 24599
rect 20453 24565 20487 24599
rect 21833 24565 21867 24599
rect 22017 24565 22051 24599
rect 23673 24565 23707 24599
rect 13737 24361 13771 24395
rect 16037 24361 16071 24395
rect 16221 24361 16255 24395
rect 18153 24361 18187 24395
rect 18613 24361 18647 24395
rect 21557 24361 21591 24395
rect 24961 24361 24995 24395
rect 25605 24361 25639 24395
rect 26065 24361 26099 24395
rect 24041 24293 24075 24327
rect 16497 24225 16531 24259
rect 19717 24225 19751 24259
rect 20729 24225 20763 24259
rect 24777 24225 24811 24259
rect 25513 24225 25547 24259
rect 12357 24157 12391 24191
rect 14933 24157 14967 24191
rect 15209 24157 15243 24191
rect 16773 24157 16807 24191
rect 18521 24157 18555 24191
rect 18889 24157 18923 24191
rect 19441 24157 19475 24191
rect 20545 24157 20579 24191
rect 20913 24157 20947 24191
rect 21281 24157 21315 24191
rect 22017 24157 22051 24191
rect 22201 24157 22235 24191
rect 22661 24157 22695 24191
rect 24685 24157 24719 24191
rect 24961 24157 24995 24191
rect 25605 24157 25639 24191
rect 26065 24157 26099 24191
rect 26249 24157 26283 24191
rect 12624 24089 12658 24123
rect 15117 24089 15151 24123
rect 15853 24089 15887 24123
rect 16069 24089 16103 24123
rect 17601 24089 17635 24123
rect 17785 24089 17819 24123
rect 17877 24089 17911 24123
rect 18429 24089 18463 24123
rect 18797 24089 18831 24123
rect 22928 24089 22962 24123
rect 24593 24089 24627 24123
rect 25329 24089 25363 24123
rect 14749 24021 14783 24055
rect 15485 24021 15519 24055
rect 17969 24021 18003 24055
rect 22109 24021 22143 24055
rect 25789 24021 25823 24055
rect 23305 23817 23339 23851
rect 26617 23817 26651 23851
rect 20913 23749 20947 23783
rect 24685 23749 24719 23783
rect 24869 23749 24903 23783
rect 14473 23681 14507 23715
rect 14657 23681 14691 23715
rect 14749 23681 14783 23715
rect 14841 23681 14875 23715
rect 15393 23681 15427 23715
rect 15577 23681 15611 23715
rect 15669 23681 15703 23715
rect 15761 23681 15795 23715
rect 16681 23681 16715 23715
rect 16957 23681 16991 23715
rect 18153 23681 18187 23715
rect 18420 23681 18454 23715
rect 19809 23681 19843 23715
rect 20361 23681 20395 23715
rect 20545 23681 20579 23715
rect 21005 23681 21039 23715
rect 21281 23681 21315 23715
rect 21465 23681 21499 23715
rect 22937 23681 22971 23715
rect 23397 23681 23431 23715
rect 23857 23681 23891 23715
rect 24133 23681 24167 23715
rect 25504 23681 25538 23715
rect 27813 23681 27847 23715
rect 28273 23681 28307 23715
rect 21833 23613 21867 23647
rect 22109 23613 22143 23647
rect 23673 23613 23707 23647
rect 23949 23613 23983 23647
rect 24041 23613 24075 23647
rect 25237 23613 25271 23647
rect 19533 23545 19567 23579
rect 20545 23545 20579 23579
rect 21373 23545 21407 23579
rect 23213 23545 23247 23579
rect 24501 23545 24535 23579
rect 28089 23545 28123 23579
rect 1409 23477 1443 23511
rect 15117 23477 15151 23511
rect 16037 23477 16071 23511
rect 17785 23477 17819 23511
rect 19901 23477 19935 23511
rect 23075 23477 23109 23511
rect 13001 23273 13035 23307
rect 14749 23273 14783 23307
rect 15301 23273 15335 23307
rect 18797 23273 18831 23307
rect 21097 23273 21131 23307
rect 24593 23273 24627 23307
rect 25421 23273 25455 23307
rect 17049 23205 17083 23239
rect 19533 23205 19567 23239
rect 23397 23205 23431 23239
rect 26433 23205 26467 23239
rect 15669 23137 15703 23171
rect 18245 23137 18279 23171
rect 20177 23137 20211 23171
rect 22293 23137 22327 23171
rect 25605 23137 25639 23171
rect 26065 23137 26099 23171
rect 14657 23069 14691 23103
rect 14841 23069 14875 23103
rect 15209 23069 15243 23103
rect 15393 23069 15427 23103
rect 15936 23069 15970 23103
rect 18153 23069 18187 23103
rect 20729 23069 20763 23103
rect 21741 23069 21775 23103
rect 22201 23069 22235 23103
rect 22385 23069 22419 23103
rect 23673 23069 23707 23103
rect 24961 23069 24995 23103
rect 25145 23069 25179 23103
rect 25697 23069 25731 23103
rect 25973 23069 26007 23103
rect 26341 23069 26375 23103
rect 13093 23001 13127 23035
rect 19692 23001 19726 23035
rect 20545 23001 20579 23035
rect 21925 23001 21959 23035
rect 23397 23001 23431 23035
rect 24501 23001 24535 23035
rect 18521 22933 18555 22967
rect 19809 22933 19843 22967
rect 19901 22933 19935 22967
rect 23581 22933 23615 22967
rect 25053 22933 25087 22967
rect 16221 22729 16255 22763
rect 17509 22729 17543 22763
rect 19809 22729 19843 22763
rect 23765 22729 23799 22763
rect 26157 22729 26191 22763
rect 15086 22661 15120 22695
rect 20913 22661 20947 22695
rect 24409 22661 24443 22695
rect 14309 22593 14343 22627
rect 14565 22593 14599 22627
rect 14841 22593 14875 22627
rect 17141 22593 17175 22627
rect 19441 22593 19475 22627
rect 20821 22593 20855 22627
rect 21005 22593 21039 22627
rect 21925 22593 21959 22627
rect 22192 22593 22226 22627
rect 24685 22593 24719 22627
rect 24869 22593 24903 22627
rect 25605 22593 25639 22627
rect 26065 22593 26099 22627
rect 27252 22593 27286 22627
rect 17233 22525 17267 22559
rect 19349 22525 19383 22559
rect 23949 22525 23983 22559
rect 24041 22525 24075 22559
rect 26985 22525 27019 22559
rect 23305 22457 23339 22491
rect 24685 22457 24719 22491
rect 12265 22389 12299 22423
rect 13185 22389 13219 22423
rect 25513 22389 25547 22423
rect 28365 22389 28399 22423
rect 19625 22185 19659 22219
rect 23397 22185 23431 22219
rect 23949 22185 23983 22219
rect 27261 22185 27295 22219
rect 17233 22117 17267 22151
rect 28365 22117 28399 22151
rect 14749 22049 14783 22083
rect 16957 22049 16991 22083
rect 17785 22049 17819 22083
rect 18061 22049 18095 22083
rect 25053 22049 25087 22083
rect 26065 22049 26099 22083
rect 26249 22049 26283 22083
rect 26893 22049 26927 22083
rect 1409 21981 1443 22015
rect 12173 21981 12207 22015
rect 14105 21981 14139 22015
rect 14289 21981 14323 22015
rect 15853 21981 15887 22015
rect 16865 21981 16899 22015
rect 17693 21981 17727 22015
rect 19809 21981 19843 22015
rect 19901 21981 19935 22015
rect 19993 21981 20027 22015
rect 20085 21981 20119 22015
rect 20453 21981 20487 22015
rect 23581 21981 23615 22015
rect 23673 21981 23707 22015
rect 24041 21981 24075 22015
rect 24409 21981 24443 22015
rect 24572 21975 24606 22009
rect 24685 21981 24719 22015
rect 24777 21981 24811 22015
rect 26525 21981 26559 22015
rect 26801 21981 26835 22015
rect 27077 21981 27111 22015
rect 11989 21913 12023 21947
rect 12725 21913 12759 21947
rect 12909 21913 12943 21947
rect 20720 21913 20754 21947
rect 25513 21913 25547 21947
rect 12541 21845 12575 21879
rect 14473 21845 14507 21879
rect 15669 21845 15703 21879
rect 21833 21845 21867 21879
rect 25421 21845 25455 21879
rect 26433 21845 26467 21879
rect 13645 21641 13679 21675
rect 14013 21641 14047 21675
rect 19809 21641 19843 21675
rect 15108 21573 15142 21607
rect 18521 21573 18555 21607
rect 24041 21573 24075 21607
rect 25421 21573 25455 21607
rect 25605 21573 25639 21607
rect 12521 21505 12555 21539
rect 14197 21505 14231 21539
rect 14381 21505 14415 21539
rect 14841 21505 14875 21539
rect 17785 21505 17819 21539
rect 18245 21505 18279 21539
rect 18337 21505 18371 21539
rect 18613 21505 18647 21539
rect 18705 21505 18739 21539
rect 19073 21505 19107 21539
rect 19257 21505 19291 21539
rect 19349 21505 19383 21539
rect 19625 21505 19659 21539
rect 20361 21505 20395 21539
rect 20545 21505 20579 21539
rect 20637 21505 20671 21539
rect 20729 21505 20763 21539
rect 22100 21505 22134 21539
rect 23581 21505 23615 21539
rect 23765 21505 23799 21539
rect 23857 21505 23891 21539
rect 24317 21505 24351 21539
rect 24961 21505 24995 21539
rect 25145 21505 25179 21539
rect 26433 21505 26467 21539
rect 12265 21437 12299 21471
rect 14473 21437 14507 21471
rect 18797 21437 18831 21471
rect 19441 21437 19475 21471
rect 21833 21437 21867 21471
rect 24409 21437 24443 21471
rect 21005 21369 21039 21403
rect 23673 21369 23707 21403
rect 24961 21369 24995 21403
rect 16221 21301 16255 21335
rect 17601 21301 17635 21335
rect 23213 21301 23247 21335
rect 24317 21301 24351 21335
rect 24685 21301 24719 21335
rect 26341 21301 26375 21335
rect 28365 21301 28399 21335
rect 12173 21097 12207 21131
rect 15761 21097 15795 21131
rect 22293 21097 22327 21131
rect 22661 21097 22695 21131
rect 24041 21097 24075 21131
rect 24685 21097 24719 21131
rect 11897 21029 11931 21063
rect 13553 21029 13587 21063
rect 17141 21029 17175 21063
rect 18889 21029 18923 21063
rect 21281 21029 21315 21063
rect 22753 21029 22787 21063
rect 23397 21029 23431 21063
rect 26709 21029 26743 21063
rect 15025 20961 15059 20995
rect 22845 20961 22879 20995
rect 25237 20961 25271 20995
rect 25697 20961 25731 20995
rect 25789 20961 25823 20995
rect 26157 20961 26191 20995
rect 12449 20893 12483 20927
rect 12541 20893 12575 20927
rect 12633 20893 12667 20927
rect 12817 20893 12851 20927
rect 13369 20893 13403 20927
rect 14361 20893 14395 20927
rect 14473 20893 14507 20927
rect 14565 20893 14599 20927
rect 14749 20893 14783 20927
rect 15945 20893 15979 20927
rect 16129 20893 16163 20927
rect 16405 20893 16439 20927
rect 17509 20893 17543 20927
rect 17765 20893 17799 20927
rect 19533 20893 19567 20927
rect 20637 20893 20671 20927
rect 20729 20893 20763 20927
rect 20821 20893 20855 20927
rect 21005 20893 21039 20927
rect 21649 20893 21683 20927
rect 21833 20893 21867 20927
rect 21925 20893 21959 20927
rect 22063 20893 22097 20927
rect 22569 20893 22603 20927
rect 23857 20893 23891 20927
rect 24041 20893 24075 20927
rect 24777 20893 24811 20927
rect 24869 20893 24903 20927
rect 25329 20893 25363 20927
rect 25881 20893 25915 20927
rect 25973 20893 26007 20927
rect 26433 20893 26467 20927
rect 26525 20893 26559 20927
rect 26709 20893 26743 20927
rect 26985 20893 27019 20927
rect 27241 20893 27275 20927
rect 15209 20825 15243 20859
rect 15393 20825 15427 20859
rect 23213 20825 23247 20859
rect 14105 20757 14139 20791
rect 16865 20757 16899 20791
rect 19625 20757 19659 20791
rect 20085 20757 20119 20791
rect 20361 20757 20395 20791
rect 24501 20757 24535 20791
rect 28365 20757 28399 20791
rect 12909 20553 12943 20587
rect 16313 20553 16347 20587
rect 18061 20553 18095 20587
rect 21465 20553 21499 20587
rect 26357 20553 26391 20587
rect 26525 20553 26559 20587
rect 13369 20485 13403 20519
rect 13553 20485 13587 20519
rect 14096 20485 14130 20519
rect 19809 20485 19843 20519
rect 26157 20485 26191 20519
rect 9321 20417 9355 20451
rect 11796 20417 11830 20451
rect 13829 20417 13863 20451
rect 15945 20417 15979 20451
rect 17325 20417 17359 20451
rect 17417 20417 17451 20451
rect 18245 20417 18279 20451
rect 18337 20417 18371 20451
rect 19257 20417 19291 20451
rect 19625 20417 19659 20451
rect 20352 20417 20386 20451
rect 23121 20417 23155 20451
rect 23397 20417 23431 20451
rect 24593 20417 24627 20451
rect 25329 20417 25363 20451
rect 25605 20417 25639 20451
rect 27241 20417 27275 20451
rect 9505 20349 9539 20383
rect 11529 20349 11563 20383
rect 15761 20349 15795 20383
rect 15853 20349 15887 20383
rect 17141 20349 17175 20383
rect 20085 20349 20119 20383
rect 23673 20349 23707 20383
rect 24869 20349 24903 20383
rect 25421 20349 25455 20383
rect 26985 20349 27019 20383
rect 17785 20281 17819 20315
rect 25145 20281 25179 20315
rect 9137 20213 9171 20247
rect 13185 20213 13219 20247
rect 15209 20213 15243 20247
rect 16681 20213 16715 20247
rect 18705 20213 18739 20247
rect 19165 20213 19199 20247
rect 25605 20213 25639 20247
rect 26341 20213 26375 20247
rect 28365 20213 28399 20247
rect 11805 20009 11839 20043
rect 17785 20009 17819 20043
rect 21097 20009 21131 20043
rect 22937 20009 22971 20043
rect 23397 20009 23431 20043
rect 26801 20009 26835 20043
rect 13093 19873 13127 19907
rect 19257 19873 19291 19907
rect 21741 19873 21775 19907
rect 23213 19873 23247 19907
rect 8401 19805 8435 19839
rect 8953 19805 8987 19839
rect 12061 19805 12095 19839
rect 12186 19802 12220 19836
rect 12286 19805 12320 19839
rect 12449 19805 12483 19839
rect 12725 19805 12759 19839
rect 13277 19805 13311 19839
rect 14657 19805 14691 19839
rect 14933 19805 14967 19839
rect 15209 19805 15243 19839
rect 15393 19805 15427 19839
rect 15485 19805 15519 19839
rect 15577 19805 15611 19839
rect 16405 19805 16439 19839
rect 18429 19805 18463 19839
rect 18521 19805 18555 19839
rect 18705 19805 18739 19839
rect 21465 19805 21499 19839
rect 21557 19805 21591 19839
rect 22201 19805 22235 19839
rect 22385 19805 22419 19839
rect 23489 19805 23523 19839
rect 23857 19805 23891 19839
rect 24041 19805 24075 19839
rect 24501 19805 24535 19839
rect 24685 19805 24719 19839
rect 24869 19805 24903 19839
rect 25329 19805 25363 19839
rect 25789 19805 25823 19839
rect 26065 19805 26099 19839
rect 26249 19805 26283 19839
rect 26525 19805 26559 19839
rect 28365 19805 28399 19839
rect 9198 19737 9232 19771
rect 11345 19737 11379 19771
rect 11529 19737 11563 19771
rect 15853 19737 15887 19771
rect 16672 19737 16706 19771
rect 18889 19737 18923 19771
rect 19502 19737 19536 19771
rect 22017 19737 22051 19771
rect 26801 19737 26835 19771
rect 8585 19669 8619 19703
rect 10333 19669 10367 19703
rect 13461 19669 13495 19703
rect 18153 19669 18187 19703
rect 20637 19669 20671 19703
rect 23949 19669 23983 19703
rect 24501 19669 24535 19703
rect 25421 19669 25455 19703
rect 25881 19669 25915 19703
rect 26617 19669 26651 19703
rect 9689 19465 9723 19499
rect 10057 19465 10091 19499
rect 10793 19465 10827 19499
rect 15485 19465 15519 19499
rect 18153 19465 18187 19499
rect 21373 19465 21407 19499
rect 25421 19465 25455 19499
rect 25605 19465 25639 19499
rect 14381 19397 14415 19431
rect 16313 19397 16347 19431
rect 18245 19397 18279 19431
rect 20177 19397 20211 19431
rect 21925 19397 21959 19431
rect 24593 19397 24627 19431
rect 25329 19397 25363 19431
rect 26617 19397 26651 19431
rect 27230 19397 27264 19431
rect 8493 19329 8527 19363
rect 9045 19329 9079 19363
rect 10149 19329 10183 19363
rect 11529 19329 11563 19363
rect 11713 19329 11747 19363
rect 12449 19329 12483 19363
rect 12633 19329 12667 19363
rect 14197 19329 14231 19363
rect 14841 19329 14875 19363
rect 15025 19329 15059 19363
rect 15117 19329 15151 19363
rect 15209 19329 15243 19363
rect 16129 19329 16163 19363
rect 16681 19329 16715 19363
rect 17141 19329 17175 19363
rect 17325 19329 17359 19363
rect 18705 19329 18739 19363
rect 18797 19329 18831 19363
rect 18981 19329 19015 19363
rect 19533 19329 19567 19363
rect 20545 19329 20579 19363
rect 20637 19329 20671 19363
rect 20821 19329 20855 19363
rect 21005 19329 21039 19363
rect 21281 19329 21315 19363
rect 21465 19329 21499 19363
rect 21833 19329 21867 19363
rect 22017 19329 22051 19363
rect 22385 19329 22419 19363
rect 22661 19329 22695 19363
rect 23949 19329 23983 19363
rect 25237 19329 25271 19363
rect 25605 19329 25639 19363
rect 26433 19329 26467 19363
rect 26985 19329 27019 19363
rect 8033 19261 8067 19295
rect 8861 19261 8895 19295
rect 10333 19261 10367 19295
rect 13921 19261 13955 19295
rect 14565 19261 14599 19295
rect 15945 19261 15979 19295
rect 17509 19261 17543 19295
rect 19993 19261 20027 19295
rect 24225 19261 24259 19295
rect 26157 19261 26191 19295
rect 8309 19193 8343 19227
rect 18981 19193 19015 19227
rect 24777 19193 24811 19227
rect 9229 19125 9263 19159
rect 11897 19125 11931 19159
rect 12817 19125 12851 19159
rect 13185 19125 13219 19159
rect 16865 19125 16899 19159
rect 19625 19125 19659 19159
rect 23765 19125 23799 19159
rect 24133 19125 24167 19159
rect 26249 19125 26283 19159
rect 28365 19125 28399 19159
rect 9229 18921 9263 18955
rect 11897 18921 11931 18955
rect 13737 18921 13771 18955
rect 14565 18921 14599 18955
rect 15761 18921 15795 18955
rect 16037 18921 16071 18955
rect 17049 18921 17083 18955
rect 18889 18921 18923 18955
rect 19625 18921 19659 18955
rect 22201 18921 22235 18955
rect 22385 18921 22419 18955
rect 24041 18921 24075 18955
rect 24409 18921 24443 18955
rect 25973 18921 26007 18955
rect 26249 18921 26283 18955
rect 27813 18921 27847 18955
rect 28181 18921 28215 18955
rect 20637 18853 20671 18887
rect 26893 18853 26927 18887
rect 9781 18785 9815 18819
rect 12357 18785 12391 18819
rect 14841 18785 14875 18819
rect 16589 18785 16623 18819
rect 17509 18785 17543 18819
rect 20545 18785 20579 18819
rect 22661 18785 22695 18819
rect 27445 18785 27479 18819
rect 7113 18717 7147 18751
rect 7573 18717 7607 18751
rect 9597 18717 9631 18751
rect 10517 18717 10551 18751
rect 14381 18717 14415 18751
rect 15025 18717 15059 18751
rect 15577 18717 15611 18751
rect 17233 18717 17267 18751
rect 17765 18717 17799 18751
rect 20453 18717 20487 18751
rect 20729 18717 20763 18751
rect 20913 18717 20947 18751
rect 21833 18717 21867 18751
rect 22928 18717 22962 18751
rect 24665 18717 24699 18751
rect 24790 18711 24824 18745
rect 24890 18717 24924 18751
rect 25053 18717 25087 18751
rect 25697 18717 25731 18751
rect 25973 18717 26007 18751
rect 26525 18717 26559 18751
rect 26985 18717 27019 18751
rect 27537 18717 27571 18751
rect 28089 18717 28123 18751
rect 28181 18717 28215 18751
rect 7389 18649 7423 18683
rect 10784 18649 10818 18683
rect 12624 18649 12658 18683
rect 14197 18649 14231 18683
rect 16497 18649 16531 18683
rect 19533 18649 19567 18683
rect 26709 18649 26743 18683
rect 6929 18581 6963 18615
rect 9689 18581 9723 18615
rect 15209 18581 15243 18615
rect 16405 18581 16439 18615
rect 22201 18581 22235 18615
rect 25789 18581 25823 18615
rect 26617 18581 26651 18615
rect 8033 18377 8067 18411
rect 8769 18377 8803 18411
rect 11529 18377 11563 18411
rect 13093 18377 13127 18411
rect 15669 18377 15703 18411
rect 16865 18377 16899 18411
rect 17233 18377 17267 18411
rect 17693 18377 17727 18411
rect 22937 18377 22971 18411
rect 24593 18377 24627 18411
rect 24685 18377 24719 18411
rect 6920 18309 6954 18343
rect 16773 18309 16807 18343
rect 19257 18309 19291 18343
rect 2533 18241 2567 18275
rect 8677 18241 8711 18275
rect 9505 18241 9539 18275
rect 10048 18241 10082 18275
rect 11759 18241 11793 18275
rect 11894 18241 11928 18275
rect 11994 18241 12028 18275
rect 12173 18241 12207 18275
rect 12449 18241 12483 18275
rect 12633 18241 12667 18275
rect 12728 18241 12762 18275
rect 12837 18241 12871 18275
rect 13553 18241 13587 18275
rect 13737 18241 13771 18275
rect 14381 18241 14415 18275
rect 14473 18241 14507 18275
rect 14565 18241 14599 18275
rect 14749 18241 14783 18275
rect 15025 18241 15059 18275
rect 15209 18241 15243 18275
rect 15301 18241 15335 18275
rect 15393 18241 15427 18275
rect 15945 18241 15979 18275
rect 16129 18241 16163 18275
rect 17601 18241 17635 18275
rect 18613 18241 18647 18275
rect 19533 18241 19567 18275
rect 20177 18241 20211 18275
rect 20453 18241 20487 18275
rect 21005 18241 21039 18275
rect 22109 18241 22143 18275
rect 23489 18241 23523 18275
rect 24317 18241 24351 18275
rect 24777 18241 24811 18275
rect 26157 18241 26191 18275
rect 26341 18241 26375 18275
rect 27169 18241 27203 18275
rect 28365 18241 28399 18275
rect 2789 18173 2823 18207
rect 6653 18173 6687 18207
rect 8953 18173 8987 18207
rect 9781 18173 9815 18207
rect 13829 18173 13863 18207
rect 14105 18173 14139 18207
rect 17877 18173 17911 18207
rect 19349 18173 19383 18207
rect 20269 18173 20303 18207
rect 22017 18173 22051 18207
rect 26249 18173 26283 18207
rect 26433 18173 26467 18207
rect 27077 18173 27111 18207
rect 13369 18105 13403 18139
rect 19717 18105 19751 18139
rect 20637 18105 20671 18139
rect 23305 18105 23339 18139
rect 1409 18037 1443 18071
rect 8309 18037 8343 18071
rect 9321 18037 9355 18071
rect 11161 18037 11195 18071
rect 16313 18037 16347 18071
rect 18245 18037 18279 18071
rect 19349 18037 19383 18071
rect 20177 18037 20211 18071
rect 21189 18037 21223 18071
rect 25973 18037 26007 18071
rect 28181 18037 28215 18071
rect 6929 17833 6963 17867
rect 15209 17833 15243 17867
rect 15853 17833 15887 17867
rect 18521 17833 18555 17867
rect 24409 17833 24443 17867
rect 28365 17833 28399 17867
rect 1409 17765 1443 17799
rect 22017 17765 22051 17799
rect 23121 17765 23155 17799
rect 25421 17765 25455 17799
rect 26065 17765 26099 17799
rect 11713 17697 11747 17731
rect 11989 17697 12023 17731
rect 15577 17697 15611 17731
rect 17141 17697 17175 17731
rect 19257 17697 19291 17731
rect 21465 17697 21499 17731
rect 24777 17697 24811 17731
rect 7113 17629 7147 17663
rect 7205 17629 7239 17663
rect 7941 17629 7975 17663
rect 8493 17629 8527 17663
rect 8953 17629 8987 17663
rect 9220 17629 9254 17663
rect 12265 17629 12299 17663
rect 12541 17629 12575 17663
rect 13553 17629 13587 17663
rect 13737 17629 13771 17663
rect 14381 17629 14415 17663
rect 14473 17629 14507 17663
rect 14565 17629 14599 17663
rect 14749 17629 14783 17663
rect 15117 17629 15151 17663
rect 15393 17629 15427 17663
rect 16037 17629 16071 17663
rect 16221 17629 16255 17663
rect 16313 17629 16347 17663
rect 16589 17629 16623 17663
rect 16681 17629 16715 17663
rect 19533 17629 19567 17663
rect 20545 17629 20579 17663
rect 20729 17629 20763 17663
rect 21373 17629 21407 17663
rect 22017 17629 22051 17663
rect 22201 17629 22235 17663
rect 22845 17629 22879 17663
rect 23121 17629 23155 17663
rect 24593 17629 24627 17663
rect 24685 17629 24719 17663
rect 24869 17629 24903 17663
rect 25237 17629 25271 17663
rect 25789 17629 25823 17663
rect 25881 17629 25915 17663
rect 26341 17629 26375 17663
rect 26525 17629 26559 17663
rect 26985 17629 27019 17663
rect 27241 17629 27275 17663
rect 16865 17561 16899 17595
rect 17386 17561 17420 17595
rect 25329 17561 25363 17595
rect 25513 17561 25547 17595
rect 26065 17561 26099 17595
rect 7849 17493 7883 17527
rect 8401 17493 8435 17527
rect 10333 17493 10367 17527
rect 10793 17493 10827 17527
rect 13369 17493 13403 17527
rect 14105 17493 14139 17527
rect 16589 17493 16623 17527
rect 18797 17493 18831 17527
rect 20913 17493 20947 17527
rect 21741 17493 21775 17527
rect 26341 17493 26375 17527
rect 7389 17289 7423 17323
rect 11529 17289 11563 17323
rect 12449 17289 12483 17323
rect 15577 17289 15611 17323
rect 16681 17289 16715 17323
rect 19533 17289 19567 17323
rect 26985 17289 27019 17323
rect 28181 17289 28215 17323
rect 10793 17221 10827 17255
rect 13645 17221 13679 17255
rect 20269 17221 20303 17255
rect 20821 17221 20855 17255
rect 26617 17221 26651 17255
rect 27445 17221 27479 17255
rect 6009 17153 6043 17187
rect 6377 17153 6411 17187
rect 6561 17153 6595 17187
rect 6745 17153 6779 17187
rect 8668 17153 8702 17187
rect 10977 17153 11011 17187
rect 11161 17153 11195 17187
rect 11785 17153 11819 17187
rect 11894 17153 11928 17187
rect 11989 17153 12023 17187
rect 12173 17153 12207 17187
rect 12633 17153 12667 17187
rect 13093 17153 13127 17187
rect 13369 17153 13403 17187
rect 13829 17153 13863 17187
rect 14473 17153 14507 17187
rect 14657 17153 14691 17187
rect 14933 17153 14967 17187
rect 15117 17153 15151 17187
rect 15209 17153 15243 17187
rect 15301 17153 15335 17187
rect 16037 17153 16071 17187
rect 16221 17153 16255 17187
rect 16313 17153 16347 17187
rect 17049 17153 17083 17187
rect 17877 17153 17911 17187
rect 17969 17153 18003 17187
rect 19073 17153 19107 17187
rect 19349 17153 19383 17187
rect 19533 17153 19567 17187
rect 20085 17153 20119 17187
rect 20729 17153 20763 17187
rect 20913 17153 20947 17187
rect 22293 17153 22327 17187
rect 22937 17153 22971 17187
rect 23213 17153 23247 17187
rect 24593 17153 24627 17187
rect 24869 17153 24903 17187
rect 25421 17153 25455 17187
rect 26157 17153 26191 17187
rect 27813 17153 27847 17187
rect 28365 17153 28399 17187
rect 7481 17085 7515 17119
rect 7665 17085 7699 17119
rect 8401 17085 8435 17119
rect 17141 17085 17175 17119
rect 17325 17085 17359 17119
rect 19211 17085 19245 17119
rect 22201 17085 22235 17119
rect 22661 17085 22695 17119
rect 24685 17085 24719 17119
rect 24777 17085 24811 17119
rect 26249 17085 26283 17119
rect 7021 17017 7055 17051
rect 12909 17017 12943 17051
rect 13277 17017 13311 17051
rect 17693 17017 17727 17051
rect 20453 17017 20487 17051
rect 25053 17017 25087 17051
rect 27077 17017 27111 17051
rect 5825 16949 5859 16983
rect 9781 16949 9815 16983
rect 10517 16949 10551 16983
rect 14013 16949 14047 16983
rect 14289 16949 14323 16983
rect 15853 16949 15887 16983
rect 18429 16949 18463 16983
rect 18797 16949 18831 16983
rect 23305 16949 23339 16983
rect 23489 16949 23523 16983
rect 25513 16949 25547 16983
rect 25973 16949 26007 16983
rect 8953 16745 8987 16779
rect 11345 16745 11379 16779
rect 13093 16745 13127 16779
rect 13461 16745 13495 16779
rect 28273 16745 28307 16779
rect 16313 16677 16347 16711
rect 17233 16677 17267 16711
rect 20361 16677 20395 16711
rect 22017 16677 22051 16711
rect 25789 16677 25823 16711
rect 26433 16677 26467 16711
rect 2789 16609 2823 16643
rect 5733 16609 5767 16643
rect 8309 16609 8343 16643
rect 8401 16609 8435 16643
rect 9965 16609 9999 16643
rect 12817 16609 12851 16643
rect 13553 16609 13587 16643
rect 14105 16609 14139 16643
rect 17509 16609 17543 16643
rect 19257 16609 19291 16643
rect 20085 16609 20119 16643
rect 6000 16541 6034 16575
rect 9137 16541 9171 16575
rect 11851 16541 11885 16575
rect 11986 16538 12020 16572
rect 12081 16541 12115 16575
rect 12265 16541 12299 16575
rect 13277 16541 13311 16575
rect 14381 16541 14415 16575
rect 14473 16541 14507 16575
rect 14565 16541 14599 16575
rect 14749 16541 14783 16575
rect 17049 16541 17083 16575
rect 19993 16541 20027 16575
rect 21741 16541 21775 16575
rect 24409 16541 24443 16575
rect 24593 16541 24627 16575
rect 25237 16541 25271 16575
rect 26157 16541 26191 16575
rect 26249 16541 26283 16575
rect 26893 16541 26927 16575
rect 2544 16473 2578 16507
rect 10232 16473 10266 16507
rect 11621 16473 11655 16507
rect 15025 16473 15059 16507
rect 17776 16473 17810 16507
rect 19441 16473 19475 16507
rect 22017 16473 22051 16507
rect 26433 16473 26467 16507
rect 27138 16473 27172 16507
rect 1409 16405 1443 16439
rect 7113 16405 7147 16439
rect 7849 16405 7883 16439
rect 8217 16405 8251 16439
rect 18889 16405 18923 16439
rect 21833 16405 21867 16439
rect 24501 16405 24535 16439
rect 25421 16405 25455 16439
rect 8401 16201 8435 16235
rect 9965 16201 9999 16235
rect 11161 16201 11195 16235
rect 12909 16201 12943 16235
rect 16957 16201 16991 16235
rect 18521 16201 18555 16235
rect 18889 16201 18923 16235
rect 19809 16201 19843 16235
rect 21465 16201 21499 16235
rect 26249 16201 26283 16235
rect 22946 16133 22980 16167
rect 27230 16133 27264 16167
rect 1409 16065 1443 16099
rect 5641 16065 5675 16099
rect 7573 16065 7607 16099
rect 8217 16065 8251 16099
rect 9045 16065 9079 16099
rect 9873 16065 9907 16099
rect 11796 16065 11830 16099
rect 13369 16065 13403 16099
rect 13553 16065 13587 16099
rect 14657 16065 14691 16099
rect 15761 16065 15795 16099
rect 16037 16065 16071 16099
rect 17049 16065 17083 16099
rect 17877 16065 17911 16099
rect 18429 16065 18463 16099
rect 19073 16065 19107 16099
rect 19625 16065 19659 16099
rect 20637 16065 20671 16099
rect 20821 16065 20855 16099
rect 20913 16065 20947 16099
rect 21281 16065 21315 16099
rect 21465 16065 21499 16099
rect 23489 16065 23523 16099
rect 23581 16065 23615 16099
rect 23765 16065 23799 16099
rect 24041 16065 24075 16099
rect 24297 16065 24331 16099
rect 25789 16065 25823 16099
rect 25881 16065 25915 16099
rect 25973 16065 26007 16099
rect 26157 16065 26191 16099
rect 26249 16065 26283 16099
rect 26985 16065 27019 16099
rect 7389 15997 7423 16031
rect 8033 15997 8067 16031
rect 8861 15997 8895 16031
rect 10057 15997 10091 16031
rect 11529 15997 11563 16031
rect 13645 15997 13679 16031
rect 14933 15997 14967 16031
rect 16865 15997 16899 16031
rect 17693 15997 17727 16031
rect 18061 15997 18095 16031
rect 19441 15997 19475 16031
rect 23213 15997 23247 16031
rect 9505 15929 9539 15963
rect 17417 15929 17451 15963
rect 21833 15929 21867 15963
rect 23765 15929 23799 15963
rect 5457 15861 5491 15895
rect 7757 15861 7791 15895
rect 9229 15861 9263 15895
rect 10701 15861 10735 15895
rect 13185 15861 13219 15895
rect 20085 15861 20119 15895
rect 20453 15861 20487 15895
rect 25421 15861 25455 15895
rect 28365 15861 28399 15895
rect 11069 15657 11103 15691
rect 11989 15657 12023 15691
rect 15025 15657 15059 15691
rect 16037 15657 16071 15691
rect 16773 15657 16807 15691
rect 21649 15657 21683 15691
rect 24409 15657 24443 15691
rect 24869 15657 24903 15691
rect 25513 15657 25547 15691
rect 27353 15657 27387 15691
rect 11713 15589 11747 15623
rect 16405 15589 16439 15623
rect 25881 15589 25915 15623
rect 27261 15589 27295 15623
rect 5181 15521 5215 15555
rect 8585 15521 8619 15555
rect 9689 15521 9723 15555
rect 17233 15521 17267 15555
rect 18153 15521 18187 15555
rect 24685 15521 24719 15555
rect 26433 15521 26467 15555
rect 27445 15521 27479 15555
rect 5448 15453 5482 15487
rect 9137 15453 9171 15487
rect 11345 15453 11379 15487
rect 11529 15453 11563 15487
rect 12265 15453 12299 15487
rect 12357 15453 12391 15487
rect 12449 15453 12483 15487
rect 12633 15453 12667 15487
rect 13093 15453 13127 15487
rect 13186 15453 13220 15487
rect 13461 15453 13495 15487
rect 13599 15453 13633 15487
rect 14381 15453 14415 15487
rect 14565 15453 14599 15487
rect 14657 15453 14691 15487
rect 14749 15453 14783 15487
rect 15761 15453 15795 15487
rect 15853 15453 15887 15487
rect 16589 15453 16623 15487
rect 16681 15453 16715 15487
rect 17325 15453 17359 15487
rect 18061 15453 18095 15487
rect 18797 15453 18831 15487
rect 19533 15453 19567 15487
rect 19993 15453 20027 15487
rect 21833 15453 21867 15487
rect 21925 15453 21959 15487
rect 22109 15453 22143 15487
rect 22201 15453 22235 15487
rect 24961 15453 24995 15487
rect 25513 15453 25547 15487
rect 25697 15453 25731 15487
rect 26525 15453 26559 15487
rect 27169 15453 27203 15487
rect 8340 15385 8374 15419
rect 9956 15385 9990 15419
rect 13369 15385 13403 15419
rect 15485 15385 15519 15419
rect 15669 15385 15703 15419
rect 16865 15385 16899 15419
rect 17969 15385 18003 15419
rect 20260 15385 20294 15419
rect 6561 15317 6595 15351
rect 7205 15317 7239 15351
rect 8953 15317 8987 15351
rect 13737 15317 13771 15351
rect 17601 15317 17635 15351
rect 18613 15317 18647 15351
rect 19349 15317 19383 15351
rect 21373 15317 21407 15351
rect 26893 15317 26927 15351
rect 28273 15317 28307 15351
rect 11161 15113 11195 15147
rect 14013 15113 14047 15147
rect 14933 15113 14967 15147
rect 15485 15113 15519 15147
rect 17233 15113 17267 15147
rect 20361 15113 20395 15147
rect 21281 15113 21315 15147
rect 21833 15113 21867 15147
rect 22569 15113 22603 15147
rect 5549 15045 5583 15079
rect 7941 15045 7975 15079
rect 12817 15045 12851 15079
rect 15945 15045 15979 15079
rect 20177 15045 20211 15079
rect 5733 14977 5767 15011
rect 6745 14977 6779 15011
rect 8033 14977 8067 15011
rect 9413 14977 9447 15011
rect 9597 14977 9631 15011
rect 9965 14977 9999 15011
rect 10609 14977 10643 15011
rect 12081 14977 12115 15011
rect 12449 14977 12483 15011
rect 12542 14977 12576 15011
rect 12725 14977 12759 15011
rect 12914 14977 12948 15011
rect 13369 14977 13403 15011
rect 13462 14977 13496 15011
rect 13645 14977 13679 15011
rect 13737 14977 13771 15011
rect 13834 14977 13868 15011
rect 14289 14977 14323 15011
rect 14382 14977 14416 15011
rect 14565 14977 14599 15011
rect 14657 14977 14691 15011
rect 14754 14977 14788 15011
rect 16681 14977 16715 15011
rect 17049 14977 17083 15011
rect 17601 14977 17635 15011
rect 18604 14977 18638 15011
rect 20453 14977 20487 15011
rect 21281 14977 21315 15011
rect 21465 14977 21499 15011
rect 22017 14977 22051 15011
rect 22201 14977 22235 15011
rect 22661 14977 22695 15011
rect 23285 14977 23319 15011
rect 24685 14977 24719 15011
rect 24869 14977 24903 15011
rect 27252 14977 27286 15011
rect 5273 14909 5307 14943
rect 5917 14909 5951 14943
rect 6837 14909 6871 14943
rect 6929 14909 6963 14943
rect 8217 14909 8251 14943
rect 9229 14909 9263 14943
rect 15393 14909 15427 14943
rect 17509 14909 17543 14943
rect 18337 14909 18371 14943
rect 23029 14909 23063 14943
rect 25329 14909 25363 14943
rect 25605 14909 25639 14943
rect 26985 14909 27019 14943
rect 6377 14841 6411 14875
rect 7573 14841 7607 14875
rect 10425 14841 10459 14875
rect 11621 14841 11655 14875
rect 13093 14841 13127 14875
rect 15945 14841 15979 14875
rect 20177 14841 20211 14875
rect 10149 14773 10183 14807
rect 11989 14773 12023 14807
rect 15209 14773 15243 14807
rect 19717 14773 19751 14807
rect 20821 14773 20855 14807
rect 24409 14773 24443 14807
rect 24869 14773 24903 14807
rect 25053 14773 25087 14807
rect 28365 14773 28399 14807
rect 16405 14569 16439 14603
rect 18245 14569 18279 14603
rect 25329 14569 25363 14603
rect 26065 14569 26099 14603
rect 27445 14569 27479 14603
rect 13277 14501 13311 14535
rect 16957 14501 16991 14535
rect 20361 14501 20395 14535
rect 23673 14501 23707 14535
rect 23949 14501 23983 14535
rect 7389 14433 7423 14467
rect 9689 14433 9723 14467
rect 10241 14433 10275 14467
rect 12449 14433 12483 14467
rect 14381 14433 14415 14467
rect 18613 14433 18647 14467
rect 19625 14433 19659 14467
rect 21557 14433 21591 14467
rect 22845 14433 22879 14467
rect 25145 14433 25179 14467
rect 25973 14433 26007 14467
rect 7573 14365 7607 14399
rect 7757 14365 7791 14399
rect 8217 14365 8251 14399
rect 9965 14365 9999 14399
rect 10497 14365 10531 14399
rect 12173 14365 12207 14399
rect 14105 14365 14139 14399
rect 15485 14365 15519 14399
rect 15945 14365 15979 14399
rect 16313 14365 16347 14399
rect 16497 14365 16531 14399
rect 17138 14359 17172 14393
rect 17233 14365 17267 14399
rect 17877 14365 17911 14399
rect 18521 14365 18555 14399
rect 18705 14365 18739 14399
rect 19441 14365 19475 14399
rect 19717 14365 19751 14399
rect 19993 14365 20027 14399
rect 20177 14365 20211 14399
rect 20453 14365 20487 14399
rect 21097 14365 21131 14399
rect 21741 14365 21775 14399
rect 22017 14365 22051 14399
rect 22201 14365 22235 14399
rect 22569 14365 22603 14399
rect 22661 14365 22695 14399
rect 23208 14343 23242 14377
rect 23305 14365 23339 14399
rect 23581 14365 23615 14399
rect 23673 14365 23707 14399
rect 25053 14365 25087 14399
rect 25329 14365 25363 14399
rect 26157 14365 26191 14399
rect 26801 14365 26835 14399
rect 26985 14365 27019 14399
rect 27077 14365 27111 14399
rect 27215 14365 27249 14399
rect 27721 14365 27755 14399
rect 28089 14365 28123 14399
rect 13461 14297 13495 14331
rect 18061 14297 18095 14331
rect 23397 14297 23431 14331
rect 25881 14297 25915 14331
rect 27905 14297 27939 14331
rect 6101 14229 6135 14263
rect 8033 14229 8067 14263
rect 11621 14229 11655 14263
rect 15301 14229 15335 14263
rect 16129 14229 16163 14263
rect 19257 14229 19291 14263
rect 20821 14229 20855 14263
rect 22845 14229 22879 14263
rect 25513 14229 25547 14263
rect 26341 14229 26375 14263
rect 5273 14025 5307 14059
rect 6377 14025 6411 14059
rect 8953 14025 8987 14059
rect 9229 14025 9263 14059
rect 9597 14025 9631 14059
rect 17785 14025 17819 14059
rect 18245 14025 18279 14059
rect 20085 14025 20119 14059
rect 22569 14025 22603 14059
rect 23305 14025 23339 14059
rect 25237 14025 25271 14059
rect 27445 14025 27479 14059
rect 7840 13957 7874 13991
rect 10333 13957 10367 13991
rect 10517 13957 10551 13991
rect 15301 13957 15335 13991
rect 15485 13957 15519 13991
rect 16037 13957 16071 13991
rect 17049 13957 17083 13991
rect 18972 13957 19006 13991
rect 24409 13957 24443 13991
rect 24777 13957 24811 13991
rect 26341 13957 26375 13991
rect 5089 13889 5123 13923
rect 5549 13889 5583 13923
rect 5733 13889 5767 13923
rect 6745 13889 6779 13923
rect 9689 13889 9723 13923
rect 10977 13889 11011 13923
rect 11621 13889 11655 13923
rect 12725 13889 12759 13923
rect 13001 13889 13035 13923
rect 13094 13889 13128 13923
rect 13277 13889 13311 13923
rect 13369 13889 13403 13923
rect 13507 13889 13541 13923
rect 17417 13889 17451 13923
rect 17877 13889 17911 13923
rect 18429 13889 18463 13923
rect 18705 13889 18739 13923
rect 20453 13889 20487 13923
rect 20545 13889 20579 13923
rect 20729 13889 20763 13923
rect 20821 13889 20855 13923
rect 21281 13889 21315 13923
rect 21465 13889 21499 13923
rect 21822 13889 21856 13923
rect 22149 13889 22183 13923
rect 22937 13889 22971 13923
rect 23765 13889 23799 13923
rect 23949 13889 23983 13923
rect 24225 13889 24259 13923
rect 24501 13889 24535 13923
rect 25053 13889 25087 13923
rect 26157 13889 26191 13923
rect 26249 13889 26283 13923
rect 26525 13889 26559 13923
rect 26985 13889 27019 13923
rect 28273 13889 28307 13923
rect 5917 13821 5951 13855
rect 6837 13821 6871 13855
rect 6929 13821 6963 13855
rect 7573 13821 7607 13855
rect 9781 13821 9815 13855
rect 12449 13821 12483 13855
rect 14473 13821 14507 13855
rect 14749 13821 14783 13855
rect 15577 13821 15611 13855
rect 22017 13821 22051 13855
rect 22845 13821 22879 13855
rect 23581 13821 23615 13855
rect 24869 13821 24903 13855
rect 11161 13753 11195 13787
rect 16037 13753 16071 13787
rect 16865 13753 16899 13787
rect 28089 13753 28123 13787
rect 13645 13685 13679 13719
rect 17049 13685 17083 13719
rect 21005 13685 21039 13719
rect 21465 13685 21499 13719
rect 21833 13685 21867 13719
rect 22293 13685 22327 13719
rect 22753 13685 22787 13719
rect 24225 13685 24259 13719
rect 25053 13685 25087 13719
rect 25973 13685 26007 13719
rect 27169 13685 27203 13719
rect 7205 13481 7239 13515
rect 7665 13481 7699 13515
rect 13737 13481 13771 13515
rect 18337 13481 18371 13515
rect 21741 13481 21775 13515
rect 23857 13481 23891 13515
rect 23949 13481 23983 13515
rect 24409 13481 24443 13515
rect 24777 13481 24811 13515
rect 26433 13481 26467 13515
rect 28365 13481 28399 13515
rect 6653 13413 6687 13447
rect 16221 13413 16255 13447
rect 18705 13413 18739 13447
rect 5273 13345 5307 13379
rect 8125 13345 8159 13379
rect 8217 13345 8251 13379
rect 9045 13345 9079 13379
rect 14381 13345 14415 13379
rect 15669 13345 15703 13379
rect 17049 13345 17083 13379
rect 17233 13345 17267 13379
rect 19257 13345 19291 13379
rect 20361 13345 20395 13379
rect 22385 13345 22419 13379
rect 24041 13345 24075 13379
rect 26985 13345 27019 13379
rect 5540 13277 5574 13311
rect 8033 13277 8067 13311
rect 9229 13277 9263 13311
rect 9689 13277 9723 13311
rect 11345 13277 11379 13311
rect 13093 13277 13127 13311
rect 13186 13277 13220 13311
rect 13369 13277 13403 13311
rect 13599 13277 13633 13311
rect 14105 13277 14139 13311
rect 17141 13277 17175 13311
rect 17693 13277 17727 13311
rect 17785 13277 17819 13311
rect 17877 13277 17911 13311
rect 19533 13277 19567 13311
rect 22201 13277 22235 13311
rect 22661 13277 22695 13311
rect 22937 13277 22971 13311
rect 23765 13277 23799 13311
rect 24409 13277 24443 13311
rect 24501 13277 24535 13311
rect 26065 13277 26099 13311
rect 26249 13277 26283 13311
rect 7297 13209 7331 13243
rect 9956 13209 9990 13243
rect 11612 13209 11646 13243
rect 13461 13209 13495 13243
rect 16221 13209 16255 13243
rect 20606 13209 20640 13243
rect 25513 13209 25547 13243
rect 25697 13209 25731 13243
rect 27252 13209 27286 13243
rect 9413 13141 9447 13175
rect 11069 13141 11103 13175
rect 12725 13141 12759 13175
rect 15485 13141 15519 13175
rect 15761 13141 15795 13175
rect 16865 13141 16899 13175
rect 18061 13141 18095 13175
rect 6745 12937 6779 12971
rect 9965 12937 9999 12971
rect 10977 12937 11011 12971
rect 11529 12937 11563 12971
rect 12633 12937 12667 12971
rect 12725 12937 12759 12971
rect 14289 12937 14323 12971
rect 15209 12937 15243 12971
rect 19717 12937 19751 12971
rect 20459 12937 20493 12971
rect 21373 12937 21407 12971
rect 22569 12937 22603 12971
rect 25605 12937 25639 12971
rect 25881 12937 25915 12971
rect 28365 12937 28399 12971
rect 7389 12869 7423 12903
rect 10333 12869 10367 12903
rect 13921 12869 13955 12903
rect 14841 12869 14875 12903
rect 17417 12869 17451 12903
rect 20361 12869 20395 12903
rect 20545 12869 20579 12903
rect 21925 12869 21959 12903
rect 22477 12869 22511 12903
rect 24492 12869 24526 12903
rect 27230 12869 27264 12903
rect 4997 12801 5031 12835
rect 5457 12801 5491 12835
rect 5641 12801 5675 12835
rect 7849 12801 7883 12835
rect 8105 12801 8139 12835
rect 9689 12801 9723 12835
rect 11161 12801 11195 12835
rect 11713 12801 11747 12835
rect 13645 12801 13679 12835
rect 13738 12801 13772 12835
rect 14013 12801 14047 12835
rect 14110 12801 14144 12835
rect 14565 12801 14599 12835
rect 14658 12801 14692 12835
rect 14933 12801 14967 12835
rect 15071 12801 15105 12835
rect 15669 12801 15703 12835
rect 15853 12801 15887 12835
rect 16313 12801 16347 12835
rect 16865 12801 16899 12835
rect 17877 12801 17911 12835
rect 18705 12801 18739 12835
rect 19165 12801 19199 12835
rect 19809 12801 19843 12835
rect 20637 12801 20671 12835
rect 20913 12801 20947 12835
rect 21097 12801 21131 12835
rect 21833 12801 21867 12835
rect 22017 12801 22051 12835
rect 24225 12801 24259 12835
rect 5825 12733 5859 12767
rect 6837 12733 6871 12767
rect 6929 12733 6963 12767
rect 10425 12733 10459 12767
rect 10609 12733 10643 12767
rect 11989 12733 12023 12767
rect 12909 12733 12943 12767
rect 15761 12733 15795 12767
rect 16957 12733 16991 12767
rect 17969 12733 18003 12767
rect 18981 12733 19015 12767
rect 22937 12733 22971 12767
rect 23213 12733 23247 12767
rect 26985 12733 27019 12767
rect 6377 12665 6411 12699
rect 9229 12665 9263 12699
rect 9505 12665 9539 12699
rect 16681 12665 16715 12699
rect 17417 12665 17451 12699
rect 18521 12665 18555 12699
rect 19349 12665 19383 12699
rect 5181 12597 5215 12631
rect 11897 12597 11931 12631
rect 12265 12597 12299 12631
rect 13277 12597 13311 12631
rect 16129 12597 16163 12631
rect 18061 12597 18095 12631
rect 18245 12597 18279 12631
rect 20913 12597 20947 12631
rect 13645 12393 13679 12427
rect 16405 12393 16439 12427
rect 18153 12393 18187 12427
rect 18797 12393 18831 12427
rect 21097 12393 21131 12427
rect 22109 12393 22143 12427
rect 27261 12393 27295 12427
rect 6561 12325 6595 12359
rect 8953 12325 8987 12359
rect 10241 12325 10275 12359
rect 20637 12325 20671 12359
rect 22477 12325 22511 12359
rect 24409 12325 24443 12359
rect 25789 12325 25823 12359
rect 5181 12257 5215 12291
rect 7389 12257 7423 12291
rect 9505 12257 9539 12291
rect 10885 12257 10919 12291
rect 13093 12257 13127 12291
rect 14105 12257 14139 12291
rect 15301 12257 15335 12291
rect 16195 12257 16229 12291
rect 16957 12257 16991 12291
rect 18153 12257 18187 12291
rect 25973 12257 26007 12291
rect 26249 12257 26283 12291
rect 28365 12257 28399 12291
rect 5437 12189 5471 12223
rect 8125 12189 8159 12223
rect 8309 12189 8343 12223
rect 9321 12189 9355 12223
rect 11069 12189 11103 12223
rect 11897 12189 11931 12223
rect 11989 12189 12023 12223
rect 14289 12189 14323 12223
rect 16037 12189 16071 12223
rect 16405 12189 16439 12223
rect 16589 12189 16623 12223
rect 17233 12189 17267 12223
rect 18337 12189 18371 12223
rect 19257 12189 19291 12223
rect 21741 12189 21775 12223
rect 21925 12189 21959 12223
rect 22201 12189 22235 12223
rect 22615 12189 22649 12223
rect 23028 12189 23062 12223
rect 23121 12189 23155 12223
rect 23397 12189 23431 12223
rect 23581 12189 23615 12223
rect 24685 12189 24719 12223
rect 25697 12189 25731 12223
rect 27077 12189 27111 12223
rect 7205 12121 7239 12155
rect 9413 12121 9447 12155
rect 10057 12121 10091 12155
rect 13553 12121 13587 12155
rect 14473 12121 14507 12155
rect 15117 12121 15151 12155
rect 18061 12121 18095 12155
rect 19524 12121 19558 12155
rect 20913 12121 20947 12155
rect 21129 12121 21163 12155
rect 22753 12121 22787 12155
rect 22845 12121 22879 12155
rect 24409 12121 24443 12155
rect 25053 12121 25087 12155
rect 25237 12121 25271 12155
rect 6837 12053 6871 12087
rect 7297 12053 7331 12087
rect 7941 12053 7975 12087
rect 10517 12053 10551 12087
rect 11529 12053 11563 12087
rect 12173 12053 12207 12087
rect 12449 12053 12483 12087
rect 12817 12053 12851 12087
rect 12909 12053 12943 12087
rect 14749 12053 14783 12087
rect 15209 12053 15243 12087
rect 18521 12053 18555 12087
rect 21281 12053 21315 12087
rect 21557 12053 21591 12087
rect 23489 12053 23523 12087
rect 23857 12053 23891 12087
rect 24593 12053 24627 12087
rect 25697 12053 25731 12087
rect 6009 11849 6043 11883
rect 7941 11849 7975 11883
rect 11529 11849 11563 11883
rect 15669 11849 15703 11883
rect 16313 11849 16347 11883
rect 16681 11849 16715 11883
rect 19257 11849 19291 11883
rect 24501 11849 24535 11883
rect 9413 11781 9447 11815
rect 18705 11781 18739 11815
rect 21925 11781 21959 11815
rect 22109 11781 22143 11815
rect 6469 11713 6503 11747
rect 6653 11713 6687 11747
rect 6837 11713 6871 11747
rect 7113 11713 7147 11747
rect 7757 11713 7791 11747
rect 8585 11713 8619 11747
rect 10037 11713 10071 11747
rect 12164 11713 12198 11747
rect 13553 11713 13587 11747
rect 14289 11713 14323 11747
rect 14556 11713 14590 11747
rect 16129 11713 16163 11747
rect 16313 11713 16347 11747
rect 17693 11713 17727 11747
rect 18521 11713 18555 11747
rect 19441 11713 19475 11747
rect 19901 11713 19935 11747
rect 21005 11713 21039 11747
rect 21465 11713 21499 11747
rect 22569 11713 22603 11747
rect 22845 11713 22879 11747
rect 23029 11713 23063 11747
rect 23581 11713 23615 11747
rect 24593 11713 24627 11747
rect 25513 11713 25547 11747
rect 8677 11645 8711 11679
rect 8769 11645 8803 11679
rect 9781 11645 9815 11679
rect 11897 11645 11931 11679
rect 17141 11645 17175 11679
rect 17417 11645 17451 11679
rect 21373 11645 21407 11679
rect 22753 11645 22787 11679
rect 23673 11645 23707 11679
rect 24225 11645 24259 11679
rect 25421 11645 25455 11679
rect 25881 11645 25915 11679
rect 9229 11577 9263 11611
rect 16773 11577 16807 11611
rect 19717 11577 19751 11611
rect 22661 11577 22695 11611
rect 24317 11577 24351 11611
rect 7297 11509 7331 11543
rect 8217 11509 8251 11543
rect 11161 11509 11195 11543
rect 13277 11509 13311 11543
rect 13645 11509 13679 11543
rect 14013 11509 14047 11543
rect 18797 11509 18831 11543
rect 20269 11509 20303 11543
rect 20821 11509 20855 11543
rect 22385 11509 22419 11543
rect 23581 11509 23615 11543
rect 23949 11509 23983 11543
rect 24409 11509 24443 11543
rect 6285 11305 6319 11339
rect 8953 11305 8987 11339
rect 14841 11305 14875 11339
rect 17233 11305 17267 11339
rect 17969 11305 18003 11339
rect 22017 11305 22051 11339
rect 22293 11305 22327 11339
rect 23121 11305 23155 11339
rect 23397 11305 23431 11339
rect 23949 11305 23983 11339
rect 24685 11305 24719 11339
rect 25973 11305 26007 11339
rect 9505 11237 9539 11271
rect 10517 11237 10551 11271
rect 13369 11237 13403 11271
rect 16221 11237 16255 11271
rect 16681 11237 16715 11271
rect 19349 11237 19383 11271
rect 24777 11237 24811 11271
rect 7665 11169 7699 11203
rect 11161 11169 11195 11203
rect 12817 11169 12851 11203
rect 18613 11169 18647 11203
rect 23397 11169 23431 11203
rect 24593 11169 24627 11203
rect 1409 11101 1443 11135
rect 7398 11101 7432 11135
rect 8033 11101 8067 11135
rect 8217 11101 8251 11135
rect 9321 11101 9355 11135
rect 9781 11101 9815 11135
rect 9965 11101 9999 11135
rect 10057 11101 10091 11135
rect 10885 11101 10919 11135
rect 12081 11101 12115 11135
rect 12357 11101 12391 11135
rect 13001 11101 13035 11135
rect 13553 11101 13587 11135
rect 14197 11101 14231 11135
rect 14381 11101 14415 11135
rect 14473 11101 14507 11135
rect 14565 11101 14599 11135
rect 15301 11101 15335 11135
rect 15394 11101 15428 11135
rect 15669 11101 15703 11135
rect 15766 11101 15800 11135
rect 18245 11101 18279 11135
rect 18429 11101 18463 11135
rect 19717 11101 19751 11135
rect 20637 11101 20671 11135
rect 20904 11101 20938 11135
rect 22661 11101 22695 11135
rect 22845 11101 22879 11135
rect 23673 11101 23707 11135
rect 24869 11101 24903 11135
rect 27353 11101 27387 11135
rect 28365 11101 28399 11135
rect 8401 11033 8435 11067
rect 15577 11033 15611 11067
rect 17417 11033 17451 11067
rect 17601 11033 17635 11067
rect 19901 11033 19935 11067
rect 20085 11033 20119 11067
rect 22753 11033 22787 11067
rect 25145 11033 25179 11067
rect 25329 11033 25363 11067
rect 27086 11033 27120 11067
rect 10977 10965 11011 10999
rect 15945 10965 15979 10999
rect 9229 10761 9263 10795
rect 10333 10761 10367 10795
rect 16865 10761 16899 10795
rect 23305 10761 23339 10795
rect 25421 10761 25455 10795
rect 27261 10761 27295 10795
rect 11069 10693 11103 10727
rect 12081 10693 12115 10727
rect 12265 10693 12299 10727
rect 17509 10693 17543 10727
rect 22192 10693 22226 10727
rect 26157 10693 26191 10727
rect 26341 10693 26375 10727
rect 7849 10625 7883 10659
rect 8116 10625 8150 10659
rect 9781 10625 9815 10659
rect 11713 10625 11747 10659
rect 12725 10625 12759 10659
rect 13185 10625 13219 10659
rect 14013 10625 14047 10659
rect 14105 10625 14139 10659
rect 15025 10625 15059 10659
rect 15669 10625 15703 10659
rect 16681 10625 16715 10659
rect 17693 10625 17727 10659
rect 19082 10625 19116 10659
rect 20260 10625 20294 10659
rect 24041 10625 24075 10659
rect 24308 10625 24342 10659
rect 25973 10625 26007 10659
rect 27353 10625 27387 10659
rect 27905 10625 27939 10659
rect 9965 10557 9999 10591
rect 13001 10557 13035 10591
rect 13369 10557 13403 10591
rect 14197 10557 14231 10591
rect 15761 10557 15795 10591
rect 15945 10557 15979 10591
rect 19349 10557 19383 10591
rect 19993 10557 20027 10591
rect 21925 10557 21959 10591
rect 10793 10489 10827 10523
rect 12541 10489 12575 10523
rect 13645 10489 13679 10523
rect 9597 10421 9631 10455
rect 11529 10421 11563 10455
rect 15301 10421 15335 10455
rect 17325 10421 17359 10455
rect 17969 10421 18003 10455
rect 19625 10421 19659 10455
rect 21373 10421 21407 10455
rect 27721 10421 27755 10455
rect 12541 10217 12575 10251
rect 14841 10217 14875 10251
rect 15577 10217 15611 10251
rect 16037 10217 16071 10251
rect 17693 10217 17727 10251
rect 18889 10217 18923 10251
rect 19625 10217 19659 10251
rect 20637 10217 20671 10251
rect 25789 10217 25823 10251
rect 8217 10081 8251 10115
rect 9321 10081 9355 10115
rect 11161 10081 11195 10115
rect 13369 10081 13403 10115
rect 15209 10081 15243 10115
rect 17417 10081 17451 10115
rect 18337 10081 18371 10115
rect 20085 10081 20119 10115
rect 20177 10081 20211 10115
rect 21557 10081 21591 10115
rect 22753 10081 22787 10115
rect 26341 10081 26375 10115
rect 1869 10013 1903 10047
rect 8401 10013 8435 10047
rect 11428 10013 11462 10047
rect 13277 10013 13311 10047
rect 14197 10013 14231 10047
rect 14290 10013 14324 10047
rect 14565 10013 14599 10047
rect 14703 10013 14737 10047
rect 15393 10013 15427 10047
rect 17150 10013 17184 10047
rect 18705 10013 18739 10047
rect 19993 10013 20027 10047
rect 20821 10013 20855 10047
rect 21097 10013 21131 10047
rect 23765 10013 23799 10047
rect 25329 10013 25363 10047
rect 26801 10013 26835 10047
rect 27068 10013 27102 10047
rect 1685 9945 1719 9979
rect 2145 9945 2179 9979
rect 9588 9945 9622 9979
rect 14473 9945 14507 9979
rect 18153 9945 18187 9979
rect 23581 9945 23615 9979
rect 24685 9945 24719 9979
rect 24869 9945 24903 9979
rect 26157 9945 26191 9979
rect 10701 9877 10735 9911
rect 12817 9877 12851 9911
rect 13185 9877 13219 9911
rect 18061 9877 18095 9911
rect 19349 9877 19383 9911
rect 21281 9877 21315 9911
rect 22109 9877 22143 9911
rect 22477 9877 22511 9911
rect 22569 9877 22603 9911
rect 23949 9877 23983 9911
rect 25513 9877 25547 9911
rect 26249 9877 26283 9911
rect 28181 9877 28215 9911
rect 8585 9673 8619 9707
rect 9597 9673 9631 9707
rect 10057 9673 10091 9707
rect 10517 9673 10551 9707
rect 11529 9673 11563 9707
rect 12173 9673 12207 9707
rect 14289 9673 14323 9707
rect 15669 9673 15703 9707
rect 19073 9673 19107 9707
rect 22845 9673 22879 9707
rect 12633 9605 12667 9639
rect 13176 9605 13210 9639
rect 14565 9605 14599 9639
rect 15301 9605 15335 9639
rect 18061 9605 18095 9639
rect 18797 9605 18831 9639
rect 25412 9605 25446 9639
rect 28089 9605 28123 9639
rect 8769 9537 8803 9571
rect 9781 9537 9815 9571
rect 10425 9537 10459 9571
rect 11713 9537 11747 9571
rect 11897 9537 11931 9571
rect 16129 9537 16163 9571
rect 16221 9537 16255 9571
rect 17325 9537 17359 9571
rect 18429 9537 18463 9571
rect 18613 9537 18647 9571
rect 19441 9537 19475 9571
rect 21198 9537 21232 9571
rect 21465 9537 21499 9571
rect 22477 9537 22511 9571
rect 24602 9537 24636 9571
rect 27813 9537 27847 9571
rect 28273 9537 28307 9571
rect 10701 9469 10735 9503
rect 12909 9469 12943 9503
rect 15025 9469 15059 9503
rect 15209 9469 15243 9503
rect 19533 9469 19567 9503
rect 19717 9469 19751 9503
rect 22201 9469 22235 9503
rect 22385 9469 22419 9503
rect 24869 9469 24903 9503
rect 25145 9469 25179 9503
rect 17877 9401 17911 9435
rect 23489 9401 23523 9435
rect 26525 9401 26559 9435
rect 9229 9333 9263 9367
rect 15945 9333 15979 9367
rect 16681 9333 16715 9367
rect 17509 9333 17543 9367
rect 20085 9333 20119 9367
rect 16405 9129 16439 9163
rect 17049 9129 17083 9163
rect 18705 9129 18739 9163
rect 23305 9129 23339 9163
rect 25329 9129 25363 9163
rect 10333 9061 10367 9095
rect 22661 9061 22695 9095
rect 8953 8993 8987 9027
rect 11069 8993 11103 9027
rect 11253 8993 11287 9027
rect 13185 8993 13219 9027
rect 15025 8993 15059 9027
rect 19717 8993 19751 9027
rect 19901 8993 19935 9027
rect 23765 8993 23799 9027
rect 23949 8993 23983 9027
rect 25881 8993 25915 9027
rect 26709 8993 26743 9027
rect 8401 8925 8435 8959
rect 10977 8925 11011 8959
rect 12081 8925 12115 8959
rect 12909 8925 12943 8959
rect 13553 8925 13587 8959
rect 14105 8925 14139 8959
rect 14289 8925 14323 8959
rect 14473 8925 14507 8959
rect 16681 8925 16715 8959
rect 16865 8925 16899 8959
rect 17325 8925 17359 8959
rect 17592 8925 17626 8959
rect 21281 8925 21315 8959
rect 23673 8925 23707 8959
rect 24593 8925 24627 8959
rect 26525 8925 26559 8959
rect 9198 8857 9232 8891
rect 13001 8857 13035 8891
rect 14381 8857 14415 8891
rect 15270 8857 15304 8891
rect 20637 8857 20671 8891
rect 20821 8857 20855 8891
rect 21548 8857 21582 8891
rect 24409 8857 24443 8891
rect 25697 8857 25731 8891
rect 26341 8857 26375 8891
rect 8585 8789 8619 8823
rect 10609 8789 10643 8823
rect 11897 8789 11931 8823
rect 12541 8789 12575 8823
rect 13737 8789 13771 8823
rect 14657 8789 14691 8823
rect 19257 8789 19291 8823
rect 19993 8789 20027 8823
rect 20361 8789 20395 8823
rect 21005 8789 21039 8823
rect 25789 8789 25823 8823
rect 9413 8585 9447 8619
rect 13001 8585 13035 8619
rect 13645 8585 13679 8619
rect 14289 8585 14323 8619
rect 16865 8585 16899 8619
rect 17325 8585 17359 8619
rect 18521 8585 18555 8619
rect 19901 8585 19935 8619
rect 21833 8585 21867 8619
rect 24041 8585 24075 8619
rect 14657 8517 14691 8551
rect 15485 8517 15519 8551
rect 20913 8517 20947 8551
rect 22937 8517 22971 8551
rect 23489 8517 23523 8551
rect 25513 8517 25547 8551
rect 1409 8449 1443 8483
rect 9597 8449 9631 8483
rect 10793 8449 10827 8483
rect 10885 8449 10919 8483
rect 11621 8449 11655 8483
rect 11888 8449 11922 8483
rect 14427 8449 14461 8483
rect 14565 8449 14599 8483
rect 14785 8449 14819 8483
rect 14933 8449 14967 8483
rect 15301 8449 15335 8483
rect 16129 8449 16163 8483
rect 17233 8449 17267 8483
rect 18061 8449 18095 8483
rect 18337 8449 18371 8483
rect 19165 8449 19199 8483
rect 19809 8449 19843 8483
rect 20637 8449 20671 8483
rect 22017 8449 22051 8483
rect 23857 8449 23891 8483
rect 24685 8449 24719 8483
rect 27905 8449 27939 8483
rect 28365 8449 28399 8483
rect 9781 8381 9815 8415
rect 10149 8381 10183 8415
rect 10977 8381 11011 8415
rect 13737 8381 13771 8415
rect 13921 8381 13955 8415
rect 15945 8381 15979 8415
rect 17509 8381 17543 8415
rect 18153 8381 18187 8415
rect 20085 8381 20119 8415
rect 23305 8381 23339 8415
rect 24409 8381 24443 8415
rect 24593 8381 24627 8415
rect 25329 8381 25363 8415
rect 1593 8313 1627 8347
rect 16313 8313 16347 8347
rect 18981 8313 19015 8347
rect 25053 8313 25087 8347
rect 10425 8245 10459 8279
rect 13277 8245 13311 8279
rect 18337 8245 18371 8279
rect 19441 8245 19475 8279
rect 20453 8245 20487 8279
rect 22845 8245 22879 8279
rect 28181 8245 28215 8279
rect 12909 8041 12943 8075
rect 13461 8041 13495 8075
rect 14105 8041 14139 8075
rect 15117 8041 15151 8075
rect 20085 8041 20119 8075
rect 11529 7973 11563 8007
rect 11989 7973 12023 8007
rect 21741 7973 21775 8007
rect 24041 7973 24075 8007
rect 10149 7905 10183 7939
rect 14473 7905 14507 7939
rect 19533 7905 19567 7939
rect 20361 7905 20395 7939
rect 22661 7905 22695 7939
rect 9689 7837 9723 7871
rect 12173 7837 12207 7871
rect 12357 7837 12391 7871
rect 13001 7837 13035 7871
rect 14657 7837 14691 7871
rect 16497 7837 16531 7871
rect 16957 7837 16991 7871
rect 18889 7837 18923 7871
rect 20617 7837 20651 7871
rect 26065 7837 26099 7871
rect 26525 7837 26559 7871
rect 10394 7769 10428 7803
rect 16230 7769 16264 7803
rect 17202 7769 17236 7803
rect 19625 7769 19659 7803
rect 22906 7769 22940 7803
rect 25820 7769 25854 7803
rect 9873 7701 9907 7735
rect 14841 7701 14875 7735
rect 18337 7701 18371 7735
rect 18705 7701 18739 7735
rect 19717 7701 19751 7735
rect 24685 7701 24719 7735
rect 26341 7701 26375 7735
rect 10057 7497 10091 7531
rect 15117 7497 15151 7531
rect 16313 7497 16347 7531
rect 16957 7497 16991 7531
rect 17233 7497 17267 7531
rect 17693 7497 17727 7531
rect 22109 7497 22143 7531
rect 22845 7497 22879 7531
rect 24961 7497 24995 7531
rect 25421 7497 25455 7531
rect 22753 7429 22787 7463
rect 10241 7361 10275 7395
rect 10333 7361 10367 7395
rect 12265 7361 12299 7395
rect 12357 7361 12391 7395
rect 13369 7361 13403 7395
rect 14197 7361 14231 7395
rect 14289 7361 14323 7395
rect 15485 7361 15519 7395
rect 16129 7361 16163 7395
rect 16773 7361 16807 7395
rect 17601 7361 17635 7395
rect 18521 7361 18555 7395
rect 18788 7361 18822 7395
rect 21925 7361 21959 7395
rect 25329 7361 25363 7395
rect 27813 7361 27847 7395
rect 28365 7361 28399 7395
rect 13185 7293 13219 7327
rect 14381 7293 14415 7327
rect 15577 7293 15611 7327
rect 15669 7293 15703 7327
rect 17877 7293 17911 7327
rect 22937 7293 22971 7327
rect 25605 7293 25639 7327
rect 13829 7225 13863 7259
rect 12541 7157 12575 7191
rect 13553 7157 13587 7191
rect 19901 7157 19935 7191
rect 22385 7157 22419 7191
rect 28181 7157 28215 7191
rect 22201 6953 22235 6987
rect 14105 6817 14139 6851
rect 16957 6817 16991 6851
rect 18429 6817 18463 6851
rect 21557 6817 21591 6851
rect 22753 6817 22787 6851
rect 24869 6817 24903 6851
rect 24961 6817 24995 6851
rect 11897 6749 11931 6783
rect 13553 6749 13587 6783
rect 17877 6749 17911 6783
rect 18061 6749 18095 6783
rect 19441 6749 19475 6783
rect 21373 6749 21407 6783
rect 22569 6749 22603 6783
rect 23581 6749 23615 6783
rect 23765 6749 23799 6783
rect 12164 6681 12198 6715
rect 14350 6681 14384 6715
rect 16681 6681 16715 6715
rect 24777 6681 24811 6715
rect 25421 6681 25455 6715
rect 13277 6613 13311 6647
rect 13737 6613 13771 6647
rect 15485 6613 15519 6647
rect 15945 6613 15979 6647
rect 16313 6613 16347 6647
rect 16773 6613 16807 6647
rect 17693 6613 17727 6647
rect 19257 6613 19291 6647
rect 21005 6613 21039 6647
rect 21465 6613 21499 6647
rect 22661 6613 22695 6647
rect 23949 6613 23983 6647
rect 24409 6613 24443 6647
rect 12265 6409 12299 6443
rect 16773 6409 16807 6443
rect 20821 6409 20855 6443
rect 25513 6409 25547 6443
rect 12449 6273 12483 6307
rect 15485 6273 15519 6307
rect 15945 6273 15979 6307
rect 16129 6273 16163 6307
rect 16221 6273 16255 6307
rect 17049 6273 17083 6307
rect 17509 6273 17543 6307
rect 17765 6273 17799 6307
rect 19809 6273 19843 6307
rect 19901 6273 19935 6307
rect 20913 6273 20947 6307
rect 22569 6273 22603 6307
rect 23213 6273 23247 6307
rect 23673 6273 23707 6307
rect 24133 6273 24167 6307
rect 24389 6273 24423 6307
rect 19993 6205 20027 6239
rect 21097 6205 21131 6239
rect 22661 6205 22695 6239
rect 22845 6205 22879 6239
rect 14749 6137 14783 6171
rect 17233 6137 17267 6171
rect 18889 6137 18923 6171
rect 23857 6137 23891 6171
rect 15669 6069 15703 6103
rect 19441 6069 19475 6103
rect 20453 6069 20487 6103
rect 22201 6069 22235 6103
rect 23397 6069 23431 6103
rect 17693 5865 17727 5899
rect 19349 5865 19383 5899
rect 21925 5865 21959 5899
rect 22201 5865 22235 5899
rect 17233 5797 17267 5831
rect 13737 5729 13771 5763
rect 18153 5729 18187 5763
rect 18337 5729 18371 5763
rect 19993 5729 20027 5763
rect 20545 5729 20579 5763
rect 23581 5729 23615 5763
rect 13470 5661 13504 5695
rect 15853 5661 15887 5695
rect 19717 5661 19751 5695
rect 23314 5661 23348 5695
rect 28089 5661 28123 5695
rect 16098 5593 16132 5627
rect 19809 5593 19843 5627
rect 20812 5593 20846 5627
rect 12357 5525 12391 5559
rect 18061 5525 18095 5559
rect 28273 5525 28307 5559
rect 17601 5321 17635 5355
rect 20821 5321 20855 5355
rect 22201 5321 22235 5355
rect 22569 5321 22603 5355
rect 22109 5253 22143 5287
rect 18981 5185 19015 5219
rect 19248 5185 19282 5219
rect 20637 5185 20671 5219
rect 22017 5117 22051 5151
rect 20361 5049 20395 5083
rect 1409 4573 1443 4607
rect 27905 4573 27939 4607
rect 28365 4573 28399 4607
rect 28181 4437 28215 4471
rect 16865 3145 16899 3179
rect 17969 3145 18003 3179
rect 1685 3009 1719 3043
rect 17325 3009 17359 3043
rect 17601 3009 17635 3043
rect 17785 3009 17819 3043
rect 1501 2805 1535 2839
rect 17233 2805 17267 2839
rect 28365 2805 28399 2839
rect 5641 2601 5675 2635
rect 15669 2601 15703 2635
rect 18153 2601 18187 2635
rect 24593 2601 24627 2635
rect 2881 2533 2915 2567
rect 8033 2533 8067 2567
rect 1685 2397 1719 2431
rect 2697 2397 2731 2431
rect 3249 2397 3283 2431
rect 6561 2397 6595 2431
rect 7849 2397 7883 2431
rect 8309 2397 8343 2431
rect 10425 2397 10459 2431
rect 15853 2397 15887 2431
rect 16129 2397 16163 2431
rect 18337 2397 18371 2431
rect 18613 2397 18647 2431
rect 20729 2397 20763 2431
rect 24777 2397 24811 2431
rect 25053 2397 25087 2431
rect 25881 2397 25915 2431
rect 27169 2397 27203 2431
rect 28365 2397 28399 2431
rect 5365 2329 5399 2363
rect 1501 2261 1535 2295
rect 4997 2261 5031 2295
rect 20913 2261 20947 2295
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 5582 27770
rect 5634 27718 5646 27770
rect 5698 27718 5710 27770
rect 5762 27718 5774 27770
rect 5826 27718 5838 27770
rect 5890 27718 14846 27770
rect 14898 27718 14910 27770
rect 14962 27718 14974 27770
rect 15026 27718 15038 27770
rect 15090 27718 15102 27770
rect 15154 27718 24110 27770
rect 24162 27718 24174 27770
rect 24226 27718 24238 27770
rect 24290 27718 24302 27770
rect 24354 27718 24366 27770
rect 24418 27718 28888 27770
rect 1104 27696 28888 27718
rect 2038 27588 2044 27600
rect 1999 27560 2044 27588
rect 2038 27548 2044 27560
rect 2096 27548 2102 27600
rect 3326 27588 3332 27600
rect 3287 27560 3332 27588
rect 3326 27548 3332 27560
rect 3384 27548 3390 27600
rect 6178 27548 6184 27600
rect 6236 27588 6242 27600
rect 6365 27591 6423 27597
rect 6365 27588 6377 27591
rect 6236 27560 6377 27588
rect 6236 27548 6242 27560
rect 6365 27557 6377 27560
rect 6411 27557 6423 27591
rect 12342 27588 12348 27600
rect 12303 27560 12348 27588
rect 6365 27551 6423 27557
rect 12342 27548 12348 27560
rect 12400 27548 12406 27600
rect 13814 27548 13820 27600
rect 13872 27588 13878 27600
rect 14277 27591 14335 27597
rect 14277 27588 14289 27591
rect 13872 27560 14289 27588
rect 13872 27548 13878 27560
rect 14277 27557 14289 27560
rect 14323 27557 14335 27591
rect 14277 27551 14335 27557
rect 14734 27548 14740 27600
rect 14792 27588 14798 27600
rect 15105 27591 15163 27597
rect 15105 27588 15117 27591
rect 14792 27560 15117 27588
rect 14792 27548 14798 27560
rect 15105 27557 15117 27560
rect 15151 27557 15163 27591
rect 15105 27551 15163 27557
rect 16114 27548 16120 27600
rect 16172 27588 16178 27600
rect 16853 27591 16911 27597
rect 16853 27588 16865 27591
rect 16172 27560 16865 27588
rect 16172 27548 16178 27560
rect 16853 27557 16865 27560
rect 16899 27557 16911 27591
rect 16853 27551 16911 27557
rect 18690 27548 18696 27600
rect 18748 27588 18754 27600
rect 19245 27591 19303 27597
rect 19245 27588 19257 27591
rect 18748 27560 19257 27588
rect 18748 27548 18754 27560
rect 19245 27557 19257 27560
rect 19291 27557 19303 27591
rect 19245 27551 19303 27557
rect 19978 27548 19984 27600
rect 20036 27588 20042 27600
rect 20349 27591 20407 27597
rect 20349 27588 20361 27591
rect 20036 27560 20361 27588
rect 20036 27548 20042 27560
rect 20349 27557 20361 27560
rect 20395 27557 20407 27591
rect 20349 27551 20407 27557
rect 21266 27548 21272 27600
rect 21324 27588 21330 27600
rect 21821 27591 21879 27597
rect 21821 27588 21833 27591
rect 21324 27560 21833 27588
rect 21324 27548 21330 27560
rect 21821 27557 21833 27560
rect 21867 27557 21879 27591
rect 21821 27551 21879 27557
rect 24949 27591 25007 27597
rect 24949 27557 24961 27591
rect 24995 27588 25007 27591
rect 25130 27588 25136 27600
rect 24995 27560 25136 27588
rect 24995 27557 25007 27560
rect 24949 27551 25007 27557
rect 25130 27548 25136 27560
rect 25188 27548 25194 27600
rect 26510 27588 26516 27600
rect 26471 27560 26516 27588
rect 26510 27548 26516 27560
rect 26568 27548 26574 27600
rect 28074 27588 28080 27600
rect 28035 27560 28080 27588
rect 28074 27548 28080 27560
rect 28132 27548 28138 27600
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27412 1458 27464
rect 3344 27452 3372 27548
rect 19797 27523 19855 27529
rect 19797 27489 19809 27523
rect 19843 27520 19855 27523
rect 21082 27520 21088 27532
rect 19843 27492 21088 27520
rect 19843 27489 19855 27492
rect 19797 27483 19855 27489
rect 21082 27480 21088 27492
rect 21140 27480 21146 27532
rect 4065 27455 4123 27461
rect 4065 27452 4077 27455
rect 3344 27424 4077 27452
rect 4065 27421 4077 27424
rect 4111 27421 4123 27455
rect 4065 27415 4123 27421
rect 13722 27412 13728 27464
rect 13780 27452 13786 27464
rect 14093 27455 14151 27461
rect 14093 27452 14105 27455
rect 13780 27424 14105 27452
rect 13780 27412 13786 27424
rect 14093 27421 14105 27424
rect 14139 27421 14151 27455
rect 14093 27415 14151 27421
rect 14642 27412 14648 27464
rect 14700 27452 14706 27464
rect 14921 27455 14979 27461
rect 14921 27452 14933 27455
rect 14700 27424 14933 27452
rect 14700 27412 14706 27424
rect 14921 27421 14933 27424
rect 14967 27421 14979 27455
rect 14921 27415 14979 27421
rect 16298 27412 16304 27464
rect 16356 27452 16362 27464
rect 16669 27455 16727 27461
rect 16669 27452 16681 27455
rect 16356 27424 16681 27452
rect 16356 27412 16362 27424
rect 16669 27421 16681 27424
rect 16715 27421 16727 27455
rect 16669 27415 16727 27421
rect 18046 27412 18052 27464
rect 18104 27452 18110 27464
rect 18141 27455 18199 27461
rect 18141 27452 18153 27455
rect 18104 27424 18153 27452
rect 18104 27412 18110 27424
rect 18141 27421 18153 27424
rect 18187 27421 18199 27455
rect 18141 27415 18199 27421
rect 19981 27455 20039 27461
rect 19981 27421 19993 27455
rect 20027 27421 20039 27455
rect 19981 27415 20039 27421
rect 20073 27455 20131 27461
rect 20073 27421 20085 27455
rect 20119 27452 20131 27455
rect 20622 27452 20628 27464
rect 20119 27424 20628 27452
rect 20119 27421 20131 27424
rect 20073 27415 20131 27421
rect 4430 27384 4436 27396
rect 4391 27356 4436 27384
rect 4430 27344 4436 27356
rect 4488 27344 4494 27396
rect 19996 27384 20024 27415
rect 20622 27412 20628 27424
rect 20680 27412 20686 27464
rect 25148 27452 25176 27548
rect 25317 27455 25375 27461
rect 25317 27452 25329 27455
rect 25148 27424 25329 27452
rect 25317 27421 25329 27424
rect 25363 27421 25375 27455
rect 26528 27452 26556 27548
rect 27249 27455 27307 27461
rect 27249 27452 27261 27455
rect 26528 27424 27261 27452
rect 25317 27415 25375 27421
rect 27249 27421 27261 27424
rect 27295 27421 27307 27455
rect 27890 27452 27896 27464
rect 27851 27424 27896 27452
rect 27249 27415 27307 27421
rect 27890 27412 27896 27424
rect 27948 27412 27954 27464
rect 20990 27384 20996 27396
rect 19996 27356 20996 27384
rect 20990 27344 20996 27356
rect 21048 27344 21054 27396
rect 25685 27387 25743 27393
rect 25685 27353 25697 27387
rect 25731 27384 25743 27387
rect 25866 27384 25872 27396
rect 25731 27356 25872 27384
rect 25731 27353 25743 27356
rect 25685 27347 25743 27353
rect 25866 27344 25872 27356
rect 25924 27344 25930 27396
rect 1578 27316 1584 27328
rect 1539 27288 1584 27316
rect 1578 27276 1584 27288
rect 1636 27276 1642 27328
rect 17954 27316 17960 27328
rect 17915 27288 17960 27316
rect 17954 27276 17960 27288
rect 18012 27276 18018 27328
rect 19797 27319 19855 27325
rect 19797 27285 19809 27319
rect 19843 27316 19855 27319
rect 20254 27316 20260 27328
rect 19843 27288 20260 27316
rect 19843 27285 19855 27288
rect 19797 27279 19855 27285
rect 20254 27276 20260 27288
rect 20312 27276 20318 27328
rect 27338 27316 27344 27328
rect 27299 27288 27344 27316
rect 27338 27276 27344 27288
rect 27396 27276 27402 27328
rect 1104 27226 28888 27248
rect 1104 27174 10214 27226
rect 10266 27174 10278 27226
rect 10330 27174 10342 27226
rect 10394 27174 10406 27226
rect 10458 27174 10470 27226
rect 10522 27174 19478 27226
rect 19530 27174 19542 27226
rect 19594 27174 19606 27226
rect 19658 27174 19670 27226
rect 19722 27174 19734 27226
rect 19786 27174 28888 27226
rect 1104 27152 28888 27174
rect 1486 27072 1492 27124
rect 1544 27112 1550 27124
rect 1857 27115 1915 27121
rect 1857 27112 1869 27115
rect 1544 27084 1869 27112
rect 1544 27072 1550 27084
rect 1857 27081 1869 27084
rect 1903 27081 1915 27115
rect 14642 27112 14648 27124
rect 14603 27084 14648 27112
rect 1857 27075 1915 27081
rect 14642 27072 14648 27084
rect 14700 27072 14706 27124
rect 16298 27112 16304 27124
rect 16259 27084 16304 27112
rect 16298 27072 16304 27084
rect 16356 27072 16362 27124
rect 20809 27115 20867 27121
rect 20809 27081 20821 27115
rect 20855 27081 20867 27115
rect 20809 27075 20867 27081
rect 21453 27115 21511 27121
rect 21453 27081 21465 27115
rect 21499 27112 21511 27115
rect 21499 27084 22094 27112
rect 21499 27081 21511 27084
rect 21453 27075 21511 27081
rect 14734 27044 14740 27056
rect 13280 27016 14740 27044
rect 1394 26976 1400 26988
rect 1355 26948 1400 26976
rect 1394 26936 1400 26948
rect 1452 26936 1458 26988
rect 13280 26985 13308 27016
rect 14734 27004 14740 27016
rect 14792 27044 14798 27056
rect 15188 27047 15246 27053
rect 14792 27016 14964 27044
rect 14792 27004 14798 27016
rect 13265 26979 13323 26985
rect 13265 26945 13277 26979
rect 13311 26945 13323 26979
rect 13265 26939 13323 26945
rect 13532 26979 13590 26985
rect 13532 26945 13544 26979
rect 13578 26976 13590 26979
rect 13998 26976 14004 26988
rect 13578 26948 14004 26976
rect 13578 26945 13590 26948
rect 13532 26939 13590 26945
rect 13998 26936 14004 26948
rect 14056 26936 14062 26988
rect 14936 26985 14964 27016
rect 15188 27013 15200 27047
rect 15234 27044 15246 27047
rect 15378 27044 15384 27056
rect 15234 27016 15384 27044
rect 15234 27013 15246 27016
rect 15188 27007 15246 27013
rect 15378 27004 15384 27016
rect 15436 27004 15442 27056
rect 17764 27047 17822 27053
rect 17764 27013 17776 27047
rect 17810 27044 17822 27047
rect 17954 27044 17960 27056
rect 17810 27016 17960 27044
rect 17810 27013 17822 27016
rect 17764 27007 17822 27013
rect 17954 27004 17960 27016
rect 18012 27004 18018 27056
rect 20288 27047 20346 27053
rect 20288 27013 20300 27047
rect 20334 27044 20346 27047
rect 20824 27044 20852 27075
rect 20334 27016 20852 27044
rect 22066 27044 22094 27084
rect 23842 27072 23848 27124
rect 23900 27112 23906 27124
rect 24029 27115 24087 27121
rect 24029 27112 24041 27115
rect 23900 27084 24041 27112
rect 23900 27072 23906 27084
rect 24029 27081 24041 27084
rect 24075 27081 24087 27115
rect 24029 27075 24087 27081
rect 26605 27115 26663 27121
rect 26605 27081 26617 27115
rect 26651 27112 26663 27115
rect 27890 27112 27896 27124
rect 26651 27084 27896 27112
rect 26651 27081 26663 27084
rect 26605 27075 26663 27081
rect 22934 27047 22992 27053
rect 22934 27044 22946 27047
rect 22066 27016 22946 27044
rect 20334 27013 20346 27016
rect 20288 27007 20346 27013
rect 22934 27013 22946 27016
rect 22980 27013 22992 27047
rect 24044 27044 24072 27075
rect 27890 27072 27896 27084
rect 27948 27072 27954 27124
rect 24489 27047 24547 27053
rect 24489 27044 24501 27047
rect 24044 27016 24501 27044
rect 22934 27007 22992 27013
rect 24489 27013 24501 27016
rect 24535 27013 24547 27047
rect 26142 27044 26148 27056
rect 24489 27007 24547 27013
rect 25240 27016 26148 27044
rect 14921 26979 14979 26985
rect 14921 26945 14933 26979
rect 14967 26945 14979 26979
rect 14921 26939 14979 26945
rect 20438 26936 20444 26988
rect 20496 26976 20502 26988
rect 20993 26979 21051 26985
rect 20993 26976 21005 26979
rect 20496 26948 21005 26976
rect 20496 26936 20502 26948
rect 20993 26945 21005 26948
rect 21039 26945 21051 26979
rect 20993 26939 21051 26945
rect 21269 26979 21327 26985
rect 21269 26945 21281 26979
rect 21315 26976 21327 26979
rect 21726 26976 21732 26988
rect 21315 26948 21732 26976
rect 21315 26945 21327 26948
rect 21269 26939 21327 26945
rect 21726 26936 21732 26948
rect 21784 26936 21790 26988
rect 17494 26908 17500 26920
rect 17455 26880 17500 26908
rect 17494 26868 17500 26880
rect 17552 26868 17558 26920
rect 20533 26911 20591 26917
rect 20533 26877 20545 26911
rect 20579 26877 20591 26911
rect 20533 26871 20591 26877
rect 23201 26911 23259 26917
rect 23201 26877 23213 26911
rect 23247 26908 23259 26911
rect 23382 26908 23388 26920
rect 23247 26880 23388 26908
rect 23247 26877 23259 26880
rect 23201 26871 23259 26877
rect 19153 26843 19211 26849
rect 19153 26809 19165 26843
rect 19199 26840 19211 26843
rect 19518 26840 19524 26852
rect 19199 26812 19524 26840
rect 19199 26809 19211 26812
rect 19153 26803 19211 26809
rect 19518 26800 19524 26812
rect 19576 26800 19582 26852
rect 18877 26775 18935 26781
rect 18877 26741 18889 26775
rect 18923 26772 18935 26775
rect 19058 26772 19064 26784
rect 18923 26744 19064 26772
rect 18923 26741 18935 26744
rect 18877 26735 18935 26741
rect 19058 26732 19064 26744
rect 19116 26732 19122 26784
rect 19334 26732 19340 26784
rect 19392 26772 19398 26784
rect 20548 26772 20576 26871
rect 23382 26868 23388 26880
rect 23440 26908 23446 26920
rect 25240 26917 25268 27016
rect 26142 27004 26148 27016
rect 26200 27044 26206 27056
rect 26200 27016 27016 27044
rect 26200 27004 26206 27016
rect 25498 26985 25504 26988
rect 25492 26976 25504 26985
rect 25459 26948 25504 26976
rect 25492 26939 25504 26948
rect 25498 26936 25504 26939
rect 25556 26936 25562 26988
rect 26988 26985 27016 27016
rect 26973 26979 27031 26985
rect 26973 26945 26985 26979
rect 27019 26945 27031 26979
rect 27229 26979 27287 26985
rect 27229 26976 27241 26979
rect 26973 26939 27031 26945
rect 27080 26948 27241 26976
rect 25225 26911 25283 26917
rect 25225 26908 25237 26911
rect 23440 26880 25237 26908
rect 23440 26868 23446 26880
rect 25225 26877 25237 26880
rect 25271 26877 25283 26911
rect 25225 26871 25283 26877
rect 26694 26868 26700 26920
rect 26752 26908 26758 26920
rect 27080 26908 27108 26948
rect 27229 26945 27241 26948
rect 27275 26945 27287 26979
rect 27229 26939 27287 26945
rect 26752 26880 27108 26908
rect 26752 26868 26758 26880
rect 24670 26840 24676 26852
rect 24631 26812 24676 26840
rect 24670 26800 24676 26812
rect 24728 26800 24734 26852
rect 19392 26744 20576 26772
rect 21821 26775 21879 26781
rect 19392 26732 19398 26744
rect 21821 26741 21833 26775
rect 21867 26772 21879 26775
rect 22186 26772 22192 26784
rect 21867 26744 22192 26772
rect 21867 26741 21879 26744
rect 21821 26735 21879 26741
rect 22186 26732 22192 26744
rect 22244 26732 22250 26784
rect 28350 26772 28356 26784
rect 28311 26744 28356 26772
rect 28350 26732 28356 26744
rect 28408 26732 28414 26784
rect 1104 26682 28888 26704
rect 1104 26630 5582 26682
rect 5634 26630 5646 26682
rect 5698 26630 5710 26682
rect 5762 26630 5774 26682
rect 5826 26630 5838 26682
rect 5890 26630 14846 26682
rect 14898 26630 14910 26682
rect 14962 26630 14974 26682
rect 15026 26630 15038 26682
rect 15090 26630 15102 26682
rect 15154 26630 24110 26682
rect 24162 26630 24174 26682
rect 24226 26630 24238 26682
rect 24290 26630 24302 26682
rect 24354 26630 24366 26682
rect 24418 26630 28888 26682
rect 1104 26608 28888 26630
rect 18046 26568 18052 26580
rect 18007 26540 18052 26568
rect 18046 26528 18052 26540
rect 18104 26528 18110 26580
rect 18230 26568 18236 26580
rect 18191 26540 18236 26568
rect 18230 26528 18236 26540
rect 18288 26528 18294 26580
rect 19337 26571 19395 26577
rect 19337 26537 19349 26571
rect 19383 26568 19395 26571
rect 20257 26571 20315 26577
rect 20257 26568 20269 26571
rect 19383 26540 20269 26568
rect 19383 26537 19395 26540
rect 19337 26531 19395 26537
rect 20257 26537 20269 26540
rect 20303 26537 20315 26571
rect 20438 26568 20444 26580
rect 20399 26540 20444 26568
rect 20257 26531 20315 26537
rect 20438 26528 20444 26540
rect 20496 26528 20502 26580
rect 21453 26571 21511 26577
rect 21453 26537 21465 26571
rect 21499 26568 21511 26571
rect 21913 26571 21971 26577
rect 21913 26568 21925 26571
rect 21499 26540 21925 26568
rect 21499 26537 21511 26540
rect 21453 26531 21511 26537
rect 21913 26537 21925 26540
rect 21959 26537 21971 26571
rect 21913 26531 21971 26537
rect 27522 26528 27528 26580
rect 27580 26568 27586 26580
rect 28169 26571 28227 26577
rect 28169 26568 28181 26571
rect 27580 26540 28181 26568
rect 27580 26528 27586 26540
rect 28169 26537 28181 26540
rect 28215 26537 28227 26571
rect 28169 26531 28227 26537
rect 21726 26500 21732 26512
rect 21687 26472 21732 26500
rect 21726 26460 21732 26472
rect 21784 26460 21790 26512
rect 19444 26404 20116 26432
rect 1670 26364 1676 26376
rect 1583 26336 1676 26364
rect 1670 26324 1676 26336
rect 1728 26364 1734 26376
rect 2133 26367 2191 26373
rect 2133 26364 2145 26367
rect 1728 26336 2145 26364
rect 1728 26324 1734 26336
rect 2133 26333 2145 26336
rect 2179 26333 2191 26367
rect 2133 26327 2191 26333
rect 16117 26367 16175 26373
rect 16117 26333 16129 26367
rect 16163 26364 16175 26367
rect 17494 26364 17500 26376
rect 16163 26336 17500 26364
rect 16163 26333 16175 26336
rect 16117 26327 16175 26333
rect 17494 26324 17500 26336
rect 17552 26364 17558 26376
rect 19334 26364 19340 26376
rect 17552 26336 19340 26364
rect 17552 26324 17558 26336
rect 19334 26324 19340 26336
rect 19392 26324 19398 26376
rect 1762 26256 1768 26308
rect 1820 26296 1826 26308
rect 1857 26299 1915 26305
rect 1857 26296 1869 26299
rect 1820 26268 1869 26296
rect 1820 26256 1826 26268
rect 1857 26265 1869 26268
rect 1903 26265 1915 26299
rect 1857 26259 1915 26265
rect 16384 26299 16442 26305
rect 16384 26265 16396 26299
rect 16430 26296 16442 26299
rect 16666 26296 16672 26308
rect 16430 26268 16672 26296
rect 16430 26265 16442 26268
rect 16384 26259 16442 26265
rect 16666 26256 16672 26268
rect 16724 26256 16730 26308
rect 18217 26299 18275 26305
rect 18217 26265 18229 26299
rect 18263 26296 18275 26299
rect 18322 26296 18328 26308
rect 18263 26268 18328 26296
rect 18263 26265 18275 26268
rect 18217 26259 18275 26265
rect 18322 26256 18328 26268
rect 18380 26256 18386 26308
rect 18414 26256 18420 26308
rect 18472 26296 18478 26308
rect 19444 26296 19472 26404
rect 19518 26324 19524 26376
rect 19576 26364 19582 26376
rect 19797 26367 19855 26373
rect 19576 26336 19669 26364
rect 19576 26324 19582 26336
rect 19797 26333 19809 26367
rect 19843 26364 19855 26367
rect 19978 26364 19984 26376
rect 19843 26336 19984 26364
rect 19843 26333 19855 26336
rect 19797 26327 19855 26333
rect 19978 26324 19984 26336
rect 20036 26324 20042 26376
rect 20088 26364 20116 26404
rect 20990 26364 20996 26376
rect 20088 26336 20392 26364
rect 20951 26336 20996 26364
rect 18472 26268 19472 26296
rect 19536 26296 19564 26324
rect 19886 26296 19892 26308
rect 19536 26268 19892 26296
rect 18472 26256 18478 26268
rect 19886 26256 19892 26268
rect 19944 26256 19950 26308
rect 20088 26305 20116 26336
rect 20073 26299 20131 26305
rect 20073 26265 20085 26299
rect 20119 26265 20131 26299
rect 20073 26259 20131 26265
rect 20254 26256 20260 26308
rect 20312 26305 20318 26308
rect 20312 26299 20331 26305
rect 20319 26265 20331 26299
rect 20364 26296 20392 26336
rect 20990 26324 20996 26336
rect 21048 26324 21054 26376
rect 21269 26367 21327 26373
rect 21269 26333 21281 26367
rect 21315 26364 21327 26367
rect 22186 26364 22192 26376
rect 21315 26336 22192 26364
rect 21315 26333 21327 26336
rect 21269 26327 21327 26333
rect 22186 26324 22192 26336
rect 22244 26324 22250 26376
rect 28350 26364 28356 26376
rect 28311 26336 28356 26364
rect 28350 26324 28356 26336
rect 28408 26324 28414 26376
rect 22097 26299 22155 26305
rect 22097 26296 22109 26299
rect 20364 26268 22109 26296
rect 20312 26259 20331 26265
rect 22097 26265 22109 26268
rect 22143 26265 22155 26299
rect 25130 26296 25136 26308
rect 25091 26268 25136 26296
rect 22097 26259 22155 26265
rect 20312 26256 20318 26259
rect 25130 26256 25136 26268
rect 25188 26256 25194 26308
rect 26694 26256 26700 26308
rect 26752 26296 26758 26308
rect 26789 26299 26847 26305
rect 26789 26296 26801 26299
rect 26752 26268 26801 26296
rect 26752 26256 26758 26268
rect 26789 26265 26801 26268
rect 26835 26265 26847 26299
rect 26789 26259 26847 26265
rect 17497 26231 17555 26237
rect 17497 26197 17509 26231
rect 17543 26228 17555 26231
rect 17586 26228 17592 26240
rect 17543 26200 17592 26228
rect 17543 26197 17555 26200
rect 17497 26191 17555 26197
rect 17586 26188 17592 26200
rect 17644 26188 17650 26240
rect 19705 26231 19763 26237
rect 19705 26197 19717 26231
rect 19751 26228 19763 26231
rect 21082 26228 21088 26240
rect 19751 26200 21088 26228
rect 19751 26197 19763 26200
rect 19705 26191 19763 26197
rect 21082 26188 21088 26200
rect 21140 26188 21146 26240
rect 21910 26237 21916 26240
rect 21897 26231 21916 26237
rect 21897 26197 21909 26231
rect 21897 26191 21916 26197
rect 21910 26188 21916 26191
rect 21968 26188 21974 26240
rect 1104 26138 28888 26160
rect 1104 26086 10214 26138
rect 10266 26086 10278 26138
rect 10330 26086 10342 26138
rect 10394 26086 10406 26138
rect 10458 26086 10470 26138
rect 10522 26086 19478 26138
rect 19530 26086 19542 26138
rect 19594 26086 19606 26138
rect 19658 26086 19670 26138
rect 19722 26086 19734 26138
rect 19786 26086 28888 26138
rect 1104 26064 28888 26086
rect 16666 26024 16672 26036
rect 16627 25996 16672 26024
rect 16666 25984 16672 25996
rect 16724 25984 16730 26036
rect 17310 26024 17316 26036
rect 16868 25996 17316 26024
rect 16301 25959 16359 25965
rect 16301 25925 16313 25959
rect 16347 25956 16359 25959
rect 16868 25956 16896 25996
rect 17310 25984 17316 25996
rect 17368 25984 17374 26036
rect 18230 25984 18236 26036
rect 18288 26024 18294 26036
rect 18325 26027 18383 26033
rect 18325 26024 18337 26027
rect 18288 25996 18337 26024
rect 18288 25984 18294 25996
rect 18325 25993 18337 25996
rect 18371 25993 18383 26027
rect 18325 25987 18383 25993
rect 18506 25984 18512 26036
rect 18564 26024 18570 26036
rect 20254 26024 20260 26036
rect 18564 25996 20260 26024
rect 18564 25984 18570 25996
rect 20254 25984 20260 25996
rect 20312 25984 20318 26036
rect 21450 25984 21456 26036
rect 21508 26024 21514 26036
rect 21910 26024 21916 26036
rect 21508 25996 21916 26024
rect 21508 25984 21514 25996
rect 21910 25984 21916 25996
rect 21968 26024 21974 26036
rect 22557 26027 22615 26033
rect 22557 26024 22569 26027
rect 21968 25996 22569 26024
rect 21968 25984 21974 25996
rect 22557 25993 22569 25996
rect 22603 25993 22615 26027
rect 22557 25987 22615 25993
rect 16347 25928 16896 25956
rect 16960 25928 17724 25956
rect 16347 25925 16359 25928
rect 16301 25919 16359 25925
rect 15470 25888 15476 25900
rect 15431 25860 15476 25888
rect 15470 25848 15476 25860
rect 15528 25848 15534 25900
rect 16960 25897 16988 25928
rect 17696 25900 17724 25928
rect 16945 25891 17003 25897
rect 16945 25857 16957 25891
rect 16991 25857 17003 25891
rect 16945 25851 17003 25857
rect 17037 25891 17095 25897
rect 17037 25857 17049 25891
rect 17083 25857 17095 25891
rect 17037 25851 17095 25857
rect 17052 25752 17080 25851
rect 17126 25848 17132 25900
rect 17184 25888 17190 25900
rect 17184 25860 17229 25888
rect 17184 25848 17190 25860
rect 17310 25848 17316 25900
rect 17368 25888 17374 25900
rect 17368 25860 17413 25888
rect 17368 25848 17374 25860
rect 17494 25848 17500 25900
rect 17552 25888 17558 25900
rect 17589 25891 17647 25897
rect 17589 25888 17601 25891
rect 17552 25860 17601 25888
rect 17552 25848 17558 25860
rect 17589 25857 17601 25860
rect 17635 25857 17647 25891
rect 17589 25851 17647 25857
rect 17678 25848 17684 25900
rect 17736 25888 17742 25900
rect 17773 25891 17831 25897
rect 17773 25888 17785 25891
rect 17736 25860 17785 25888
rect 17736 25848 17742 25860
rect 17773 25857 17785 25860
rect 17819 25857 17831 25891
rect 18524 25888 18552 25984
rect 19150 25916 19156 25968
rect 19208 25956 19214 25968
rect 19245 25959 19303 25965
rect 19245 25956 19257 25959
rect 19208 25928 19257 25956
rect 19208 25916 19214 25928
rect 19245 25925 19257 25928
rect 19291 25925 19303 25959
rect 19445 25959 19503 25965
rect 19445 25956 19457 25959
rect 19245 25919 19303 25925
rect 19352 25928 19457 25956
rect 18590 25891 18648 25897
rect 18590 25888 18602 25891
rect 18524 25860 18602 25888
rect 17773 25851 17831 25857
rect 18590 25857 18602 25860
rect 18636 25857 18648 25891
rect 18590 25851 18648 25857
rect 18690 25848 18696 25900
rect 18748 25888 18754 25900
rect 18748 25860 18793 25888
rect 18748 25848 18754 25860
rect 19058 25848 19064 25900
rect 19116 25888 19122 25900
rect 19352 25888 19380 25928
rect 19445 25925 19457 25928
rect 19491 25925 19503 25959
rect 19445 25919 19503 25925
rect 20714 25916 20720 25968
rect 20772 25956 20778 25968
rect 22186 25956 22192 25968
rect 20772 25928 22192 25956
rect 20772 25916 20778 25928
rect 19116 25860 19380 25888
rect 20073 25891 20131 25897
rect 19116 25848 19122 25860
rect 20073 25857 20085 25891
rect 20119 25888 20131 25891
rect 20119 25860 20760 25888
rect 20119 25857 20131 25860
rect 20073 25851 20131 25857
rect 18322 25780 18328 25832
rect 18380 25820 18386 25832
rect 18509 25823 18567 25829
rect 18509 25820 18521 25823
rect 18380 25792 18521 25820
rect 18380 25780 18386 25792
rect 18509 25789 18521 25792
rect 18555 25789 18567 25823
rect 18509 25783 18567 25789
rect 18785 25823 18843 25829
rect 18785 25789 18797 25823
rect 18831 25820 18843 25823
rect 19150 25820 19156 25832
rect 18831 25792 19156 25820
rect 18831 25789 18843 25792
rect 18785 25783 18843 25789
rect 19150 25780 19156 25792
rect 19208 25780 19214 25832
rect 19889 25823 19947 25829
rect 19889 25820 19901 25823
rect 19260 25792 19901 25820
rect 17052 25724 17724 25752
rect 15286 25684 15292 25696
rect 15247 25656 15292 25684
rect 15286 25644 15292 25656
rect 15344 25644 15350 25696
rect 17218 25644 17224 25696
rect 17276 25684 17282 25696
rect 17589 25687 17647 25693
rect 17589 25684 17601 25687
rect 17276 25656 17601 25684
rect 17276 25644 17282 25656
rect 17589 25653 17601 25656
rect 17635 25653 17647 25687
rect 17696 25684 17724 25724
rect 18690 25712 18696 25764
rect 18748 25712 18754 25764
rect 18966 25712 18972 25764
rect 19024 25752 19030 25764
rect 19260 25752 19288 25792
rect 19889 25789 19901 25792
rect 19935 25789 19947 25823
rect 19889 25783 19947 25789
rect 19978 25780 19984 25832
rect 20036 25780 20042 25832
rect 20254 25780 20260 25832
rect 20312 25820 20318 25832
rect 20732 25829 20760 25860
rect 20990 25848 20996 25900
rect 21048 25888 21054 25900
rect 21928 25897 21956 25928
rect 22186 25916 22192 25928
rect 22244 25916 22250 25968
rect 22281 25959 22339 25965
rect 22281 25925 22293 25959
rect 22327 25956 22339 25959
rect 25682 25956 25688 25968
rect 22327 25928 22784 25956
rect 25643 25928 25688 25956
rect 22327 25925 22339 25928
rect 22281 25919 22339 25925
rect 21821 25891 21879 25897
rect 21821 25888 21833 25891
rect 21048 25860 21833 25888
rect 21048 25848 21054 25860
rect 21821 25857 21833 25860
rect 21867 25857 21879 25891
rect 21821 25851 21879 25857
rect 21913 25891 21971 25897
rect 21913 25857 21925 25891
rect 21959 25857 21971 25891
rect 22094 25888 22100 25900
rect 22055 25860 22100 25888
rect 21913 25851 21971 25857
rect 22094 25848 22100 25860
rect 22152 25848 22158 25900
rect 22756 25897 22784 25928
rect 25682 25916 25688 25928
rect 25740 25916 25746 25968
rect 23750 25897 23756 25900
rect 22557 25891 22615 25897
rect 22557 25857 22569 25891
rect 22603 25857 22615 25891
rect 22557 25851 22615 25857
rect 22741 25891 22799 25897
rect 22741 25857 22753 25891
rect 22787 25857 22799 25891
rect 22741 25851 22799 25857
rect 23744 25851 23756 25897
rect 23808 25888 23814 25900
rect 25406 25888 25412 25900
rect 23808 25860 23844 25888
rect 25367 25860 25412 25888
rect 20441 25823 20499 25829
rect 20441 25820 20453 25823
rect 20312 25792 20453 25820
rect 20312 25780 20318 25792
rect 20441 25789 20453 25792
rect 20487 25789 20499 25823
rect 20441 25783 20499 25789
rect 20717 25823 20775 25829
rect 20717 25789 20729 25823
rect 20763 25820 20775 25823
rect 21082 25820 21088 25832
rect 20763 25792 21088 25820
rect 20763 25789 20775 25792
rect 20717 25783 20775 25789
rect 21082 25780 21088 25792
rect 21140 25820 21146 25832
rect 22572 25820 22600 25851
rect 23750 25848 23756 25851
rect 23808 25848 23814 25860
rect 25406 25848 25412 25860
rect 25464 25848 25470 25900
rect 25590 25888 25596 25900
rect 25551 25860 25596 25888
rect 25590 25848 25596 25860
rect 25648 25848 25654 25900
rect 25774 25888 25780 25900
rect 25735 25860 25780 25888
rect 25774 25848 25780 25860
rect 25832 25848 25838 25900
rect 21140 25792 22600 25820
rect 21140 25780 21146 25792
rect 23382 25780 23388 25832
rect 23440 25820 23446 25832
rect 23477 25823 23535 25829
rect 23477 25820 23489 25823
rect 23440 25792 23489 25820
rect 23440 25780 23446 25792
rect 23477 25789 23489 25792
rect 23523 25789 23535 25823
rect 23477 25783 23535 25789
rect 19024 25724 19288 25752
rect 19613 25755 19671 25761
rect 19024 25712 19030 25724
rect 19613 25721 19625 25755
rect 19659 25752 19671 25755
rect 19996 25752 20024 25780
rect 20530 25752 20536 25764
rect 19659 25724 20536 25752
rect 19659 25721 19671 25724
rect 19613 25715 19671 25721
rect 20530 25712 20536 25724
rect 20588 25712 20594 25764
rect 20622 25712 20628 25764
rect 20680 25752 20686 25764
rect 22094 25752 22100 25764
rect 20680 25724 22100 25752
rect 20680 25712 20686 25724
rect 22094 25712 22100 25724
rect 22152 25712 22158 25764
rect 18598 25684 18604 25696
rect 17696 25656 18604 25684
rect 17589 25647 17647 25653
rect 18598 25644 18604 25656
rect 18656 25644 18662 25696
rect 18708 25684 18736 25712
rect 19429 25687 19487 25693
rect 19429 25684 19441 25687
rect 18708 25656 19441 25684
rect 19429 25653 19441 25656
rect 19475 25684 19487 25687
rect 19518 25684 19524 25696
rect 19475 25656 19524 25684
rect 19475 25653 19487 25656
rect 19429 25647 19487 25653
rect 19518 25644 19524 25656
rect 19576 25644 19582 25696
rect 24762 25644 24768 25696
rect 24820 25684 24826 25696
rect 24857 25687 24915 25693
rect 24857 25684 24869 25687
rect 24820 25656 24869 25684
rect 24820 25644 24826 25656
rect 24857 25653 24869 25656
rect 24903 25653 24915 25687
rect 25958 25684 25964 25696
rect 25919 25656 25964 25684
rect 24857 25647 24915 25653
rect 25958 25644 25964 25656
rect 26016 25644 26022 25696
rect 1104 25594 28888 25616
rect 1104 25542 5582 25594
rect 5634 25542 5646 25594
rect 5698 25542 5710 25594
rect 5762 25542 5774 25594
rect 5826 25542 5838 25594
rect 5890 25542 14846 25594
rect 14898 25542 14910 25594
rect 14962 25542 14974 25594
rect 15026 25542 15038 25594
rect 15090 25542 15102 25594
rect 15154 25542 24110 25594
rect 24162 25542 24174 25594
rect 24226 25542 24238 25594
rect 24290 25542 24302 25594
rect 24354 25542 24366 25594
rect 24418 25542 28888 25594
rect 1104 25520 28888 25542
rect 17126 25480 17132 25492
rect 17087 25452 17132 25480
rect 17126 25440 17132 25452
rect 17184 25440 17190 25492
rect 17218 25440 17224 25492
rect 17276 25480 17282 25492
rect 17276 25452 17321 25480
rect 17276 25440 17282 25452
rect 23750 25440 23756 25492
rect 23808 25480 23814 25492
rect 23845 25483 23903 25489
rect 23845 25480 23857 25483
rect 23808 25452 23857 25480
rect 23808 25440 23814 25452
rect 23845 25449 23857 25452
rect 23891 25449 23903 25483
rect 23845 25443 23903 25449
rect 25682 25440 25688 25492
rect 25740 25480 25746 25492
rect 25777 25483 25835 25489
rect 25777 25480 25789 25483
rect 25740 25452 25789 25480
rect 25740 25440 25746 25452
rect 25777 25449 25789 25452
rect 25823 25449 25835 25483
rect 25777 25443 25835 25449
rect 16574 25412 16580 25424
rect 16535 25384 16580 25412
rect 16574 25372 16580 25384
rect 16632 25372 16638 25424
rect 16850 25372 16856 25424
rect 16908 25412 16914 25424
rect 16908 25384 17807 25412
rect 16908 25372 16914 25384
rect 14734 25304 14740 25356
rect 14792 25344 14798 25356
rect 17779 25353 17807 25384
rect 18322 25372 18328 25424
rect 18380 25412 18386 25424
rect 19058 25412 19064 25424
rect 18380 25384 19064 25412
rect 18380 25372 18386 25384
rect 19058 25372 19064 25384
rect 19116 25412 19122 25424
rect 22002 25412 22008 25424
rect 19116 25384 19656 25412
rect 19116 25372 19122 25384
rect 14829 25347 14887 25353
rect 14829 25344 14841 25347
rect 14792 25316 14841 25344
rect 14792 25304 14798 25316
rect 14829 25313 14841 25316
rect 14875 25313 14887 25347
rect 14829 25307 14887 25313
rect 16485 25347 16543 25353
rect 16485 25313 16497 25347
rect 16531 25313 16543 25347
rect 17773 25347 17831 25353
rect 16485 25307 16543 25313
rect 16776 25316 17540 25344
rect 15096 25211 15154 25217
rect 15096 25177 15108 25211
rect 15142 25208 15154 25211
rect 15286 25208 15292 25220
rect 15142 25180 15292 25208
rect 15142 25177 15154 25180
rect 15096 25171 15154 25177
rect 15286 25168 15292 25180
rect 15344 25168 15350 25220
rect 16500 25208 16528 25307
rect 16666 25276 16672 25288
rect 16627 25248 16672 25276
rect 16666 25236 16672 25248
rect 16724 25236 16730 25288
rect 16776 25285 16804 25316
rect 17402 25285 17408 25288
rect 16761 25279 16819 25285
rect 16761 25245 16773 25279
rect 16807 25245 16819 25279
rect 17037 25279 17095 25285
rect 17037 25276 17049 25279
rect 16761 25239 16819 25245
rect 16960 25248 17049 25276
rect 16960 25208 16988 25248
rect 17037 25245 17049 25248
rect 17083 25276 17095 25279
rect 17359 25279 17408 25285
rect 17083 25248 17264 25276
rect 17083 25245 17095 25248
rect 17037 25239 17095 25245
rect 16500 25180 16988 25208
rect 17236 25208 17264 25248
rect 17359 25245 17371 25279
rect 17405 25245 17408 25279
rect 17359 25239 17408 25245
rect 17402 25236 17408 25239
rect 17460 25236 17466 25288
rect 17512 25285 17540 25316
rect 17773 25313 17785 25347
rect 17819 25344 17831 25347
rect 18506 25344 18512 25356
rect 17819 25316 18512 25344
rect 17819 25313 17831 25316
rect 17773 25307 17831 25313
rect 18506 25304 18512 25316
rect 18564 25304 18570 25356
rect 19628 25344 19656 25384
rect 20364 25384 22008 25412
rect 20364 25353 20392 25384
rect 22002 25372 22008 25384
rect 22060 25372 22066 25424
rect 20349 25347 20407 25353
rect 19628 25316 19748 25344
rect 17497 25279 17555 25285
rect 17497 25245 17509 25279
rect 17543 25276 17555 25279
rect 18064 25276 18184 25286
rect 19429 25279 19487 25285
rect 19429 25276 19441 25279
rect 17543 25273 17724 25276
rect 17880 25273 19441 25276
rect 17543 25258 19441 25273
rect 17543 25248 18092 25258
rect 18156 25248 19441 25258
rect 17543 25245 17555 25248
rect 17696 25245 17908 25248
rect 19429 25245 19441 25248
rect 19475 25245 19487 25279
rect 17497 25239 17555 25245
rect 19429 25239 19487 25245
rect 19444 25208 19472 25239
rect 19518 25236 19524 25288
rect 19576 25276 19582 25288
rect 19720 25285 19748 25316
rect 20349 25313 20361 25347
rect 20395 25313 20407 25347
rect 20349 25307 20407 25313
rect 20441 25347 20499 25353
rect 20441 25313 20453 25347
rect 20487 25344 20499 25347
rect 20714 25344 20720 25356
rect 20487 25316 20720 25344
rect 20487 25313 20499 25316
rect 20441 25307 20499 25313
rect 20714 25304 20720 25316
rect 20772 25304 20778 25356
rect 20809 25347 20867 25353
rect 20809 25313 20821 25347
rect 20855 25344 20867 25347
rect 22370 25344 22376 25356
rect 20855 25316 21312 25344
rect 20855 25313 20867 25316
rect 20809 25307 20867 25313
rect 19705 25279 19763 25285
rect 19576 25248 19656 25276
rect 19576 25236 19582 25248
rect 19628 25217 19656 25248
rect 19705 25245 19717 25279
rect 19751 25245 19763 25279
rect 20533 25279 20591 25285
rect 20533 25276 20545 25279
rect 19705 25239 19763 25245
rect 20364 25248 20545 25276
rect 20364 25220 20392 25248
rect 20533 25245 20545 25248
rect 20579 25245 20591 25279
rect 20533 25239 20591 25245
rect 20625 25279 20683 25285
rect 20625 25245 20637 25279
rect 20671 25276 20683 25279
rect 20898 25276 20904 25288
rect 20671 25248 20904 25276
rect 20671 25245 20683 25248
rect 20625 25239 20683 25245
rect 20898 25236 20904 25248
rect 20956 25236 20962 25288
rect 21082 25276 21088 25288
rect 21043 25248 21088 25276
rect 21082 25236 21088 25248
rect 21140 25236 21146 25288
rect 21284 25285 21312 25316
rect 21376 25316 22376 25344
rect 21376 25285 21404 25316
rect 22370 25304 22376 25316
rect 22428 25304 22434 25356
rect 24762 25304 24768 25356
rect 24820 25344 24826 25356
rect 24949 25347 25007 25353
rect 24949 25344 24961 25347
rect 24820 25316 24961 25344
rect 24820 25304 24826 25316
rect 24949 25313 24961 25316
rect 24995 25313 25007 25347
rect 24949 25307 25007 25313
rect 25774 25304 25780 25356
rect 25832 25304 25838 25356
rect 21269 25279 21327 25285
rect 21269 25245 21281 25279
rect 21315 25245 21327 25279
rect 21269 25239 21327 25245
rect 21361 25279 21419 25285
rect 21361 25245 21373 25279
rect 21407 25245 21419 25279
rect 21361 25239 21419 25245
rect 21450 25236 21456 25288
rect 21508 25276 21514 25288
rect 21508 25248 21553 25276
rect 21508 25236 21514 25248
rect 22646 25236 22652 25288
rect 22704 25276 22710 25288
rect 23382 25276 23388 25288
rect 22704 25248 23388 25276
rect 22704 25236 22710 25248
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 24029 25279 24087 25285
rect 24029 25245 24041 25279
rect 24075 25276 24087 25279
rect 24854 25276 24860 25288
rect 24075 25248 24440 25276
rect 24767 25248 24860 25276
rect 24075 25245 24087 25248
rect 24029 25239 24087 25245
rect 19613 25211 19671 25217
rect 17236 25180 18046 25208
rect 19444 25180 19533 25208
rect 16206 25140 16212 25152
rect 16167 25112 16212 25140
rect 16206 25100 16212 25112
rect 16264 25100 16270 25152
rect 16666 25100 16672 25152
rect 16724 25140 16730 25152
rect 17494 25140 17500 25152
rect 16724 25112 17500 25140
rect 16724 25100 16730 25112
rect 17494 25100 17500 25112
rect 17552 25100 17558 25152
rect 18018 25149 18046 25180
rect 18003 25143 18061 25149
rect 18003 25109 18015 25143
rect 18049 25140 18061 25143
rect 19058 25140 19064 25152
rect 18049 25112 19064 25140
rect 18049 25109 18061 25112
rect 18003 25103 18061 25109
rect 19058 25100 19064 25112
rect 19116 25100 19122 25152
rect 19242 25140 19248 25152
rect 19203 25112 19248 25140
rect 19242 25100 19248 25112
rect 19300 25100 19306 25152
rect 19505 25140 19533 25180
rect 19613 25177 19625 25211
rect 19659 25208 19671 25211
rect 20162 25208 20168 25220
rect 19659 25180 20168 25208
rect 19659 25177 19671 25180
rect 19613 25171 19671 25177
rect 20162 25168 20168 25180
rect 20220 25168 20226 25220
rect 20346 25168 20352 25220
rect 20404 25168 20410 25220
rect 21729 25211 21787 25217
rect 21729 25177 21741 25211
rect 21775 25208 21787 25211
rect 23118 25211 23176 25217
rect 23118 25208 23130 25211
rect 21775 25180 23130 25208
rect 21775 25177 21787 25180
rect 21729 25171 21787 25177
rect 23118 25177 23130 25180
rect 23164 25177 23176 25211
rect 23118 25171 23176 25177
rect 21266 25140 21272 25152
rect 19505 25112 21272 25140
rect 21266 25100 21272 25112
rect 21324 25100 21330 25152
rect 24412 25149 24440 25248
rect 24854 25236 24860 25248
rect 24912 25276 24918 25288
rect 25792 25276 25820 25304
rect 24912 25248 25820 25276
rect 24912 25236 24918 25248
rect 26142 25236 26148 25288
rect 26200 25276 26206 25288
rect 27157 25279 27215 25285
rect 27157 25276 27169 25279
rect 26200 25248 27169 25276
rect 26200 25236 26206 25248
rect 27157 25245 27169 25248
rect 27203 25245 27215 25279
rect 27157 25239 27215 25245
rect 24765 25211 24823 25217
rect 24765 25177 24777 25211
rect 24811 25208 24823 25211
rect 25406 25208 25412 25220
rect 24811 25180 25412 25208
rect 24811 25177 24823 25180
rect 24765 25171 24823 25177
rect 25406 25168 25412 25180
rect 25464 25208 25470 25220
rect 25774 25208 25780 25220
rect 25464 25180 25780 25208
rect 25464 25168 25470 25180
rect 25774 25168 25780 25180
rect 25832 25168 25838 25220
rect 25958 25168 25964 25220
rect 26016 25208 26022 25220
rect 26890 25211 26948 25217
rect 26890 25208 26902 25211
rect 26016 25180 26902 25208
rect 26016 25168 26022 25180
rect 26890 25177 26902 25180
rect 26936 25177 26948 25211
rect 26890 25171 26948 25177
rect 24397 25143 24455 25149
rect 24397 25109 24409 25143
rect 24443 25109 24455 25143
rect 24397 25103 24455 25109
rect 1104 25050 28888 25072
rect 1104 24998 10214 25050
rect 10266 24998 10278 25050
rect 10330 24998 10342 25050
rect 10394 24998 10406 25050
rect 10458 24998 10470 25050
rect 10522 24998 19478 25050
rect 19530 24998 19542 25050
rect 19594 24998 19606 25050
rect 19658 24998 19670 25050
rect 19722 24998 19734 25050
rect 19786 24998 28888 25050
rect 1104 24976 28888 24998
rect 15470 24896 15476 24948
rect 15528 24936 15534 24948
rect 15841 24939 15899 24945
rect 15841 24936 15853 24939
rect 15528 24908 15853 24936
rect 15528 24896 15534 24908
rect 15841 24905 15853 24908
rect 15887 24905 15899 24939
rect 19058 24936 19064 24948
rect 19019 24908 19064 24936
rect 15841 24899 15899 24905
rect 19058 24896 19064 24908
rect 19116 24896 19122 24948
rect 19150 24896 19156 24948
rect 19208 24936 19214 24948
rect 19705 24939 19763 24945
rect 19705 24936 19717 24939
rect 19208 24908 19717 24936
rect 19208 24896 19214 24908
rect 19705 24905 19717 24908
rect 19751 24936 19763 24939
rect 19978 24936 19984 24948
rect 19751 24908 19984 24936
rect 19751 24905 19763 24908
rect 19705 24899 19763 24905
rect 19978 24896 19984 24908
rect 20036 24896 20042 24948
rect 20073 24939 20131 24945
rect 20073 24905 20085 24939
rect 20119 24936 20131 24939
rect 20898 24936 20904 24948
rect 20119 24908 20904 24936
rect 20119 24905 20131 24908
rect 20073 24899 20131 24905
rect 20898 24896 20904 24908
rect 20956 24896 20962 24948
rect 21266 24936 21272 24948
rect 21179 24908 21272 24936
rect 21266 24896 21272 24908
rect 21324 24936 21330 24948
rect 21324 24908 22223 24936
rect 21324 24896 21330 24908
rect 16009 24871 16067 24877
rect 16009 24837 16021 24871
rect 16055 24868 16067 24871
rect 16209 24871 16267 24877
rect 16055 24837 16068 24868
rect 16009 24831 16068 24837
rect 16209 24837 16221 24871
rect 16255 24868 16267 24871
rect 16298 24868 16304 24880
rect 16255 24840 16304 24868
rect 16255 24837 16267 24840
rect 16209 24831 16267 24837
rect 15013 24803 15071 24809
rect 15013 24769 15025 24803
rect 15059 24800 15071 24803
rect 15470 24800 15476 24812
rect 15059 24772 15476 24800
rect 15059 24769 15071 24772
rect 15013 24763 15071 24769
rect 15470 24760 15476 24772
rect 15528 24760 15534 24812
rect 16040 24800 16068 24831
rect 16298 24828 16304 24840
rect 16356 24868 16362 24880
rect 18414 24868 18420 24880
rect 16356 24840 18420 24868
rect 16356 24828 16362 24840
rect 18414 24828 18420 24840
rect 18472 24828 18478 24880
rect 18877 24871 18935 24877
rect 18877 24837 18889 24871
rect 18923 24868 18935 24871
rect 20162 24868 20168 24880
rect 18923 24840 19334 24868
rect 18923 24837 18935 24840
rect 18877 24831 18935 24837
rect 16574 24800 16580 24812
rect 16040 24772 16580 24800
rect 16574 24760 16580 24772
rect 16632 24760 16638 24812
rect 17129 24803 17187 24809
rect 17129 24800 17141 24803
rect 16684 24772 17141 24800
rect 15289 24735 15347 24741
rect 15289 24701 15301 24735
rect 15335 24732 15347 24735
rect 15746 24732 15752 24744
rect 15335 24704 15752 24732
rect 15335 24701 15347 24704
rect 15289 24695 15347 24701
rect 15746 24692 15752 24704
rect 15804 24692 15810 24744
rect 15838 24692 15844 24744
rect 15896 24732 15902 24744
rect 16206 24732 16212 24744
rect 15896 24704 16212 24732
rect 15896 24692 15902 24704
rect 16206 24692 16212 24704
rect 16264 24732 16270 24744
rect 16684 24732 16712 24772
rect 17129 24769 17141 24772
rect 17175 24800 17187 24803
rect 17770 24800 17776 24812
rect 17175 24772 17776 24800
rect 17175 24769 17187 24772
rect 17129 24763 17187 24769
rect 17770 24760 17776 24772
rect 17828 24760 17834 24812
rect 19153 24803 19211 24809
rect 19153 24800 19165 24803
rect 18340 24772 19165 24800
rect 18340 24744 18368 24772
rect 19153 24769 19165 24772
rect 19199 24769 19211 24803
rect 19306 24800 19334 24840
rect 19812 24840 20168 24868
rect 19702 24800 19708 24812
rect 19306 24772 19708 24800
rect 19153 24763 19211 24769
rect 19702 24760 19708 24772
rect 19760 24800 19766 24812
rect 19812 24809 19840 24840
rect 20162 24828 20168 24840
rect 20220 24828 20226 24880
rect 22195 24868 22223 24908
rect 22370 24896 22376 24948
rect 22428 24936 22434 24948
rect 22557 24939 22615 24945
rect 22557 24936 22569 24939
rect 22428 24908 22569 24936
rect 22428 24896 22434 24908
rect 22557 24905 22569 24908
rect 22603 24905 22615 24939
rect 22557 24899 22615 24905
rect 25501 24939 25559 24945
rect 25501 24905 25513 24939
rect 25547 24936 25559 24939
rect 25590 24936 25596 24948
rect 25547 24908 25596 24936
rect 25547 24905 25559 24908
rect 25501 24899 25559 24905
rect 25590 24896 25596 24908
rect 25648 24896 25654 24948
rect 23014 24868 23020 24880
rect 22195 24840 22692 24868
rect 22927 24840 23020 24868
rect 19797 24803 19855 24809
rect 19797 24800 19809 24803
rect 19760 24772 19809 24800
rect 19760 24760 19766 24772
rect 19797 24769 19809 24772
rect 19843 24769 19855 24803
rect 19797 24763 19855 24769
rect 19889 24803 19947 24809
rect 19889 24769 19901 24803
rect 19935 24769 19947 24803
rect 20530 24800 20536 24812
rect 20491 24772 20536 24800
rect 19889 24763 19947 24769
rect 16850 24732 16856 24744
rect 16264 24704 16712 24732
rect 16811 24704 16856 24732
rect 16264 24692 16270 24704
rect 16850 24692 16856 24704
rect 16908 24692 16914 24744
rect 16945 24735 17003 24741
rect 16945 24701 16957 24735
rect 16991 24701 17003 24735
rect 16945 24695 17003 24701
rect 17037 24735 17095 24741
rect 17037 24701 17049 24735
rect 17083 24701 17095 24735
rect 17037 24695 17095 24701
rect 16482 24664 16488 24676
rect 15120 24636 16488 24664
rect 15120 24605 15148 24636
rect 16482 24624 16488 24636
rect 16540 24664 16546 24676
rect 16960 24664 16988 24695
rect 16540 24636 16988 24664
rect 16540 24624 16546 24636
rect 17052 24608 17080 24695
rect 17402 24692 17408 24744
rect 17460 24732 17466 24744
rect 18322 24732 18328 24744
rect 17460 24704 18328 24732
rect 17460 24692 17466 24704
rect 18322 24692 18328 24704
rect 18380 24692 18386 24744
rect 18414 24692 18420 24744
rect 18472 24732 18478 24744
rect 18601 24735 18659 24741
rect 18601 24732 18613 24735
rect 18472 24704 18613 24732
rect 18472 24692 18478 24704
rect 18601 24701 18613 24704
rect 18647 24732 18659 24735
rect 19904 24732 19932 24763
rect 20530 24760 20536 24772
rect 20588 24760 20594 24812
rect 20622 24760 20628 24812
rect 20680 24800 20686 24812
rect 21361 24803 21419 24809
rect 21361 24800 21373 24803
rect 20680 24772 21373 24800
rect 20680 24760 20686 24772
rect 21361 24769 21373 24772
rect 21407 24769 21419 24803
rect 21361 24763 21419 24769
rect 22186 24760 22192 24812
rect 22244 24800 22250 24812
rect 22244 24772 22289 24800
rect 22244 24760 22250 24772
rect 22370 24760 22376 24812
rect 22428 24800 22434 24812
rect 22664 24809 22692 24840
rect 23014 24828 23020 24840
rect 23072 24868 23078 24880
rect 28077 24871 28135 24877
rect 28077 24868 28089 24871
rect 23072 24840 28089 24868
rect 23072 24828 23078 24840
rect 28077 24837 28089 24840
rect 28123 24837 28135 24871
rect 28077 24831 28135 24837
rect 22465 24803 22523 24809
rect 22465 24800 22477 24803
rect 22428 24772 22477 24800
rect 22428 24760 22434 24772
rect 22465 24769 22477 24772
rect 22511 24769 22523 24803
rect 22465 24763 22523 24769
rect 22649 24803 22707 24809
rect 22649 24769 22661 24803
rect 22695 24800 22707 24803
rect 23569 24803 23627 24809
rect 23569 24800 23581 24803
rect 22695 24772 23581 24800
rect 22695 24769 22707 24772
rect 22649 24763 22707 24769
rect 23569 24769 23581 24772
rect 23615 24769 23627 24803
rect 23569 24763 23627 24769
rect 23753 24803 23811 24809
rect 23753 24769 23765 24803
rect 23799 24800 23811 24803
rect 24762 24800 24768 24812
rect 23799 24772 24768 24800
rect 23799 24769 23811 24772
rect 23753 24763 23811 24769
rect 24762 24760 24768 24772
rect 24820 24760 24826 24812
rect 25133 24803 25191 24809
rect 25133 24769 25145 24803
rect 25179 24800 25191 24803
rect 25682 24800 25688 24812
rect 25179 24772 25688 24800
rect 25179 24769 25191 24772
rect 25133 24763 25191 24769
rect 25682 24760 25688 24772
rect 25740 24760 25746 24812
rect 27801 24803 27859 24809
rect 27801 24769 27813 24803
rect 27847 24800 27859 24803
rect 28258 24800 28264 24812
rect 27847 24772 28264 24800
rect 27847 24769 27859 24772
rect 27801 24763 27859 24769
rect 28258 24760 28264 24772
rect 28316 24760 28322 24812
rect 20346 24732 20352 24744
rect 18647 24704 19932 24732
rect 19996 24704 20352 24732
rect 18647 24701 18659 24704
rect 18601 24695 18659 24701
rect 19521 24667 19579 24673
rect 19521 24633 19533 24667
rect 19567 24664 19579 24667
rect 19886 24664 19892 24676
rect 19567 24636 19892 24664
rect 19567 24633 19579 24636
rect 19521 24627 19579 24633
rect 19886 24624 19892 24636
rect 19944 24624 19950 24676
rect 15105 24599 15163 24605
rect 15105 24565 15117 24599
rect 15151 24565 15163 24599
rect 15105 24559 15163 24565
rect 15194 24556 15200 24608
rect 15252 24596 15258 24608
rect 16025 24599 16083 24605
rect 15252 24568 15297 24596
rect 15252 24556 15258 24568
rect 16025 24565 16037 24599
rect 16071 24596 16083 24599
rect 16669 24599 16727 24605
rect 16669 24596 16681 24599
rect 16071 24568 16681 24596
rect 16071 24565 16083 24568
rect 16025 24559 16083 24565
rect 16669 24565 16681 24568
rect 16715 24565 16727 24599
rect 16669 24559 16727 24565
rect 17034 24556 17040 24608
rect 17092 24556 17098 24608
rect 18598 24556 18604 24608
rect 18656 24596 18662 24608
rect 18877 24599 18935 24605
rect 18877 24596 18889 24599
rect 18656 24568 18889 24596
rect 18656 24556 18662 24568
rect 18877 24565 18889 24568
rect 18923 24565 18935 24599
rect 18877 24559 18935 24565
rect 19058 24556 19064 24608
rect 19116 24596 19122 24608
rect 19996 24596 20024 24704
rect 20346 24692 20352 24704
rect 20404 24692 20410 24744
rect 22097 24735 22155 24741
rect 22097 24701 22109 24735
rect 22143 24732 22155 24735
rect 25041 24735 25099 24741
rect 22143 24704 22232 24732
rect 22143 24701 22155 24704
rect 22097 24695 22155 24701
rect 22204 24664 22232 24704
rect 25041 24701 25053 24735
rect 25087 24732 25099 24735
rect 25087 24704 25176 24732
rect 25087 24701 25099 24704
rect 25041 24695 25099 24701
rect 25148 24676 25176 24704
rect 22462 24664 22468 24676
rect 22204 24636 22468 24664
rect 22462 24624 22468 24636
rect 22520 24664 22526 24676
rect 23014 24664 23020 24676
rect 22520 24636 23020 24664
rect 22520 24624 22526 24636
rect 23014 24624 23020 24636
rect 23072 24624 23078 24676
rect 25130 24624 25136 24676
rect 25188 24624 25194 24676
rect 20438 24596 20444 24608
rect 19116 24568 20024 24596
rect 20399 24568 20444 24596
rect 19116 24556 19122 24568
rect 20438 24556 20444 24568
rect 20496 24556 20502 24608
rect 21818 24596 21824 24608
rect 21779 24568 21824 24596
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 22002 24596 22008 24608
rect 21963 24568 22008 24596
rect 22002 24556 22008 24568
rect 22060 24596 22066 24608
rect 22370 24596 22376 24608
rect 22060 24568 22376 24596
rect 22060 24556 22066 24568
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 23661 24599 23719 24605
rect 23661 24565 23673 24599
rect 23707 24596 23719 24599
rect 23842 24596 23848 24608
rect 23707 24568 23848 24596
rect 23707 24565 23719 24568
rect 23661 24559 23719 24565
rect 23842 24556 23848 24568
rect 23900 24556 23906 24608
rect 1104 24506 28888 24528
rect 1104 24454 5582 24506
rect 5634 24454 5646 24506
rect 5698 24454 5710 24506
rect 5762 24454 5774 24506
rect 5826 24454 5838 24506
rect 5890 24454 14846 24506
rect 14898 24454 14910 24506
rect 14962 24454 14974 24506
rect 15026 24454 15038 24506
rect 15090 24454 15102 24506
rect 15154 24454 24110 24506
rect 24162 24454 24174 24506
rect 24226 24454 24238 24506
rect 24290 24454 24302 24506
rect 24354 24454 24366 24506
rect 24418 24454 28888 24506
rect 1104 24432 28888 24454
rect 13722 24392 13728 24404
rect 13683 24364 13728 24392
rect 13722 24352 13728 24364
rect 13780 24352 13786 24404
rect 15470 24352 15476 24404
rect 15528 24392 15534 24404
rect 16025 24395 16083 24401
rect 16025 24392 16037 24395
rect 15528 24364 16037 24392
rect 15528 24352 15534 24364
rect 16025 24361 16037 24364
rect 16071 24361 16083 24395
rect 16025 24355 16083 24361
rect 16209 24395 16267 24401
rect 16209 24361 16221 24395
rect 16255 24392 16267 24395
rect 16666 24392 16672 24404
rect 16255 24364 16672 24392
rect 16255 24361 16267 24364
rect 16209 24355 16267 24361
rect 15194 24284 15200 24336
rect 15252 24284 15258 24336
rect 15212 24256 15240 24284
rect 14936 24228 15240 24256
rect 12345 24191 12403 24197
rect 12345 24157 12357 24191
rect 12391 24188 12403 24191
rect 13814 24188 13820 24200
rect 12391 24160 13820 24188
rect 12391 24157 12403 24160
rect 12345 24151 12403 24157
rect 13814 24148 13820 24160
rect 13872 24188 13878 24200
rect 14734 24188 14740 24200
rect 13872 24160 14740 24188
rect 13872 24148 13878 24160
rect 14734 24148 14740 24160
rect 14792 24148 14798 24200
rect 14936 24197 14964 24228
rect 14921 24191 14979 24197
rect 14921 24157 14933 24191
rect 14967 24157 14979 24191
rect 14921 24151 14979 24157
rect 15197 24191 15255 24197
rect 15197 24157 15209 24191
rect 15243 24188 15255 24191
rect 15654 24188 15660 24200
rect 15243 24160 15660 24188
rect 15243 24157 15255 24160
rect 15197 24151 15255 24157
rect 15654 24148 15660 24160
rect 15712 24148 15718 24200
rect 16040 24188 16068 24355
rect 16666 24352 16672 24364
rect 16724 24352 16730 24404
rect 18141 24395 18199 24401
rect 18141 24361 18153 24395
rect 18187 24392 18199 24395
rect 18414 24392 18420 24404
rect 18187 24364 18420 24392
rect 18187 24361 18199 24364
rect 18141 24355 18199 24361
rect 18414 24352 18420 24364
rect 18472 24352 18478 24404
rect 18598 24392 18604 24404
rect 18559 24364 18604 24392
rect 18598 24352 18604 24364
rect 18656 24352 18662 24404
rect 20254 24352 20260 24404
rect 20312 24392 20318 24404
rect 20312 24364 20760 24392
rect 20312 24352 20318 24364
rect 18230 24284 18236 24336
rect 18288 24324 18294 24336
rect 20438 24324 20444 24336
rect 18288 24296 20444 24324
rect 18288 24284 18294 24296
rect 20438 24284 20444 24296
rect 20496 24284 20502 24336
rect 16206 24216 16212 24268
rect 16264 24256 16270 24268
rect 16485 24259 16543 24265
rect 16485 24256 16497 24259
rect 16264 24228 16497 24256
rect 16264 24216 16270 24228
rect 16485 24225 16497 24228
rect 16531 24256 16543 24259
rect 19702 24256 19708 24268
rect 16531 24228 17908 24256
rect 19663 24228 19708 24256
rect 16531 24225 16543 24228
rect 16485 24219 16543 24225
rect 16761 24191 16819 24197
rect 16761 24188 16773 24191
rect 15764 24160 16773 24188
rect 12612 24123 12670 24129
rect 12612 24089 12624 24123
rect 12658 24120 12670 24123
rect 12802 24120 12808 24132
rect 12658 24092 12808 24120
rect 12658 24089 12670 24092
rect 12612 24083 12670 24089
rect 12802 24080 12808 24092
rect 12860 24080 12866 24132
rect 14826 24080 14832 24132
rect 14884 24120 14890 24132
rect 15105 24123 15163 24129
rect 15105 24120 15117 24123
rect 14884 24092 15117 24120
rect 14884 24080 14890 24092
rect 15105 24089 15117 24092
rect 15151 24120 15163 24123
rect 15764 24120 15792 24160
rect 16761 24157 16773 24160
rect 16807 24188 16819 24191
rect 17034 24188 17040 24200
rect 16807 24160 17040 24188
rect 16807 24157 16819 24160
rect 16761 24151 16819 24157
rect 17034 24148 17040 24160
rect 17092 24148 17098 24200
rect 15151 24092 15792 24120
rect 15151 24089 15163 24092
rect 15105 24083 15163 24089
rect 15838 24080 15844 24132
rect 15896 24120 15902 24132
rect 16057 24123 16115 24129
rect 15896 24092 15941 24120
rect 15896 24080 15902 24092
rect 16057 24089 16069 24123
rect 16103 24120 16115 24123
rect 16666 24120 16672 24132
rect 16103 24092 16672 24120
rect 16103 24089 16115 24092
rect 16057 24083 16115 24089
rect 16666 24080 16672 24092
rect 16724 24080 16730 24132
rect 17586 24120 17592 24132
rect 17547 24092 17592 24120
rect 17586 24080 17592 24092
rect 17644 24080 17650 24132
rect 17770 24120 17776 24132
rect 17731 24092 17776 24120
rect 17770 24080 17776 24092
rect 17828 24080 17834 24132
rect 17880 24129 17908 24228
rect 19702 24216 19708 24228
rect 19760 24216 19766 24268
rect 20732 24265 20760 24364
rect 21082 24352 21088 24404
rect 21140 24392 21146 24404
rect 21545 24395 21603 24401
rect 21545 24392 21557 24395
rect 21140 24364 21557 24392
rect 21140 24352 21146 24364
rect 21545 24361 21557 24364
rect 21591 24361 21603 24395
rect 24949 24395 25007 24401
rect 24949 24392 24961 24395
rect 21545 24355 21603 24361
rect 22204 24364 24961 24392
rect 20717 24259 20775 24265
rect 20717 24225 20729 24259
rect 20763 24225 20775 24259
rect 20717 24219 20775 24225
rect 22204 24200 22232 24364
rect 24949 24361 24961 24364
rect 24995 24361 25007 24395
rect 24949 24355 25007 24361
rect 25593 24395 25651 24401
rect 25593 24361 25605 24395
rect 25639 24392 25651 24395
rect 25682 24392 25688 24404
rect 25639 24364 25688 24392
rect 25639 24361 25651 24364
rect 25593 24355 25651 24361
rect 24029 24327 24087 24333
rect 24029 24293 24041 24327
rect 24075 24324 24087 24327
rect 25608 24324 25636 24355
rect 25682 24352 25688 24364
rect 25740 24352 25746 24404
rect 25774 24352 25780 24404
rect 25832 24392 25838 24404
rect 26053 24395 26111 24401
rect 26053 24392 26065 24395
rect 25832 24364 26065 24392
rect 25832 24352 25838 24364
rect 26053 24361 26065 24364
rect 26099 24361 26111 24395
rect 26053 24355 26111 24361
rect 24075 24296 24716 24324
rect 24075 24293 24087 24296
rect 24029 24287 24087 24293
rect 18506 24188 18512 24200
rect 18467 24160 18512 24188
rect 18506 24148 18512 24160
rect 18564 24148 18570 24200
rect 18877 24191 18935 24197
rect 18877 24157 18889 24191
rect 18923 24188 18935 24191
rect 19242 24188 19248 24200
rect 18923 24160 19248 24188
rect 18923 24157 18935 24160
rect 18877 24151 18935 24157
rect 19242 24148 19248 24160
rect 19300 24148 19306 24200
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 20254 24188 20260 24200
rect 19475 24160 20260 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 20254 24148 20260 24160
rect 20312 24148 20318 24200
rect 20346 24148 20352 24200
rect 20404 24188 20410 24200
rect 20533 24191 20591 24197
rect 20533 24188 20545 24191
rect 20404 24160 20545 24188
rect 20404 24148 20410 24160
rect 20533 24157 20545 24160
rect 20579 24157 20591 24191
rect 20898 24188 20904 24200
rect 20859 24160 20904 24188
rect 20533 24151 20591 24157
rect 20898 24148 20904 24160
rect 20956 24148 20962 24200
rect 21266 24188 21272 24200
rect 21227 24160 21272 24188
rect 21266 24148 21272 24160
rect 21324 24148 21330 24200
rect 22002 24188 22008 24200
rect 21963 24160 22008 24188
rect 22002 24148 22008 24160
rect 22060 24148 22066 24200
rect 22186 24148 22192 24200
rect 22244 24188 22250 24200
rect 22646 24188 22652 24200
rect 22244 24160 22337 24188
rect 22607 24160 22652 24188
rect 22244 24148 22250 24160
rect 22646 24148 22652 24160
rect 22704 24148 22710 24200
rect 24688 24197 24716 24296
rect 25332 24296 25636 24324
rect 24765 24259 24823 24265
rect 24765 24225 24777 24259
rect 24811 24256 24823 24259
rect 25222 24256 25228 24268
rect 24811 24228 25228 24256
rect 24811 24225 24823 24228
rect 24765 24219 24823 24225
rect 25222 24216 25228 24228
rect 25280 24216 25286 24268
rect 24673 24191 24731 24197
rect 24673 24157 24685 24191
rect 24719 24188 24731 24191
rect 24854 24188 24860 24200
rect 24719 24160 24860 24188
rect 24719 24157 24731 24160
rect 24673 24151 24731 24157
rect 24854 24148 24860 24160
rect 24912 24148 24918 24200
rect 24949 24191 25007 24197
rect 24949 24157 24961 24191
rect 24995 24188 25007 24191
rect 25332 24188 25360 24296
rect 25406 24216 25412 24268
rect 25464 24256 25470 24268
rect 25501 24259 25559 24265
rect 25501 24256 25513 24259
rect 25464 24228 25513 24256
rect 25464 24216 25470 24228
rect 25501 24225 25513 24228
rect 25547 24256 25559 24259
rect 25547 24228 26096 24256
rect 25547 24225 25559 24228
rect 25501 24219 25559 24225
rect 26068 24197 26096 24228
rect 24995 24160 25360 24188
rect 25593 24191 25651 24197
rect 24995 24157 25007 24160
rect 24949 24151 25007 24157
rect 25593 24157 25605 24191
rect 25639 24157 25651 24191
rect 25593 24151 25651 24157
rect 26053 24191 26111 24197
rect 26053 24157 26065 24191
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 26237 24191 26295 24197
rect 26237 24157 26249 24191
rect 26283 24157 26295 24191
rect 26237 24151 26295 24157
rect 17865 24123 17923 24129
rect 17865 24089 17877 24123
rect 17911 24089 17923 24123
rect 18414 24120 18420 24132
rect 18375 24092 18420 24120
rect 17865 24083 17923 24089
rect 18414 24080 18420 24092
rect 18472 24080 18478 24132
rect 18785 24123 18843 24129
rect 18785 24089 18797 24123
rect 18831 24120 18843 24123
rect 18966 24120 18972 24132
rect 18831 24092 18972 24120
rect 18831 24089 18843 24092
rect 18785 24083 18843 24089
rect 18966 24080 18972 24092
rect 19024 24080 19030 24132
rect 22916 24123 22974 24129
rect 22916 24089 22928 24123
rect 22962 24120 22974 24123
rect 23290 24120 23296 24132
rect 22962 24092 23296 24120
rect 22962 24089 22974 24092
rect 22916 24083 22974 24089
rect 23290 24080 23296 24092
rect 23348 24080 23354 24132
rect 24581 24123 24639 24129
rect 24581 24089 24593 24123
rect 24627 24120 24639 24123
rect 24762 24120 24768 24132
rect 24627 24092 24768 24120
rect 24627 24089 24639 24092
rect 24581 24083 24639 24089
rect 24762 24080 24768 24092
rect 24820 24080 24826 24132
rect 25130 24080 25136 24132
rect 25188 24120 25194 24132
rect 25317 24123 25375 24129
rect 25317 24120 25329 24123
rect 25188 24092 25329 24120
rect 25188 24080 25194 24092
rect 25317 24089 25329 24092
rect 25363 24089 25375 24123
rect 25317 24083 25375 24089
rect 25608 24120 25636 24151
rect 26252 24120 26280 24151
rect 25608 24092 26280 24120
rect 14550 24012 14556 24064
rect 14608 24052 14614 24064
rect 14737 24055 14795 24061
rect 14737 24052 14749 24055
rect 14608 24024 14749 24052
rect 14608 24012 14614 24024
rect 14737 24021 14749 24024
rect 14783 24021 14795 24055
rect 15470 24052 15476 24064
rect 15431 24024 15476 24052
rect 14737 24015 14795 24021
rect 15470 24012 15476 24024
rect 15528 24012 15534 24064
rect 16684 24052 16712 24080
rect 17957 24055 18015 24061
rect 17957 24052 17969 24055
rect 16684 24024 17969 24052
rect 17957 24021 17969 24024
rect 18003 24021 18015 24055
rect 17957 24015 18015 24021
rect 22097 24055 22155 24061
rect 22097 24021 22109 24055
rect 22143 24052 22155 24055
rect 22370 24052 22376 24064
rect 22143 24024 22376 24052
rect 22143 24021 22155 24024
rect 22097 24015 22155 24021
rect 22370 24012 22376 24024
rect 22428 24012 22434 24064
rect 24486 24012 24492 24064
rect 24544 24052 24550 24064
rect 25608 24052 25636 24092
rect 25774 24052 25780 24064
rect 24544 24024 25636 24052
rect 25735 24024 25780 24052
rect 24544 24012 24550 24024
rect 25774 24012 25780 24024
rect 25832 24012 25838 24064
rect 1104 23962 28888 23984
rect 1104 23910 10214 23962
rect 10266 23910 10278 23962
rect 10330 23910 10342 23962
rect 10394 23910 10406 23962
rect 10458 23910 10470 23962
rect 10522 23910 19478 23962
rect 19530 23910 19542 23962
rect 19594 23910 19606 23962
rect 19658 23910 19670 23962
rect 19722 23910 19734 23962
rect 19786 23910 28888 23962
rect 1104 23888 28888 23910
rect 20346 23848 20352 23860
rect 15672 23820 20352 23848
rect 14476 23752 15424 23780
rect 14476 23721 14504 23752
rect 14461 23715 14519 23721
rect 14461 23681 14473 23715
rect 14507 23681 14519 23715
rect 14642 23712 14648 23724
rect 14603 23684 14648 23712
rect 14461 23675 14519 23681
rect 14642 23672 14648 23684
rect 14700 23672 14706 23724
rect 14737 23715 14795 23721
rect 14737 23681 14749 23715
rect 14783 23681 14795 23715
rect 14737 23675 14795 23681
rect 14752 23644 14780 23675
rect 14826 23672 14832 23724
rect 14884 23712 14890 23724
rect 15396 23721 15424 23752
rect 15381 23715 15439 23721
rect 14884 23684 14929 23712
rect 14884 23672 14890 23684
rect 15381 23681 15393 23715
rect 15427 23681 15439 23715
rect 15562 23712 15568 23724
rect 15523 23684 15568 23712
rect 15381 23675 15439 23681
rect 14476 23616 14780 23644
rect 15396 23644 15424 23675
rect 15562 23672 15568 23684
rect 15620 23672 15626 23724
rect 15672 23721 15700 23820
rect 20346 23808 20352 23820
rect 20404 23808 20410 23860
rect 23290 23848 23296 23860
rect 23251 23820 23296 23848
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 25222 23808 25228 23860
rect 25280 23848 25286 23860
rect 25958 23848 25964 23860
rect 25280 23820 25964 23848
rect 25280 23808 25286 23820
rect 25958 23808 25964 23820
rect 26016 23848 26022 23860
rect 26605 23851 26663 23857
rect 26605 23848 26617 23851
rect 26016 23820 26617 23848
rect 26016 23808 26022 23820
rect 26605 23817 26617 23820
rect 26651 23817 26663 23851
rect 26605 23811 26663 23817
rect 16482 23740 16488 23792
rect 16540 23780 16546 23792
rect 19334 23780 19340 23792
rect 16540 23752 16988 23780
rect 16540 23740 16546 23752
rect 15657 23715 15715 23721
rect 15657 23681 15669 23715
rect 15703 23681 15715 23715
rect 15657 23675 15715 23681
rect 15746 23672 15752 23724
rect 15804 23712 15810 23724
rect 16500 23712 16528 23740
rect 16666 23712 16672 23724
rect 15804 23684 16528 23712
rect 16627 23684 16672 23712
rect 15804 23672 15810 23684
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 16960 23721 16988 23752
rect 18156 23752 19340 23780
rect 18156 23724 18184 23752
rect 19334 23740 19340 23752
rect 19392 23780 19398 23792
rect 20438 23780 20444 23792
rect 19392 23752 20444 23780
rect 19392 23740 19398 23752
rect 20438 23740 20444 23752
rect 20496 23740 20502 23792
rect 20714 23740 20720 23792
rect 20772 23780 20778 23792
rect 20901 23783 20959 23789
rect 20901 23780 20913 23783
rect 20772 23752 20913 23780
rect 20772 23740 20778 23752
rect 20901 23749 20913 23752
rect 20947 23780 20959 23783
rect 22002 23780 22008 23792
rect 20947 23752 22008 23780
rect 20947 23749 20959 23752
rect 20901 23743 20959 23749
rect 22002 23740 22008 23752
rect 22060 23780 22066 23792
rect 24486 23780 24492 23792
rect 22060 23752 24492 23780
rect 22060 23740 22066 23752
rect 16945 23715 17003 23721
rect 16945 23681 16957 23715
rect 16991 23681 17003 23715
rect 18138 23712 18144 23724
rect 18051 23684 18144 23712
rect 16945 23675 17003 23681
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 18414 23721 18420 23724
rect 18408 23712 18420 23721
rect 18375 23684 18420 23712
rect 18408 23675 18420 23684
rect 18414 23672 18420 23675
rect 18472 23672 18478 23724
rect 19797 23715 19855 23721
rect 19797 23681 19809 23715
rect 19843 23712 19855 23715
rect 19978 23712 19984 23724
rect 19843 23684 19984 23712
rect 19843 23681 19855 23684
rect 19797 23675 19855 23681
rect 19978 23672 19984 23684
rect 20036 23672 20042 23724
rect 20349 23715 20407 23721
rect 20349 23681 20361 23715
rect 20395 23681 20407 23715
rect 20530 23712 20536 23724
rect 20491 23684 20536 23712
rect 20349 23675 20407 23681
rect 15470 23644 15476 23656
rect 15396 23616 15476 23644
rect 14476 23588 14504 23616
rect 15470 23604 15476 23616
rect 15528 23644 15534 23656
rect 20364 23644 20392 23675
rect 20530 23672 20536 23684
rect 20588 23672 20594 23724
rect 20993 23715 21051 23721
rect 20993 23681 21005 23715
rect 21039 23712 21051 23715
rect 21269 23715 21327 23721
rect 21269 23712 21281 23715
rect 21039 23684 21281 23712
rect 21039 23681 21051 23684
rect 20993 23675 21051 23681
rect 21269 23681 21281 23684
rect 21315 23681 21327 23715
rect 21269 23675 21327 23681
rect 21453 23715 21511 23721
rect 21453 23681 21465 23715
rect 21499 23712 21511 23715
rect 22186 23712 22192 23724
rect 21499 23684 22192 23712
rect 21499 23681 21511 23684
rect 21453 23675 21511 23681
rect 21008 23644 21036 23675
rect 15528 23616 16896 23644
rect 20364 23616 21036 23644
rect 21284 23644 21312 23675
rect 22186 23672 22192 23684
rect 22244 23672 22250 23724
rect 22940 23721 22968 23752
rect 24486 23740 24492 23752
rect 24544 23740 24550 23792
rect 24673 23783 24731 23789
rect 24673 23749 24685 23783
rect 24719 23780 24731 23783
rect 24762 23780 24768 23792
rect 24719 23752 24768 23780
rect 24719 23749 24731 23752
rect 24673 23743 24731 23749
rect 24762 23740 24768 23752
rect 24820 23740 24826 23792
rect 24854 23740 24860 23792
rect 24912 23780 24918 23792
rect 26142 23780 26148 23792
rect 24912 23752 26148 23780
rect 24912 23740 24918 23752
rect 26142 23740 26148 23752
rect 26200 23740 26206 23792
rect 22925 23715 22983 23721
rect 22925 23681 22937 23715
rect 22971 23681 22983 23715
rect 22925 23675 22983 23681
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23712 23443 23715
rect 23842 23712 23848 23724
rect 23431 23684 23704 23712
rect 23803 23684 23848 23712
rect 23431 23681 23443 23684
rect 23385 23675 23443 23681
rect 21726 23644 21732 23656
rect 21284 23616 21732 23644
rect 15528 23604 15534 23616
rect 14458 23536 14464 23588
rect 14516 23536 14522 23588
rect 16868 23520 16896 23616
rect 21726 23604 21732 23616
rect 21784 23644 21790 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21784 23616 21833 23644
rect 21784 23604 21790 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 22094 23644 22100 23656
rect 22055 23616 22100 23644
rect 21821 23607 21879 23613
rect 22094 23604 22100 23616
rect 22152 23604 22158 23656
rect 23676 23653 23704 23684
rect 23842 23672 23848 23684
rect 23900 23672 23906 23724
rect 24121 23715 24179 23721
rect 24121 23681 24133 23715
rect 24167 23712 24179 23715
rect 25038 23712 25044 23724
rect 24167 23684 25044 23712
rect 24167 23681 24179 23684
rect 24121 23675 24179 23681
rect 25038 23672 25044 23684
rect 25096 23672 25102 23724
rect 25498 23721 25504 23724
rect 25492 23675 25504 23721
rect 25556 23712 25562 23724
rect 27801 23715 27859 23721
rect 25556 23684 25592 23712
rect 25498 23672 25504 23675
rect 25556 23672 25562 23684
rect 27801 23681 27813 23715
rect 27847 23712 27859 23715
rect 28258 23712 28264 23724
rect 27847 23684 28264 23712
rect 27847 23681 27859 23684
rect 27801 23675 27859 23681
rect 28258 23672 28264 23684
rect 28316 23672 28322 23724
rect 23661 23647 23719 23653
rect 23661 23613 23673 23647
rect 23707 23613 23719 23647
rect 23661 23607 23719 23613
rect 23750 23604 23756 23656
rect 23808 23644 23814 23656
rect 23934 23644 23940 23656
rect 23808 23616 23940 23644
rect 23808 23604 23814 23616
rect 23934 23604 23940 23616
rect 23992 23604 23998 23656
rect 24029 23647 24087 23653
rect 24029 23613 24041 23647
rect 24075 23644 24087 23647
rect 24578 23644 24584 23656
rect 24075 23616 24584 23644
rect 24075 23613 24087 23616
rect 24029 23607 24087 23613
rect 24578 23604 24584 23616
rect 24636 23604 24642 23656
rect 25222 23644 25228 23656
rect 25183 23616 25228 23644
rect 25222 23604 25228 23616
rect 25280 23604 25286 23656
rect 19521 23579 19579 23585
rect 19521 23545 19533 23579
rect 19567 23576 19579 23579
rect 20254 23576 20260 23588
rect 19567 23548 20260 23576
rect 19567 23545 19579 23548
rect 19521 23539 19579 23545
rect 20254 23536 20260 23548
rect 20312 23536 20318 23588
rect 20346 23536 20352 23588
rect 20404 23576 20410 23588
rect 20533 23579 20591 23585
rect 20533 23576 20545 23579
rect 20404 23548 20545 23576
rect 20404 23536 20410 23548
rect 20533 23545 20545 23548
rect 20579 23545 20591 23579
rect 20533 23539 20591 23545
rect 20806 23536 20812 23588
rect 20864 23576 20870 23588
rect 21361 23579 21419 23585
rect 21361 23576 21373 23579
rect 20864 23548 21373 23576
rect 20864 23536 20870 23548
rect 21361 23545 21373 23548
rect 21407 23545 21419 23579
rect 21361 23539 21419 23545
rect 23201 23579 23259 23585
rect 23201 23545 23213 23579
rect 23247 23576 23259 23579
rect 24489 23579 24547 23585
rect 24489 23576 24501 23579
rect 23247 23548 24501 23576
rect 23247 23545 23259 23548
rect 23201 23539 23259 23545
rect 24489 23545 24501 23548
rect 24535 23576 24547 23579
rect 25130 23576 25136 23588
rect 24535 23548 25136 23576
rect 24535 23545 24547 23548
rect 24489 23539 24547 23545
rect 25130 23536 25136 23548
rect 25188 23536 25194 23588
rect 27982 23536 27988 23588
rect 28040 23576 28046 23588
rect 28077 23579 28135 23585
rect 28077 23576 28089 23579
rect 28040 23548 28089 23576
rect 28040 23536 28046 23548
rect 28077 23545 28089 23548
rect 28123 23545 28135 23579
rect 28077 23539 28135 23545
rect 1394 23508 1400 23520
rect 1355 23480 1400 23508
rect 1394 23468 1400 23480
rect 1452 23468 1458 23520
rect 14734 23468 14740 23520
rect 14792 23508 14798 23520
rect 15105 23511 15163 23517
rect 15105 23508 15117 23511
rect 14792 23480 15117 23508
rect 14792 23468 14798 23480
rect 15105 23477 15117 23480
rect 15151 23477 15163 23511
rect 15105 23471 15163 23477
rect 15930 23468 15936 23520
rect 15988 23508 15994 23520
rect 16025 23511 16083 23517
rect 16025 23508 16037 23511
rect 15988 23480 16037 23508
rect 15988 23468 15994 23480
rect 16025 23477 16037 23480
rect 16071 23477 16083 23511
rect 16025 23471 16083 23477
rect 16850 23468 16856 23520
rect 16908 23508 16914 23520
rect 17773 23511 17831 23517
rect 17773 23508 17785 23511
rect 16908 23480 17785 23508
rect 16908 23468 16914 23480
rect 17773 23477 17785 23480
rect 17819 23477 17831 23511
rect 17773 23471 17831 23477
rect 19889 23511 19947 23517
rect 19889 23477 19901 23511
rect 19935 23508 19947 23511
rect 20070 23508 20076 23520
rect 19935 23480 20076 23508
rect 19935 23477 19947 23480
rect 19889 23471 19947 23477
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 21910 23468 21916 23520
rect 21968 23508 21974 23520
rect 23063 23511 23121 23517
rect 23063 23508 23075 23511
rect 21968 23480 23075 23508
rect 21968 23468 21974 23480
rect 23063 23477 23075 23480
rect 23109 23477 23121 23511
rect 23063 23471 23121 23477
rect 1104 23418 28888 23440
rect 1104 23366 5582 23418
rect 5634 23366 5646 23418
rect 5698 23366 5710 23418
rect 5762 23366 5774 23418
rect 5826 23366 5838 23418
rect 5890 23366 14846 23418
rect 14898 23366 14910 23418
rect 14962 23366 14974 23418
rect 15026 23366 15038 23418
rect 15090 23366 15102 23418
rect 15154 23366 24110 23418
rect 24162 23366 24174 23418
rect 24226 23366 24238 23418
rect 24290 23366 24302 23418
rect 24354 23366 24366 23418
rect 24418 23366 28888 23418
rect 1104 23344 28888 23366
rect 12989 23307 13047 23313
rect 12989 23273 13001 23307
rect 13035 23304 13047 23307
rect 13814 23304 13820 23316
rect 13035 23276 13820 23304
rect 13035 23273 13047 23276
rect 12989 23267 13047 23273
rect 13814 23264 13820 23276
rect 13872 23264 13878 23316
rect 14642 23264 14648 23316
rect 14700 23304 14706 23316
rect 14737 23307 14795 23313
rect 14737 23304 14749 23307
rect 14700 23276 14749 23304
rect 14700 23264 14706 23276
rect 14737 23273 14749 23276
rect 14783 23273 14795 23307
rect 14737 23267 14795 23273
rect 15289 23307 15347 23313
rect 15289 23273 15301 23307
rect 15335 23304 15347 23307
rect 15562 23304 15568 23316
rect 15335 23276 15568 23304
rect 15335 23273 15347 23276
rect 15289 23267 15347 23273
rect 15562 23264 15568 23276
rect 15620 23264 15626 23316
rect 18138 23304 18144 23316
rect 15672 23276 18144 23304
rect 14458 23128 14464 23180
rect 14516 23168 14522 23180
rect 15672 23177 15700 23276
rect 18138 23264 18144 23276
rect 18196 23264 18202 23316
rect 18506 23264 18512 23316
rect 18564 23304 18570 23316
rect 18782 23304 18788 23316
rect 18564 23276 18788 23304
rect 18564 23264 18570 23276
rect 18782 23264 18788 23276
rect 18840 23264 18846 23316
rect 20530 23264 20536 23316
rect 20588 23304 20594 23316
rect 21085 23307 21143 23313
rect 21085 23304 21097 23307
rect 20588 23276 21097 23304
rect 20588 23264 20594 23276
rect 21085 23273 21097 23276
rect 21131 23304 21143 23307
rect 22462 23304 22468 23316
rect 21131 23276 22468 23304
rect 21131 23273 21143 23276
rect 21085 23267 21143 23273
rect 22462 23264 22468 23276
rect 22520 23264 22526 23316
rect 22646 23264 22652 23316
rect 22704 23304 22710 23316
rect 24581 23307 24639 23313
rect 24581 23304 24593 23307
rect 22704 23276 24593 23304
rect 22704 23264 22710 23276
rect 24581 23273 24593 23276
rect 24627 23304 24639 23307
rect 25222 23304 25228 23316
rect 24627 23276 25228 23304
rect 24627 23273 24639 23276
rect 24581 23267 24639 23273
rect 25222 23264 25228 23276
rect 25280 23264 25286 23316
rect 25409 23307 25467 23313
rect 25409 23273 25421 23307
rect 25455 23304 25467 23307
rect 25498 23304 25504 23316
rect 25455 23276 25504 23304
rect 25455 23273 25467 23276
rect 25409 23267 25467 23273
rect 25498 23264 25504 23276
rect 25556 23264 25562 23316
rect 16666 23196 16672 23248
rect 16724 23236 16730 23248
rect 17037 23239 17095 23245
rect 17037 23236 17049 23239
rect 16724 23208 17049 23236
rect 16724 23196 16730 23208
rect 17037 23205 17049 23208
rect 17083 23205 17095 23239
rect 17037 23199 17095 23205
rect 19521 23239 19579 23245
rect 19521 23205 19533 23239
rect 19567 23236 19579 23239
rect 19978 23236 19984 23248
rect 19567 23208 19984 23236
rect 19567 23205 19579 23208
rect 19521 23199 19579 23205
rect 15657 23171 15715 23177
rect 14516 23140 14872 23168
rect 14516 23128 14522 23140
rect 14550 23060 14556 23112
rect 14608 23100 14614 23112
rect 14844 23109 14872 23140
rect 15657 23137 15669 23171
rect 15703 23137 15715 23171
rect 15657 23131 15715 23137
rect 14645 23103 14703 23109
rect 14645 23100 14657 23103
rect 14608 23072 14657 23100
rect 14608 23060 14614 23072
rect 14645 23069 14657 23072
rect 14691 23069 14703 23103
rect 14645 23063 14703 23069
rect 14829 23103 14887 23109
rect 14829 23069 14841 23103
rect 14875 23100 14887 23103
rect 15197 23103 15255 23109
rect 15197 23100 15209 23103
rect 14875 23072 15209 23100
rect 14875 23069 14887 23072
rect 14829 23063 14887 23069
rect 15197 23069 15209 23072
rect 15243 23069 15255 23103
rect 15197 23063 15255 23069
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23100 15439 23103
rect 15746 23100 15752 23112
rect 15427 23072 15752 23100
rect 15427 23069 15439 23072
rect 15381 23063 15439 23069
rect 13081 23035 13139 23041
rect 13081 23001 13093 23035
rect 13127 23032 13139 23035
rect 13354 23032 13360 23044
rect 13127 23004 13360 23032
rect 13127 23001 13139 23004
rect 13081 22995 13139 23001
rect 13354 22992 13360 23004
rect 13412 22992 13418 23044
rect 15212 23032 15240 23063
rect 15746 23060 15752 23072
rect 15804 23060 15810 23112
rect 15930 23109 15936 23112
rect 15924 23100 15936 23109
rect 15891 23072 15936 23100
rect 15924 23063 15936 23072
rect 15930 23060 15936 23063
rect 15988 23060 15994 23112
rect 17052 23100 17080 23199
rect 19978 23196 19984 23208
rect 20036 23196 20042 23248
rect 23382 23236 23388 23248
rect 23343 23208 23388 23236
rect 23382 23196 23388 23208
rect 23440 23196 23446 23248
rect 23584 23208 24992 23236
rect 18233 23171 18291 23177
rect 18233 23137 18245 23171
rect 18279 23168 18291 23171
rect 18506 23168 18512 23180
rect 18279 23140 18512 23168
rect 18279 23137 18291 23140
rect 18233 23131 18291 23137
rect 18506 23128 18512 23140
rect 18564 23128 18570 23180
rect 20165 23171 20223 23177
rect 20165 23137 20177 23171
rect 20211 23168 20223 23171
rect 21818 23168 21824 23180
rect 20211 23140 21824 23168
rect 20211 23137 20223 23140
rect 20165 23131 20223 23137
rect 21818 23128 21824 23140
rect 21876 23128 21882 23180
rect 22281 23171 22339 23177
rect 22281 23137 22293 23171
rect 22327 23168 22339 23171
rect 23474 23168 23480 23180
rect 22327 23140 23480 23168
rect 22327 23137 22339 23140
rect 22281 23131 22339 23137
rect 23474 23128 23480 23140
rect 23532 23128 23538 23180
rect 18141 23103 18199 23109
rect 18141 23100 18153 23103
rect 17052 23072 18153 23100
rect 18141 23069 18153 23072
rect 18187 23069 18199 23103
rect 18966 23100 18972 23112
rect 18141 23063 18199 23069
rect 18248 23072 18972 23100
rect 18248 23032 18276 23072
rect 18966 23060 18972 23072
rect 19024 23060 19030 23112
rect 20438 23060 20444 23112
rect 20496 23100 20502 23112
rect 20717 23103 20775 23109
rect 20717 23100 20729 23103
rect 20496 23072 20729 23100
rect 20496 23060 20502 23072
rect 20717 23069 20729 23072
rect 20763 23069 20775 23103
rect 20717 23063 20775 23069
rect 21266 23060 21272 23112
rect 21324 23100 21330 23112
rect 21729 23103 21787 23109
rect 21729 23100 21741 23103
rect 21324 23072 21741 23100
rect 21324 23060 21330 23072
rect 21729 23069 21741 23072
rect 21775 23100 21787 23103
rect 21775 23072 22048 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 19680 23035 19738 23041
rect 19680 23032 19692 23035
rect 15212 23004 18276 23032
rect 18524 23004 19692 23032
rect 18524 22973 18552 23004
rect 19680 23001 19692 23004
rect 19726 23001 19738 23035
rect 20530 23032 20536 23044
rect 20491 23004 20536 23032
rect 19680 22995 19738 23001
rect 20530 22992 20536 23004
rect 20588 22992 20594 23044
rect 21910 23032 21916 23044
rect 21871 23004 21916 23032
rect 21910 22992 21916 23004
rect 21968 22992 21974 23044
rect 22020 23032 22048 23072
rect 22094 23060 22100 23112
rect 22152 23100 22158 23112
rect 22189 23103 22247 23109
rect 22189 23100 22201 23103
rect 22152 23072 22201 23100
rect 22152 23060 22158 23072
rect 22189 23069 22201 23072
rect 22235 23069 22247 23103
rect 22189 23063 22247 23069
rect 22373 23103 22431 23109
rect 22373 23069 22385 23103
rect 22419 23069 22431 23103
rect 22373 23063 22431 23069
rect 22388 23032 22416 23063
rect 22462 23060 22468 23112
rect 22520 23100 22526 23112
rect 23584 23100 23612 23208
rect 24964 23168 24992 23208
rect 25038 23196 25044 23248
rect 25096 23236 25102 23248
rect 26421 23239 26479 23245
rect 26421 23236 26433 23239
rect 25096 23208 26433 23236
rect 25096 23196 25102 23208
rect 26421 23205 26433 23208
rect 26467 23205 26479 23239
rect 26421 23199 26479 23205
rect 25593 23171 25651 23177
rect 25593 23168 25605 23171
rect 24964 23140 25605 23168
rect 25593 23137 25605 23140
rect 25639 23137 25651 23171
rect 25593 23131 25651 23137
rect 25774 23128 25780 23180
rect 25832 23168 25838 23180
rect 26053 23171 26111 23177
rect 26053 23168 26065 23171
rect 25832 23140 26065 23168
rect 25832 23128 25838 23140
rect 26053 23137 26065 23140
rect 26099 23137 26111 23171
rect 26053 23131 26111 23137
rect 22520 23072 23612 23100
rect 23661 23103 23719 23109
rect 22520 23060 22526 23072
rect 23661 23069 23673 23103
rect 23707 23100 23719 23103
rect 23750 23100 23756 23112
rect 23707 23072 23756 23100
rect 23707 23069 23719 23072
rect 23661 23063 23719 23069
rect 23750 23060 23756 23072
rect 23808 23060 23814 23112
rect 23934 23060 23940 23112
rect 23992 23100 23998 23112
rect 24949 23103 25007 23109
rect 24949 23100 24961 23103
rect 23992 23072 24961 23100
rect 23992 23060 23998 23072
rect 24949 23069 24961 23072
rect 24995 23069 25007 23103
rect 24949 23063 25007 23069
rect 25133 23103 25191 23109
rect 25133 23069 25145 23103
rect 25179 23100 25191 23103
rect 25498 23100 25504 23112
rect 25179 23072 25504 23100
rect 25179 23069 25191 23072
rect 25133 23063 25191 23069
rect 25498 23060 25504 23072
rect 25556 23060 25562 23112
rect 25685 23103 25743 23109
rect 25685 23069 25697 23103
rect 25731 23069 25743 23103
rect 25958 23100 25964 23112
rect 25919 23072 25964 23100
rect 25685 23063 25743 23069
rect 22922 23032 22928 23044
rect 22020 23004 22928 23032
rect 22922 22992 22928 23004
rect 22980 22992 22986 23044
rect 23385 23035 23443 23041
rect 23385 23001 23397 23035
rect 23431 23032 23443 23035
rect 24486 23032 24492 23044
rect 23431 23004 23704 23032
rect 24447 23004 24492 23032
rect 23431 23001 23443 23004
rect 23385 22995 23443 23001
rect 23676 22976 23704 23004
rect 24486 22992 24492 23004
rect 24544 22992 24550 23044
rect 25700 23032 25728 23063
rect 25958 23060 25964 23072
rect 26016 23060 26022 23112
rect 26142 23060 26148 23112
rect 26200 23100 26206 23112
rect 26329 23103 26387 23109
rect 26329 23100 26341 23103
rect 26200 23072 26341 23100
rect 26200 23060 26206 23072
rect 26329 23069 26341 23072
rect 26375 23069 26387 23103
rect 26329 23063 26387 23069
rect 25056 23004 25728 23032
rect 18509 22967 18567 22973
rect 18509 22933 18521 22967
rect 18555 22933 18567 22967
rect 18509 22927 18567 22933
rect 18598 22924 18604 22976
rect 18656 22964 18662 22976
rect 19797 22967 19855 22973
rect 19797 22964 19809 22967
rect 18656 22936 19809 22964
rect 18656 22924 18662 22936
rect 19797 22933 19809 22936
rect 19843 22933 19855 22967
rect 19797 22927 19855 22933
rect 19886 22924 19892 22976
rect 19944 22964 19950 22976
rect 19944 22936 19989 22964
rect 19944 22924 19950 22936
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 23569 22967 23627 22973
rect 23569 22964 23581 22967
rect 23532 22936 23581 22964
rect 23532 22924 23538 22936
rect 23569 22933 23581 22936
rect 23615 22933 23627 22967
rect 23569 22927 23627 22933
rect 23658 22924 23664 22976
rect 23716 22924 23722 22976
rect 24946 22924 24952 22976
rect 25004 22964 25010 22976
rect 25056 22973 25084 23004
rect 25041 22967 25099 22973
rect 25041 22964 25053 22967
rect 25004 22936 25053 22964
rect 25004 22924 25010 22936
rect 25041 22933 25053 22936
rect 25087 22933 25099 22967
rect 25041 22927 25099 22933
rect 1104 22874 28888 22896
rect 1104 22822 10214 22874
rect 10266 22822 10278 22874
rect 10330 22822 10342 22874
rect 10394 22822 10406 22874
rect 10458 22822 10470 22874
rect 10522 22822 19478 22874
rect 19530 22822 19542 22874
rect 19594 22822 19606 22874
rect 19658 22822 19670 22874
rect 19722 22822 19734 22874
rect 19786 22822 28888 22874
rect 1104 22800 28888 22822
rect 16206 22760 16212 22772
rect 16167 22732 16212 22760
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 17497 22763 17555 22769
rect 17497 22729 17509 22763
rect 17543 22760 17555 22763
rect 18598 22760 18604 22772
rect 17543 22732 18604 22760
rect 17543 22729 17555 22732
rect 17497 22723 17555 22729
rect 18598 22720 18604 22732
rect 18656 22720 18662 22772
rect 19797 22763 19855 22769
rect 19797 22729 19809 22763
rect 19843 22760 19855 22763
rect 19886 22760 19892 22772
rect 19843 22732 19892 22760
rect 19843 22729 19855 22732
rect 19797 22723 19855 22729
rect 19886 22720 19892 22732
rect 19944 22720 19950 22772
rect 23750 22760 23756 22772
rect 23711 22732 23756 22760
rect 23750 22720 23756 22732
rect 23808 22720 23814 22772
rect 23860 22732 24532 22760
rect 13814 22652 13820 22704
rect 13872 22692 13878 22704
rect 13872 22664 14596 22692
rect 13872 22652 13878 22664
rect 14568 22633 14596 22664
rect 14734 22652 14740 22704
rect 14792 22692 14798 22704
rect 15074 22695 15132 22701
rect 15074 22692 15086 22695
rect 14792 22664 15086 22692
rect 14792 22652 14798 22664
rect 15074 22661 15086 22664
rect 15120 22661 15132 22695
rect 20901 22695 20959 22701
rect 20901 22692 20913 22695
rect 15074 22655 15132 22661
rect 17052 22664 20913 22692
rect 14297 22627 14355 22633
rect 14297 22593 14309 22627
rect 14343 22624 14355 22627
rect 14553 22627 14611 22633
rect 14343 22596 14504 22624
rect 14343 22593 14355 22596
rect 14297 22587 14355 22593
rect 14476 22556 14504 22596
rect 14553 22593 14565 22627
rect 14599 22624 14611 22627
rect 14829 22627 14887 22633
rect 14829 22624 14841 22627
rect 14599 22596 14841 22624
rect 14599 22593 14611 22596
rect 14553 22587 14611 22593
rect 14829 22593 14841 22596
rect 14875 22593 14887 22627
rect 17052 22624 17080 22664
rect 20901 22661 20913 22664
rect 20947 22661 20959 22695
rect 22646 22692 22652 22704
rect 20901 22655 20959 22661
rect 22066 22664 22652 22692
rect 14829 22587 14887 22593
rect 14936 22596 17080 22624
rect 17129 22627 17187 22633
rect 14936 22556 14964 22596
rect 17129 22593 17141 22627
rect 17175 22624 17187 22627
rect 17770 22624 17776 22636
rect 17175 22596 17776 22624
rect 17175 22593 17187 22596
rect 17129 22587 17187 22593
rect 17770 22584 17776 22596
rect 17828 22584 17834 22636
rect 19429 22627 19487 22633
rect 19429 22593 19441 22627
rect 19475 22624 19487 22627
rect 20162 22624 20168 22636
rect 19475 22596 20168 22624
rect 19475 22593 19487 22596
rect 19429 22587 19487 22593
rect 20162 22584 20168 22596
rect 20220 22584 20226 22636
rect 20806 22624 20812 22636
rect 20767 22596 20812 22624
rect 20806 22584 20812 22596
rect 20864 22584 20870 22636
rect 20993 22627 21051 22633
rect 20993 22593 21005 22627
rect 21039 22624 21051 22627
rect 21818 22624 21824 22636
rect 21039 22596 21824 22624
rect 21039 22593 21051 22596
rect 20993 22587 21051 22593
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 21913 22627 21971 22633
rect 21913 22593 21925 22627
rect 21959 22624 21971 22627
rect 22066 22624 22094 22664
rect 22646 22652 22652 22664
rect 22704 22652 22710 22704
rect 21959 22596 22094 22624
rect 22180 22627 22238 22633
rect 21959 22593 21971 22596
rect 21913 22587 21971 22593
rect 22180 22593 22192 22627
rect 22226 22624 22238 22627
rect 23382 22624 23388 22636
rect 22226 22596 23388 22624
rect 22226 22593 22238 22596
rect 22180 22587 22238 22593
rect 23382 22584 23388 22596
rect 23440 22584 23446 22636
rect 14476 22528 14964 22556
rect 17221 22559 17279 22565
rect 17221 22525 17233 22559
rect 17267 22525 17279 22559
rect 19334 22556 19340 22568
rect 19295 22528 19340 22556
rect 17221 22519 17279 22525
rect 17236 22488 17264 22519
rect 19334 22516 19340 22528
rect 19392 22516 19398 22568
rect 22922 22516 22928 22568
rect 22980 22556 22986 22568
rect 23860 22556 23888 22732
rect 23934 22652 23940 22704
rect 23992 22692 23998 22704
rect 24397 22695 24455 22701
rect 24397 22692 24409 22695
rect 23992 22664 24409 22692
rect 23992 22652 23998 22664
rect 24397 22661 24409 22664
rect 24443 22661 24455 22695
rect 24504 22692 24532 22732
rect 24578 22720 24584 22772
rect 24636 22760 24642 22772
rect 25038 22760 25044 22772
rect 24636 22732 25044 22760
rect 24636 22720 24642 22732
rect 25038 22720 25044 22732
rect 25096 22760 25102 22772
rect 26145 22763 26203 22769
rect 26145 22760 26157 22763
rect 25096 22732 26157 22760
rect 25096 22720 25102 22732
rect 26145 22729 26157 22732
rect 26191 22729 26203 22763
rect 26145 22723 26203 22729
rect 25314 22692 25320 22704
rect 24504 22664 25320 22692
rect 24397 22655 24455 22661
rect 25314 22652 25320 22664
rect 25372 22652 25378 22704
rect 24210 22584 24216 22636
rect 24268 22624 24274 22636
rect 24673 22627 24731 22633
rect 24673 22624 24685 22627
rect 24268 22596 24685 22624
rect 24268 22584 24274 22596
rect 24673 22593 24685 22596
rect 24719 22593 24731 22627
rect 24673 22587 24731 22593
rect 24857 22627 24915 22633
rect 24857 22593 24869 22627
rect 24903 22593 24915 22627
rect 25590 22624 25596 22636
rect 25551 22596 25596 22624
rect 24857 22587 24915 22593
rect 22980 22528 23888 22556
rect 23937 22559 23995 22565
rect 22980 22516 22986 22528
rect 23937 22525 23949 22559
rect 23983 22525 23995 22559
rect 23937 22519 23995 22525
rect 24029 22559 24087 22565
rect 24029 22525 24041 22559
rect 24075 22525 24087 22559
rect 24029 22519 24087 22525
rect 19886 22488 19892 22500
rect 17236 22460 19892 22488
rect 19886 22448 19892 22460
rect 19944 22448 19950 22500
rect 23293 22491 23351 22497
rect 23293 22457 23305 22491
rect 23339 22488 23351 22491
rect 23566 22488 23572 22500
rect 23339 22460 23572 22488
rect 23339 22457 23351 22460
rect 23293 22451 23351 22457
rect 23566 22448 23572 22460
rect 23624 22488 23630 22500
rect 23842 22488 23848 22500
rect 23624 22460 23848 22488
rect 23624 22448 23630 22460
rect 23842 22448 23848 22460
rect 23900 22448 23906 22500
rect 11974 22380 11980 22432
rect 12032 22420 12038 22432
rect 12253 22423 12311 22429
rect 12253 22420 12265 22423
rect 12032 22392 12265 22420
rect 12032 22380 12038 22392
rect 12253 22389 12265 22392
rect 12299 22389 12311 22423
rect 12253 22383 12311 22389
rect 12526 22380 12532 22432
rect 12584 22420 12590 22432
rect 13173 22423 13231 22429
rect 13173 22420 13185 22423
rect 12584 22392 13185 22420
rect 12584 22380 12590 22392
rect 13173 22389 13185 22392
rect 13219 22389 13231 22423
rect 23952 22420 23980 22519
rect 24044 22488 24072 22519
rect 24578 22488 24584 22500
rect 24044 22460 24584 22488
rect 24578 22448 24584 22460
rect 24636 22488 24642 22500
rect 24673 22491 24731 22497
rect 24673 22488 24685 22491
rect 24636 22460 24685 22488
rect 24636 22448 24642 22460
rect 24673 22457 24685 22460
rect 24719 22457 24731 22491
rect 24673 22451 24731 22457
rect 24762 22448 24768 22500
rect 24820 22488 24826 22500
rect 24872 22488 24900 22587
rect 25590 22584 25596 22596
rect 25648 22624 25654 22636
rect 27246 22633 27252 22636
rect 26053 22627 26111 22633
rect 26053 22624 26065 22627
rect 25648 22596 26065 22624
rect 25648 22584 25654 22596
rect 26053 22593 26065 22596
rect 26099 22593 26111 22627
rect 26053 22587 26111 22593
rect 27240 22587 27252 22633
rect 27304 22624 27310 22636
rect 27304 22596 27340 22624
rect 27246 22584 27252 22587
rect 27304 22584 27310 22596
rect 25222 22516 25228 22568
rect 25280 22556 25286 22568
rect 26973 22559 27031 22565
rect 26973 22556 26985 22559
rect 25280 22528 26985 22556
rect 25280 22516 25286 22528
rect 26973 22525 26985 22528
rect 27019 22525 27031 22559
rect 26973 22519 27031 22525
rect 26050 22488 26056 22500
rect 24820 22460 26056 22488
rect 24820 22448 24826 22460
rect 26050 22448 26056 22460
rect 26108 22488 26114 22500
rect 26108 22460 26280 22488
rect 26108 22448 26114 22460
rect 25406 22420 25412 22432
rect 23952 22392 25412 22420
rect 13173 22383 13231 22389
rect 25406 22380 25412 22392
rect 25464 22380 25470 22432
rect 25498 22380 25504 22432
rect 25556 22420 25562 22432
rect 25866 22420 25872 22432
rect 25556 22392 25872 22420
rect 25556 22380 25562 22392
rect 25866 22380 25872 22392
rect 25924 22380 25930 22432
rect 26252 22420 26280 22460
rect 28353 22423 28411 22429
rect 28353 22420 28365 22423
rect 26252 22392 28365 22420
rect 28353 22389 28365 22392
rect 28399 22389 28411 22423
rect 28353 22383 28411 22389
rect 1104 22330 28888 22352
rect 1104 22278 5582 22330
rect 5634 22278 5646 22330
rect 5698 22278 5710 22330
rect 5762 22278 5774 22330
rect 5826 22278 5838 22330
rect 5890 22278 14846 22330
rect 14898 22278 14910 22330
rect 14962 22278 14974 22330
rect 15026 22278 15038 22330
rect 15090 22278 15102 22330
rect 15154 22278 24110 22330
rect 24162 22278 24174 22330
rect 24226 22278 24238 22330
rect 24290 22278 24302 22330
rect 24354 22278 24366 22330
rect 24418 22278 28888 22330
rect 1104 22256 28888 22278
rect 19613 22219 19671 22225
rect 19613 22185 19625 22219
rect 19659 22216 19671 22219
rect 23385 22219 23443 22225
rect 19659 22188 23336 22216
rect 19659 22185 19671 22188
rect 19613 22179 19671 22185
rect 17221 22151 17279 22157
rect 17221 22117 17233 22151
rect 17267 22148 17279 22151
rect 19058 22148 19064 22160
rect 17267 22120 19064 22148
rect 17267 22117 17279 22120
rect 17221 22111 17279 22117
rect 19058 22108 19064 22120
rect 19116 22108 19122 22160
rect 19978 22108 19984 22160
rect 20036 22108 20042 22160
rect 4430 22040 4436 22092
rect 4488 22080 4494 22092
rect 14182 22080 14188 22092
rect 4488 22052 14188 22080
rect 4488 22040 4494 22052
rect 14182 22040 14188 22052
rect 14240 22080 14246 22092
rect 14737 22083 14795 22089
rect 14737 22080 14749 22083
rect 14240 22052 14749 22080
rect 14240 22040 14246 22052
rect 14737 22049 14749 22052
rect 14783 22080 14795 22083
rect 16390 22080 16396 22092
rect 14783 22052 16396 22080
rect 14783 22049 14795 22052
rect 14737 22043 14795 22049
rect 16390 22040 16396 22052
rect 16448 22040 16454 22092
rect 16945 22083 17003 22089
rect 16945 22049 16957 22083
rect 16991 22080 17003 22083
rect 17402 22080 17408 22092
rect 16991 22052 17408 22080
rect 16991 22049 17003 22052
rect 16945 22043 17003 22049
rect 17402 22040 17408 22052
rect 17460 22040 17466 22092
rect 17770 22080 17776 22092
rect 17731 22052 17776 22080
rect 17770 22040 17776 22052
rect 17828 22040 17834 22092
rect 18046 22080 18052 22092
rect 18007 22052 18052 22080
rect 18046 22040 18052 22052
rect 18104 22040 18110 22092
rect 1394 22012 1400 22024
rect 1355 21984 1400 22012
rect 1394 21972 1400 21984
rect 1452 21972 1458 22024
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 22012 12219 22015
rect 13354 22012 13360 22024
rect 12207 21984 13360 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 21981 14151 22015
rect 14274 22012 14280 22024
rect 14235 21984 14280 22012
rect 14093 21975 14151 21981
rect 11974 21944 11980 21956
rect 11935 21916 11980 21944
rect 11974 21904 11980 21916
rect 12032 21904 12038 21956
rect 12710 21944 12716 21956
rect 12671 21916 12716 21944
rect 12710 21904 12716 21916
rect 12768 21904 12774 21956
rect 12897 21947 12955 21953
rect 12897 21913 12909 21947
rect 12943 21944 12955 21947
rect 13538 21944 13544 21956
rect 12943 21916 13544 21944
rect 12943 21913 12955 21916
rect 12897 21907 12955 21913
rect 13538 21904 13544 21916
rect 13596 21904 13602 21956
rect 12529 21879 12587 21885
rect 12529 21845 12541 21879
rect 12575 21876 12587 21879
rect 12618 21876 12624 21888
rect 12575 21848 12624 21876
rect 12575 21845 12587 21848
rect 12529 21839 12587 21845
rect 12618 21836 12624 21848
rect 12676 21836 12682 21888
rect 12728 21876 12756 21904
rect 14108 21876 14136 21975
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 15746 21972 15752 22024
rect 15804 22012 15810 22024
rect 15841 22015 15899 22021
rect 15841 22012 15853 22015
rect 15804 21984 15853 22012
rect 15804 21972 15810 21984
rect 15841 21981 15853 21984
rect 15887 21981 15899 22015
rect 15841 21975 15899 21981
rect 16206 21972 16212 22024
rect 16264 22012 16270 22024
rect 16853 22015 16911 22021
rect 16853 22012 16865 22015
rect 16264 21984 16865 22012
rect 16264 21972 16270 21984
rect 16853 21981 16865 21984
rect 16899 21981 16911 22015
rect 16853 21975 16911 21981
rect 17586 21972 17592 22024
rect 17644 22012 17650 22024
rect 17681 22015 17739 22021
rect 17681 22012 17693 22015
rect 17644 21984 17693 22012
rect 17644 21972 17650 21984
rect 17681 21981 17693 21984
rect 17727 21981 17739 22015
rect 17681 21975 17739 21981
rect 18874 21972 18880 22024
rect 18932 22012 18938 22024
rect 19996 22021 20024 22108
rect 23308 22080 23336 22188
rect 23385 22185 23397 22219
rect 23431 22216 23443 22219
rect 23474 22216 23480 22228
rect 23431 22188 23480 22216
rect 23431 22185 23443 22188
rect 23385 22179 23443 22185
rect 23474 22176 23480 22188
rect 23532 22176 23538 22228
rect 23937 22219 23995 22225
rect 23937 22185 23949 22219
rect 23983 22216 23995 22219
rect 24762 22216 24768 22228
rect 23983 22188 24768 22216
rect 23983 22185 23995 22188
rect 23937 22179 23995 22185
rect 24762 22176 24768 22188
rect 24820 22176 24826 22228
rect 27246 22216 27252 22228
rect 27207 22188 27252 22216
rect 27246 22176 27252 22188
rect 27304 22176 27310 22228
rect 24578 22148 24584 22160
rect 24412 22120 24584 22148
rect 24302 22080 24308 22092
rect 23308 22052 24308 22080
rect 19797 22015 19855 22021
rect 19797 22012 19809 22015
rect 18932 21984 19809 22012
rect 18932 21972 18938 21984
rect 19797 21981 19809 21984
rect 19843 21981 19855 22015
rect 19797 21975 19855 21981
rect 19889 22015 19947 22021
rect 19889 21981 19901 22015
rect 19935 21981 19947 22015
rect 19889 21975 19947 21981
rect 19981 22015 20039 22021
rect 19981 21981 19993 22015
rect 20027 21981 20039 22015
rect 19981 21975 20039 21981
rect 20073 22015 20131 22021
rect 20073 21981 20085 22015
rect 20119 21981 20131 22015
rect 20438 22012 20444 22024
rect 20399 21984 20444 22012
rect 20073 21975 20131 21981
rect 19904 21888 19932 21975
rect 12728 21848 14136 21876
rect 14366 21836 14372 21888
rect 14424 21876 14430 21888
rect 14461 21879 14519 21885
rect 14461 21876 14473 21879
rect 14424 21848 14473 21876
rect 14424 21836 14430 21848
rect 14461 21845 14473 21848
rect 14507 21845 14519 21879
rect 15654 21876 15660 21888
rect 15615 21848 15660 21876
rect 14461 21839 14519 21845
rect 15654 21836 15660 21848
rect 15712 21836 15718 21888
rect 16482 21836 16488 21888
rect 16540 21876 16546 21888
rect 19334 21876 19340 21888
rect 16540 21848 19340 21876
rect 16540 21836 16546 21848
rect 19334 21836 19340 21848
rect 19392 21836 19398 21888
rect 19886 21836 19892 21888
rect 19944 21836 19950 21888
rect 20088 21876 20116 21975
rect 20438 21972 20444 21984
rect 20496 21972 20502 22024
rect 23566 22012 23572 22024
rect 23527 21984 23572 22012
rect 23566 21972 23572 21984
rect 23624 21972 23630 22024
rect 23658 21972 23664 22024
rect 23716 22012 23722 22024
rect 23842 22012 23848 22024
rect 23716 21984 23848 22012
rect 23716 21972 23722 21984
rect 23842 21972 23848 21984
rect 23900 21972 23906 22024
rect 24044 22021 24072 22052
rect 24302 22040 24308 22052
rect 24360 22040 24366 22092
rect 24412 22021 24440 22120
rect 24578 22108 24584 22120
rect 24636 22108 24642 22160
rect 28350 22148 28356 22160
rect 28311 22120 28356 22148
rect 28350 22108 28356 22120
rect 28408 22108 28414 22160
rect 24946 22080 24952 22092
rect 24688 22052 24952 22080
rect 24688 22021 24716 22052
rect 24946 22040 24952 22052
rect 25004 22040 25010 22092
rect 25041 22083 25099 22089
rect 25041 22049 25053 22083
rect 25087 22080 25099 22083
rect 26050 22080 26056 22092
rect 25087 22052 25912 22080
rect 26011 22052 26056 22080
rect 25087 22049 25099 22052
rect 25041 22043 25099 22049
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 21981 24087 22015
rect 24029 21975 24087 21981
rect 24397 22015 24455 22021
rect 24673 22015 24731 22021
rect 24397 21981 24409 22015
rect 24443 21981 24455 22015
rect 24560 22009 24618 22015
rect 24560 22006 24572 22009
rect 24397 21975 24455 21981
rect 24504 21978 24572 22006
rect 20714 21953 20720 21956
rect 20708 21907 20720 21953
rect 20772 21944 20778 21956
rect 20772 21916 20808 21944
rect 20714 21904 20720 21907
rect 20772 21904 20778 21916
rect 24302 21904 24308 21956
rect 24360 21944 24366 21956
rect 24504 21944 24532 21978
rect 24560 21975 24572 21978
rect 24606 21975 24618 22009
rect 24673 21981 24685 22015
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 24765 22015 24823 22021
rect 24765 21981 24777 22015
rect 24811 22006 24823 22015
rect 24854 22006 24860 22024
rect 24811 21981 24860 22006
rect 24765 21978 24860 21981
rect 24765 21975 24823 21978
rect 24560 21969 24618 21975
rect 24854 21972 24860 21978
rect 24912 21972 24918 22024
rect 25498 21944 25504 21956
rect 24360 21916 24532 21944
rect 25459 21916 25504 21944
rect 24360 21904 24366 21916
rect 25498 21904 25504 21916
rect 25556 21904 25562 21956
rect 25884 21944 25912 22052
rect 26050 22040 26056 22052
rect 26108 22040 26114 22092
rect 26237 22083 26295 22089
rect 26237 22049 26249 22083
rect 26283 22080 26295 22083
rect 26881 22083 26939 22089
rect 26881 22080 26893 22083
rect 26283 22052 26893 22080
rect 26283 22049 26295 22052
rect 26237 22043 26295 22049
rect 26881 22049 26893 22052
rect 26927 22049 26939 22083
rect 26881 22043 26939 22049
rect 25958 21972 25964 22024
rect 26016 22012 26022 22024
rect 26513 22015 26571 22021
rect 26513 22012 26525 22015
rect 26016 21984 26525 22012
rect 26016 21972 26022 21984
rect 26513 21981 26525 21984
rect 26559 21981 26571 22015
rect 26513 21975 26571 21981
rect 26789 22015 26847 22021
rect 26789 21981 26801 22015
rect 26835 21981 26847 22015
rect 27062 22012 27068 22024
rect 27023 21984 27068 22012
rect 26789 21975 26847 21981
rect 26804 21944 26832 21975
rect 27062 21972 27068 21984
rect 27120 21972 27126 22024
rect 25884 21916 26832 21944
rect 21726 21876 21732 21888
rect 20088 21848 21732 21876
rect 21726 21836 21732 21848
rect 21784 21876 21790 21888
rect 21821 21879 21879 21885
rect 21821 21876 21833 21879
rect 21784 21848 21833 21876
rect 21784 21836 21790 21848
rect 21821 21845 21833 21848
rect 21867 21845 21879 21879
rect 21821 21839 21879 21845
rect 23474 21836 23480 21888
rect 23532 21876 23538 21888
rect 24670 21876 24676 21888
rect 23532 21848 24676 21876
rect 23532 21836 23538 21848
rect 24670 21836 24676 21848
rect 24728 21836 24734 21888
rect 25409 21879 25467 21885
rect 25409 21845 25421 21879
rect 25455 21876 25467 21879
rect 25958 21876 25964 21888
rect 25455 21848 25964 21876
rect 25455 21845 25467 21848
rect 25409 21839 25467 21845
rect 25958 21836 25964 21848
rect 26016 21836 26022 21888
rect 26421 21879 26479 21885
rect 26421 21845 26433 21879
rect 26467 21876 26479 21879
rect 26510 21876 26516 21888
rect 26467 21848 26516 21876
rect 26467 21845 26479 21848
rect 26421 21839 26479 21845
rect 26510 21836 26516 21848
rect 26568 21836 26574 21888
rect 1104 21786 28888 21808
rect 1104 21734 10214 21786
rect 10266 21734 10278 21786
rect 10330 21734 10342 21786
rect 10394 21734 10406 21786
rect 10458 21734 10470 21786
rect 10522 21734 19478 21786
rect 19530 21734 19542 21786
rect 19594 21734 19606 21786
rect 19658 21734 19670 21786
rect 19722 21734 19734 21786
rect 19786 21734 28888 21786
rect 1104 21712 28888 21734
rect 12710 21632 12716 21684
rect 12768 21672 12774 21684
rect 13633 21675 13691 21681
rect 13633 21672 13645 21675
rect 12768 21644 13645 21672
rect 12768 21632 12774 21644
rect 13633 21641 13645 21644
rect 13679 21641 13691 21675
rect 13998 21672 14004 21684
rect 13959 21644 14004 21672
rect 13633 21635 13691 21641
rect 13998 21632 14004 21644
rect 14056 21632 14062 21684
rect 19797 21675 19855 21681
rect 18432 21644 19380 21672
rect 13814 21604 13820 21616
rect 12268 21576 13820 21604
rect 11514 21428 11520 21480
rect 11572 21468 11578 21480
rect 12268 21477 12296 21576
rect 13814 21564 13820 21576
rect 13872 21604 13878 21616
rect 15096 21607 15154 21613
rect 13872 21576 14872 21604
rect 13872 21564 13878 21576
rect 12342 21496 12348 21548
rect 12400 21536 12406 21548
rect 12509 21539 12567 21545
rect 12509 21536 12521 21539
rect 12400 21508 12521 21536
rect 12400 21496 12406 21508
rect 12509 21505 12521 21508
rect 12555 21505 12567 21539
rect 12509 21499 12567 21505
rect 13998 21496 14004 21548
rect 14056 21536 14062 21548
rect 14185 21539 14243 21545
rect 14185 21536 14197 21539
rect 14056 21508 14197 21536
rect 14056 21496 14062 21508
rect 14185 21505 14197 21508
rect 14231 21505 14243 21539
rect 14366 21536 14372 21548
rect 14327 21508 14372 21536
rect 14185 21499 14243 21505
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 14844 21545 14872 21576
rect 15096 21573 15108 21607
rect 15142 21604 15154 21607
rect 15654 21604 15660 21616
rect 15142 21576 15660 21604
rect 15142 21573 15154 21576
rect 15096 21567 15154 21573
rect 15654 21564 15660 21576
rect 15712 21564 15718 21616
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21505 14887 21539
rect 14829 21499 14887 21505
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 17954 21536 17960 21548
rect 17819 21508 17960 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 17954 21496 17960 21508
rect 18012 21496 18018 21548
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 18233 21539 18291 21545
rect 18233 21536 18245 21539
rect 18104 21508 18245 21536
rect 18104 21496 18110 21508
rect 18233 21505 18245 21508
rect 18279 21505 18291 21539
rect 18233 21499 18291 21505
rect 18325 21539 18383 21545
rect 18325 21505 18337 21539
rect 18371 21536 18383 21539
rect 18432 21536 18460 21644
rect 18509 21607 18567 21613
rect 18509 21573 18521 21607
rect 18555 21604 18567 21607
rect 19352 21604 19380 21644
rect 19797 21641 19809 21675
rect 19843 21672 19855 21675
rect 19886 21672 19892 21684
rect 19843 21644 19892 21672
rect 19843 21641 19855 21644
rect 19797 21635 19855 21641
rect 19886 21632 19892 21644
rect 19944 21632 19950 21684
rect 21174 21632 21180 21684
rect 21232 21672 21238 21684
rect 23474 21672 23480 21684
rect 21232 21644 23480 21672
rect 21232 21632 21238 21644
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 24762 21672 24768 21684
rect 23860 21644 24768 21672
rect 20162 21604 20168 21616
rect 18555 21576 19196 21604
rect 18555 21573 18567 21576
rect 18509 21567 18567 21573
rect 19168 21548 19196 21576
rect 19352 21576 20168 21604
rect 18371 21508 18460 21536
rect 18601 21539 18659 21545
rect 18371 21505 18383 21508
rect 18325 21499 18383 21505
rect 18601 21505 18613 21539
rect 18647 21505 18659 21539
rect 18601 21499 18659 21505
rect 12253 21471 12311 21477
rect 12253 21468 12265 21471
rect 11572 21440 12265 21468
rect 11572 21428 11578 21440
rect 12253 21437 12265 21440
rect 12299 21437 12311 21471
rect 12253 21431 12311 21437
rect 14461 21471 14519 21477
rect 14461 21437 14473 21471
rect 14507 21437 14519 21471
rect 18616 21468 18644 21499
rect 18690 21496 18696 21548
rect 18748 21536 18754 21548
rect 19058 21536 19064 21548
rect 18748 21508 18793 21536
rect 19019 21508 19064 21536
rect 18748 21496 18754 21508
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 19150 21496 19156 21548
rect 19208 21536 19214 21548
rect 19352 21545 19380 21576
rect 20162 21564 20168 21576
rect 20220 21564 20226 21616
rect 20254 21564 20260 21616
rect 20312 21604 20318 21616
rect 20806 21604 20812 21616
rect 20312 21576 20576 21604
rect 20312 21564 20318 21576
rect 19245 21539 19303 21545
rect 19245 21536 19257 21539
rect 19208 21508 19257 21536
rect 19208 21496 19214 21508
rect 19245 21505 19257 21508
rect 19291 21505 19303 21539
rect 19245 21499 19303 21505
rect 19337 21539 19395 21545
rect 19337 21505 19349 21539
rect 19383 21505 19395 21539
rect 19337 21499 19395 21505
rect 19613 21539 19671 21545
rect 19613 21505 19625 21539
rect 19659 21536 19671 21539
rect 20070 21536 20076 21548
rect 19659 21508 20076 21536
rect 19659 21505 19671 21508
rect 19613 21499 19671 21505
rect 18785 21471 18843 21477
rect 18616 21440 18736 21468
rect 14461 21431 14519 21437
rect 14476 21332 14504 21431
rect 17218 21360 17224 21412
rect 17276 21400 17282 21412
rect 18708 21400 18736 21440
rect 18785 21437 18797 21471
rect 18831 21468 18843 21471
rect 18874 21468 18880 21480
rect 18831 21440 18880 21468
rect 18831 21437 18843 21440
rect 18785 21431 18843 21437
rect 18874 21428 18880 21440
rect 18932 21428 18938 21480
rect 19429 21471 19487 21477
rect 19429 21437 19441 21471
rect 19475 21468 19487 21471
rect 19518 21468 19524 21480
rect 19475 21440 19524 21468
rect 19475 21437 19487 21440
rect 19429 21431 19487 21437
rect 19518 21428 19524 21440
rect 19576 21428 19582 21480
rect 19628 21400 19656 21499
rect 20070 21496 20076 21508
rect 20128 21496 20134 21548
rect 20346 21536 20352 21548
rect 20307 21508 20352 21536
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 20548 21545 20576 21576
rect 20640 21576 20812 21604
rect 20640 21545 20668 21576
rect 20806 21564 20812 21576
rect 20864 21564 20870 21616
rect 23860 21604 23888 21644
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 23768 21576 23888 21604
rect 24029 21607 24087 21613
rect 20533 21539 20591 21545
rect 20533 21505 20545 21539
rect 20579 21505 20591 21539
rect 20533 21499 20591 21505
rect 20625 21539 20683 21545
rect 20625 21505 20637 21539
rect 20671 21505 20683 21539
rect 20625 21499 20683 21505
rect 20717 21539 20775 21545
rect 20717 21505 20729 21539
rect 20763 21536 20775 21539
rect 21910 21536 21916 21548
rect 20763 21508 21916 21536
rect 20763 21505 20775 21508
rect 20717 21499 20775 21505
rect 21910 21496 21916 21508
rect 21968 21496 21974 21548
rect 22094 21545 22100 21548
rect 22088 21499 22100 21545
rect 22152 21536 22158 21548
rect 23768 21545 23796 21576
rect 24029 21573 24041 21607
rect 24075 21604 24087 21607
rect 25406 21604 25412 21616
rect 24075 21576 24992 21604
rect 25367 21576 25412 21604
rect 24075 21573 24087 21576
rect 24029 21567 24087 21573
rect 23569 21539 23627 21545
rect 23569 21536 23581 21539
rect 22152 21508 22188 21536
rect 23216 21508 23581 21536
rect 22094 21496 22100 21499
rect 22152 21496 22158 21508
rect 20438 21428 20444 21480
rect 20496 21468 20502 21480
rect 21821 21471 21879 21477
rect 21821 21468 21833 21471
rect 20496 21440 21833 21468
rect 20496 21428 20502 21440
rect 21821 21437 21833 21440
rect 21867 21437 21879 21471
rect 21821 21431 21879 21437
rect 17276 21372 18644 21400
rect 18708 21372 19656 21400
rect 17276 21360 17282 21372
rect 15562 21332 15568 21344
rect 14476 21304 15568 21332
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 16209 21335 16267 21341
rect 16209 21301 16221 21335
rect 16255 21332 16267 21335
rect 16482 21332 16488 21344
rect 16255 21304 16488 21332
rect 16255 21301 16267 21304
rect 16209 21295 16267 21301
rect 16482 21292 16488 21304
rect 16540 21292 16546 21344
rect 17586 21332 17592 21344
rect 17547 21304 17592 21332
rect 17586 21292 17592 21304
rect 17644 21292 17650 21344
rect 18616 21332 18644 21372
rect 19886 21360 19892 21412
rect 19944 21400 19950 21412
rect 20622 21400 20628 21412
rect 19944 21372 20628 21400
rect 19944 21360 19950 21372
rect 20622 21360 20628 21372
rect 20680 21360 20686 21412
rect 20714 21360 20720 21412
rect 20772 21400 20778 21412
rect 20993 21403 21051 21409
rect 20993 21400 21005 21403
rect 20772 21372 21005 21400
rect 20772 21360 20778 21372
rect 20993 21369 21005 21372
rect 21039 21369 21051 21403
rect 20993 21363 21051 21369
rect 21174 21332 21180 21344
rect 18616 21304 21180 21332
rect 21174 21292 21180 21304
rect 21232 21292 21238 21344
rect 22186 21292 22192 21344
rect 22244 21332 22250 21344
rect 23216 21341 23244 21508
rect 23569 21505 23581 21508
rect 23615 21505 23627 21539
rect 23569 21499 23627 21505
rect 23753 21539 23811 21545
rect 23753 21505 23765 21539
rect 23799 21505 23811 21539
rect 23753 21499 23811 21505
rect 23845 21539 23903 21545
rect 23845 21505 23857 21539
rect 23891 21536 23903 21539
rect 23934 21536 23940 21548
rect 23891 21508 23940 21536
rect 23891 21505 23903 21508
rect 23845 21499 23903 21505
rect 23584 21468 23612 21499
rect 23934 21496 23940 21508
rect 23992 21496 23998 21548
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21536 24363 21539
rect 24762 21536 24768 21548
rect 24351 21508 24768 21536
rect 24351 21505 24363 21508
rect 24305 21499 24363 21505
rect 24762 21496 24768 21508
rect 24820 21496 24826 21548
rect 24964 21545 24992 21576
rect 25406 21564 25412 21576
rect 25464 21564 25470 21616
rect 25498 21564 25504 21616
rect 25556 21604 25562 21616
rect 25593 21607 25651 21613
rect 25593 21604 25605 21607
rect 25556 21576 25605 21604
rect 25556 21564 25562 21576
rect 25593 21573 25605 21576
rect 25639 21573 25651 21607
rect 25593 21567 25651 21573
rect 24949 21539 25007 21545
rect 24949 21505 24961 21539
rect 24995 21505 25007 21539
rect 24949 21499 25007 21505
rect 25038 21496 25044 21548
rect 25096 21536 25102 21548
rect 25133 21539 25191 21545
rect 25133 21536 25145 21539
rect 25096 21508 25145 21536
rect 25096 21496 25102 21508
rect 25133 21505 25145 21508
rect 25179 21536 25191 21539
rect 26142 21536 26148 21548
rect 25179 21508 26148 21536
rect 25179 21505 25191 21508
rect 25133 21499 25191 21505
rect 26142 21496 26148 21508
rect 26200 21496 26206 21548
rect 26418 21536 26424 21548
rect 26379 21508 26424 21536
rect 26418 21496 26424 21508
rect 26476 21496 26482 21548
rect 24397 21471 24455 21477
rect 24397 21468 24409 21471
rect 23584 21440 24409 21468
rect 24397 21437 24409 21440
rect 24443 21437 24455 21471
rect 24397 21431 24455 21437
rect 23658 21400 23664 21412
rect 23619 21372 23664 21400
rect 23658 21360 23664 21372
rect 23716 21360 23722 21412
rect 23842 21360 23848 21412
rect 23900 21400 23906 21412
rect 24949 21403 25007 21409
rect 24949 21400 24961 21403
rect 23900 21372 24961 21400
rect 23900 21360 23906 21372
rect 24949 21369 24961 21372
rect 24995 21369 25007 21403
rect 24949 21363 25007 21369
rect 23201 21335 23259 21341
rect 23201 21332 23213 21335
rect 22244 21304 23213 21332
rect 22244 21292 22250 21304
rect 23201 21301 23213 21304
rect 23247 21301 23259 21335
rect 23201 21295 23259 21301
rect 23566 21292 23572 21344
rect 23624 21332 23630 21344
rect 23934 21332 23940 21344
rect 23624 21304 23940 21332
rect 23624 21292 23630 21304
rect 23934 21292 23940 21304
rect 23992 21332 23998 21344
rect 24305 21335 24363 21341
rect 24305 21332 24317 21335
rect 23992 21304 24317 21332
rect 23992 21292 23998 21304
rect 24305 21301 24317 21304
rect 24351 21301 24363 21335
rect 24670 21332 24676 21344
rect 24631 21304 24676 21332
rect 24305 21295 24363 21301
rect 24670 21292 24676 21304
rect 24728 21292 24734 21344
rect 25866 21292 25872 21344
rect 25924 21332 25930 21344
rect 26050 21332 26056 21344
rect 25924 21304 26056 21332
rect 25924 21292 25930 21304
rect 26050 21292 26056 21304
rect 26108 21292 26114 21344
rect 26326 21332 26332 21344
rect 26287 21304 26332 21332
rect 26326 21292 26332 21304
rect 26384 21292 26390 21344
rect 28350 21332 28356 21344
rect 28311 21304 28356 21332
rect 28350 21292 28356 21304
rect 28408 21292 28414 21344
rect 1104 21242 28888 21264
rect 1104 21190 5582 21242
rect 5634 21190 5646 21242
rect 5698 21190 5710 21242
rect 5762 21190 5774 21242
rect 5826 21190 5838 21242
rect 5890 21190 14846 21242
rect 14898 21190 14910 21242
rect 14962 21190 14974 21242
rect 15026 21190 15038 21242
rect 15090 21190 15102 21242
rect 15154 21190 24110 21242
rect 24162 21190 24174 21242
rect 24226 21190 24238 21242
rect 24290 21190 24302 21242
rect 24354 21190 24366 21242
rect 24418 21190 28888 21242
rect 1104 21168 28888 21190
rect 12161 21131 12219 21137
rect 12161 21097 12173 21131
rect 12207 21128 12219 21131
rect 12342 21128 12348 21140
rect 12207 21100 12348 21128
rect 12207 21097 12219 21100
rect 12161 21091 12219 21097
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 15746 21128 15752 21140
rect 13188 21100 15608 21128
rect 15707 21100 15752 21128
rect 13188 21072 13216 21100
rect 11885 21063 11943 21069
rect 11885 21029 11897 21063
rect 11931 21060 11943 21063
rect 13170 21060 13176 21072
rect 11931 21032 13176 21060
rect 11931 21029 11943 21032
rect 11885 21023 11943 21029
rect 12360 20924 12388 21032
rect 13170 21020 13176 21032
rect 13228 21020 13234 21072
rect 13541 21063 13599 21069
rect 13541 21029 13553 21063
rect 13587 21060 13599 21063
rect 13814 21060 13820 21072
rect 13587 21032 13820 21060
rect 13587 21029 13599 21032
rect 13541 21023 13599 21029
rect 13814 21020 13820 21032
rect 13872 21020 13878 21072
rect 15580 21060 15608 21100
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 20346 21128 20352 21140
rect 17328 21100 20352 21128
rect 17129 21063 17187 21069
rect 17129 21060 17141 21063
rect 13924 21032 14504 21060
rect 15580 21032 17141 21060
rect 13924 20992 13952 21032
rect 12544 20964 13952 20992
rect 12544 20933 12572 20964
rect 12437 20927 12495 20933
rect 12437 20924 12449 20927
rect 12360 20896 12449 20924
rect 12437 20893 12449 20896
rect 12483 20893 12495 20927
rect 12437 20887 12495 20893
rect 12529 20927 12587 20933
rect 12529 20893 12541 20927
rect 12575 20893 12587 20927
rect 12529 20887 12587 20893
rect 12250 20816 12256 20868
rect 12308 20856 12314 20868
rect 12544 20856 12572 20887
rect 12618 20884 12624 20936
rect 12676 20924 12682 20936
rect 12805 20927 12863 20933
rect 12676 20896 12721 20924
rect 12676 20884 12682 20896
rect 12805 20893 12817 20927
rect 12851 20924 12863 20927
rect 12894 20924 12900 20936
rect 12851 20896 12900 20924
rect 12851 20893 12863 20896
rect 12805 20887 12863 20893
rect 12894 20884 12900 20896
rect 12952 20884 12958 20936
rect 13354 20924 13360 20936
rect 13315 20896 13360 20924
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 14182 20884 14188 20936
rect 14240 20918 14246 20936
rect 14476 20933 14504 21032
rect 17129 21029 17141 21032
rect 17175 21060 17187 21063
rect 17218 21060 17224 21072
rect 17175 21032 17224 21060
rect 17175 21029 17187 21032
rect 17129 21023 17187 21029
rect 17218 21020 17224 21032
rect 17276 21020 17282 21072
rect 15013 20995 15071 21001
rect 15013 20992 15025 20995
rect 14568 20964 15025 20992
rect 14568 20933 14596 20964
rect 15013 20961 15025 20964
rect 15059 20961 15071 20995
rect 17328 20992 17356 21100
rect 20346 21088 20352 21100
rect 20404 21088 20410 21140
rect 22094 21088 22100 21140
rect 22152 21128 22158 21140
rect 22281 21131 22339 21137
rect 22281 21128 22293 21131
rect 22152 21100 22293 21128
rect 22152 21088 22158 21100
rect 22281 21097 22293 21100
rect 22327 21097 22339 21131
rect 22281 21091 22339 21097
rect 22649 21131 22707 21137
rect 22649 21097 22661 21131
rect 22695 21128 22707 21131
rect 23842 21128 23848 21140
rect 22695 21100 23848 21128
rect 22695 21097 22707 21100
rect 22649 21091 22707 21097
rect 23842 21088 23848 21100
rect 23900 21088 23906 21140
rect 24029 21131 24087 21137
rect 24029 21097 24041 21131
rect 24075 21128 24087 21131
rect 24670 21128 24676 21140
rect 24075 21100 24532 21128
rect 24631 21100 24676 21128
rect 24075 21097 24087 21100
rect 24029 21091 24087 21097
rect 18877 21063 18935 21069
rect 18877 21029 18889 21063
rect 18923 21060 18935 21063
rect 19518 21060 19524 21072
rect 18923 21032 19524 21060
rect 18923 21029 18935 21032
rect 18877 21023 18935 21029
rect 19518 21020 19524 21032
rect 19576 21020 19582 21072
rect 20070 21020 20076 21072
rect 20128 21060 20134 21072
rect 20990 21060 20996 21072
rect 20128 21032 20996 21060
rect 20128 21020 20134 21032
rect 20990 21020 20996 21032
rect 21048 21060 21054 21072
rect 21269 21063 21327 21069
rect 21269 21060 21281 21063
rect 21048 21032 21281 21060
rect 21048 21020 21054 21032
rect 21269 21029 21281 21032
rect 21315 21029 21327 21063
rect 21269 21023 21327 21029
rect 21818 21020 21824 21072
rect 21876 21060 21882 21072
rect 22741 21063 22799 21069
rect 22741 21060 22753 21063
rect 21876 21032 22753 21060
rect 21876 21020 21882 21032
rect 22741 21029 22753 21032
rect 22787 21029 22799 21063
rect 22741 21023 22799 21029
rect 23385 21063 23443 21069
rect 23385 21029 23397 21063
rect 23431 21060 23443 21063
rect 24394 21060 24400 21072
rect 23431 21032 24400 21060
rect 23431 21029 23443 21032
rect 23385 21023 23443 21029
rect 24394 21020 24400 21032
rect 24452 21020 24458 21072
rect 24504 21060 24532 21100
rect 24670 21088 24676 21100
rect 24728 21088 24734 21140
rect 25056 21100 26556 21128
rect 24854 21060 24860 21072
rect 24504 21032 24860 21060
rect 24854 21020 24860 21032
rect 24912 21020 24918 21072
rect 15013 20955 15071 20961
rect 15111 20964 17356 20992
rect 14349 20927 14407 20933
rect 14349 20918 14361 20927
rect 14240 20893 14361 20918
rect 14395 20924 14407 20927
rect 14461 20927 14519 20933
rect 14395 20893 14412 20924
rect 14240 20890 14412 20893
rect 14461 20893 14473 20927
rect 14507 20893 14519 20927
rect 14240 20884 14246 20890
rect 14349 20887 14407 20890
rect 14461 20887 14519 20893
rect 14553 20927 14611 20933
rect 14553 20893 14565 20927
rect 14599 20893 14611 20927
rect 14553 20887 14611 20893
rect 14734 20884 14740 20936
rect 14792 20924 14798 20936
rect 15111 20924 15139 20964
rect 20254 20952 20260 21004
rect 20312 20992 20318 21004
rect 21358 20992 21364 21004
rect 20312 20964 21364 20992
rect 20312 20952 20318 20964
rect 15930 20924 15936 20936
rect 14792 20896 15139 20924
rect 15891 20896 15936 20924
rect 14792 20884 14798 20896
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 16117 20927 16175 20933
rect 16117 20893 16129 20927
rect 16163 20893 16175 20927
rect 16390 20924 16396 20936
rect 16351 20896 16396 20924
rect 16117 20887 16175 20893
rect 15194 20856 15200 20868
rect 12308 20828 12572 20856
rect 15155 20828 15200 20856
rect 12308 20816 12314 20828
rect 15194 20816 15200 20828
rect 15252 20816 15258 20868
rect 15286 20816 15292 20868
rect 15344 20856 15350 20868
rect 15381 20859 15439 20865
rect 15381 20856 15393 20859
rect 15344 20828 15393 20856
rect 15344 20816 15350 20828
rect 15381 20825 15393 20828
rect 15427 20825 15439 20859
rect 16132 20856 16160 20887
rect 16390 20884 16396 20896
rect 16448 20884 16454 20936
rect 17494 20924 17500 20936
rect 17455 20896 17500 20924
rect 17494 20884 17500 20896
rect 17552 20884 17558 20936
rect 17586 20884 17592 20936
rect 17644 20924 17650 20936
rect 17753 20927 17811 20933
rect 17753 20924 17765 20927
rect 17644 20896 17765 20924
rect 17644 20884 17650 20896
rect 17753 20893 17765 20896
rect 17799 20893 17811 20927
rect 19518 20924 19524 20936
rect 19479 20896 19524 20924
rect 17753 20887 17811 20893
rect 19518 20884 19524 20896
rect 19576 20884 19582 20936
rect 20622 20924 20628 20936
rect 20583 20896 20628 20924
rect 20622 20884 20628 20896
rect 20680 20884 20686 20936
rect 20732 20933 20760 20964
rect 21358 20952 21364 20964
rect 21416 20992 21422 21004
rect 21928 20992 22068 21000
rect 22833 20995 22891 21001
rect 22833 20992 22845 20995
rect 21416 20972 22845 20992
rect 21416 20964 21956 20972
rect 22040 20964 22845 20972
rect 21416 20952 21422 20964
rect 20717 20927 20775 20933
rect 20717 20893 20729 20927
rect 20763 20893 20775 20927
rect 20717 20887 20775 20893
rect 20806 20884 20812 20936
rect 20864 20924 20870 20936
rect 20864 20896 20909 20924
rect 20864 20884 20870 20896
rect 20990 20884 20996 20936
rect 21048 20924 21054 20936
rect 21637 20927 21695 20933
rect 21637 20924 21649 20927
rect 21048 20896 21649 20924
rect 21048 20884 21054 20896
rect 21637 20893 21649 20896
rect 21683 20893 21695 20927
rect 21818 20924 21824 20936
rect 21779 20896 21824 20924
rect 21637 20887 21695 20893
rect 21818 20884 21824 20896
rect 21876 20884 21882 20936
rect 21928 20933 21956 20964
rect 22833 20961 22845 20964
rect 22879 20992 22891 20995
rect 23106 20992 23112 21004
rect 22879 20964 23112 20992
rect 22879 20961 22891 20964
rect 22833 20955 22891 20961
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 24670 20992 24676 21004
rect 24044 20964 24676 20992
rect 21913 20927 21971 20933
rect 21913 20893 21925 20927
rect 21959 20893 21971 20927
rect 21913 20887 21971 20893
rect 22051 20927 22109 20933
rect 22051 20893 22063 20927
rect 22097 20926 22109 20927
rect 22097 20924 22131 20926
rect 22186 20924 22192 20936
rect 22097 20896 22192 20924
rect 22097 20893 22109 20896
rect 22051 20887 22109 20893
rect 22186 20884 22192 20896
rect 22244 20884 22250 20936
rect 22554 20924 22560 20936
rect 22515 20896 22560 20924
rect 22554 20884 22560 20896
rect 22612 20884 22618 20936
rect 23658 20884 23664 20936
rect 23716 20924 23722 20936
rect 23842 20924 23848 20936
rect 23716 20896 23848 20924
rect 23716 20884 23722 20896
rect 23842 20884 23848 20896
rect 23900 20884 23906 20936
rect 24044 20933 24072 20964
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 24029 20927 24087 20933
rect 24029 20893 24041 20927
rect 24075 20893 24087 20927
rect 24762 20924 24768 20936
rect 24723 20896 24768 20924
rect 24029 20887 24087 20893
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 24857 20927 24915 20933
rect 24857 20893 24869 20927
rect 24903 20924 24915 20927
rect 24946 20924 24952 20936
rect 24903 20896 24952 20924
rect 24903 20893 24915 20896
rect 24857 20887 24915 20893
rect 24946 20884 24952 20896
rect 25004 20884 25010 20936
rect 18322 20856 18328 20868
rect 16132 20828 18328 20856
rect 15381 20819 15439 20825
rect 18322 20816 18328 20828
rect 18380 20816 18386 20868
rect 20438 20856 20444 20868
rect 19628 20828 20444 20856
rect 14090 20788 14096 20800
rect 14051 20760 14096 20788
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 16850 20788 16856 20800
rect 16763 20760 16856 20788
rect 16850 20748 16856 20760
rect 16908 20788 16914 20800
rect 17126 20788 17132 20800
rect 16908 20760 17132 20788
rect 16908 20748 16914 20760
rect 17126 20748 17132 20760
rect 17184 20748 17190 20800
rect 18690 20748 18696 20800
rect 18748 20788 18754 20800
rect 19628 20797 19656 20828
rect 20438 20816 20444 20828
rect 20496 20816 20502 20868
rect 23198 20856 23204 20868
rect 23159 20828 23204 20856
rect 23198 20816 23204 20828
rect 23256 20816 23262 20868
rect 23290 20816 23296 20868
rect 23348 20856 23354 20868
rect 25056 20856 25084 21100
rect 26326 21060 26332 21072
rect 25792 21032 26332 21060
rect 25225 20995 25283 21001
rect 25225 20961 25237 20995
rect 25271 20992 25283 20995
rect 25682 20992 25688 21004
rect 25271 20964 25688 20992
rect 25271 20961 25283 20964
rect 25225 20955 25283 20961
rect 25682 20952 25688 20964
rect 25740 20952 25746 21004
rect 25792 21001 25820 21032
rect 26326 21020 26332 21032
rect 26384 21020 26390 21072
rect 25777 20995 25835 21001
rect 25777 20961 25789 20995
rect 25823 20961 25835 20995
rect 25777 20955 25835 20961
rect 26145 20995 26203 21001
rect 26145 20961 26157 20995
rect 26191 20992 26203 20995
rect 26191 20964 26464 20992
rect 26191 20961 26203 20964
rect 26145 20955 26203 20961
rect 25314 20924 25320 20936
rect 25227 20896 25320 20924
rect 25314 20884 25320 20896
rect 25372 20924 25378 20936
rect 25866 20924 25872 20936
rect 25372 20896 25728 20924
rect 25827 20896 25872 20924
rect 25372 20884 25378 20896
rect 23348 20828 25084 20856
rect 25700 20856 25728 20896
rect 25866 20884 25872 20896
rect 25924 20884 25930 20936
rect 25961 20927 26019 20933
rect 25961 20893 25973 20927
rect 26007 20924 26019 20927
rect 26050 20924 26056 20936
rect 26007 20896 26056 20924
rect 26007 20893 26019 20896
rect 25961 20887 26019 20893
rect 26050 20884 26056 20896
rect 26108 20884 26114 20936
rect 26436 20933 26464 20964
rect 26528 20933 26556 21100
rect 26697 21063 26755 21069
rect 26697 21029 26709 21063
rect 26743 21029 26755 21063
rect 26697 21023 26755 21029
rect 26712 20992 26740 21023
rect 26712 20964 27108 20992
rect 26421 20927 26479 20933
rect 26421 20893 26433 20927
rect 26467 20893 26479 20927
rect 26421 20887 26479 20893
rect 26513 20927 26571 20933
rect 26513 20893 26525 20927
rect 26559 20893 26571 20927
rect 26513 20887 26571 20893
rect 26602 20884 26608 20936
rect 26660 20924 26666 20936
rect 26697 20927 26755 20933
rect 26697 20924 26709 20927
rect 26660 20896 26709 20924
rect 26660 20884 26666 20896
rect 26697 20893 26709 20896
rect 26743 20893 26755 20927
rect 26697 20887 26755 20893
rect 26878 20884 26884 20936
rect 26936 20924 26942 20936
rect 26973 20927 27031 20933
rect 26973 20924 26985 20927
rect 26936 20896 26985 20924
rect 26936 20884 26942 20896
rect 26973 20893 26985 20896
rect 27019 20893 27031 20927
rect 27080 20924 27108 20964
rect 27229 20927 27287 20933
rect 27229 20924 27241 20927
rect 27080 20896 27241 20924
rect 26973 20887 27031 20893
rect 27229 20893 27241 20896
rect 27275 20893 27287 20927
rect 27229 20887 27287 20893
rect 25700 20828 28396 20856
rect 23348 20816 23354 20828
rect 19613 20791 19671 20797
rect 19613 20788 19625 20791
rect 18748 20760 19625 20788
rect 18748 20748 18754 20760
rect 19613 20757 19625 20760
rect 19659 20757 19671 20791
rect 20070 20788 20076 20800
rect 20031 20760 20076 20788
rect 19613 20751 19671 20757
rect 20070 20748 20076 20760
rect 20128 20748 20134 20800
rect 20346 20788 20352 20800
rect 20307 20760 20352 20788
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 24489 20791 24547 20797
rect 24489 20757 24501 20791
rect 24535 20788 24547 20791
rect 25222 20788 25228 20800
rect 24535 20760 25228 20788
rect 24535 20757 24547 20760
rect 24489 20751 24547 20757
rect 25222 20748 25228 20760
rect 25280 20748 25286 20800
rect 28368 20797 28396 20828
rect 28353 20791 28411 20797
rect 28353 20757 28365 20791
rect 28399 20757 28411 20791
rect 28353 20751 28411 20757
rect 1104 20698 28888 20720
rect 1104 20646 10214 20698
rect 10266 20646 10278 20698
rect 10330 20646 10342 20698
rect 10394 20646 10406 20698
rect 10458 20646 10470 20698
rect 10522 20646 19478 20698
rect 19530 20646 19542 20698
rect 19594 20646 19606 20698
rect 19658 20646 19670 20698
rect 19722 20646 19734 20698
rect 19786 20646 28888 20698
rect 1104 20624 28888 20646
rect 12897 20587 12955 20593
rect 12897 20553 12909 20587
rect 12943 20584 12955 20587
rect 13078 20584 13084 20596
rect 12943 20556 13084 20584
rect 12943 20553 12955 20556
rect 12897 20547 12955 20553
rect 13078 20544 13084 20556
rect 13136 20584 13142 20596
rect 15286 20584 15292 20596
rect 13136 20556 13400 20584
rect 13136 20544 13142 20556
rect 13372 20525 13400 20556
rect 13556 20556 15292 20584
rect 13556 20528 13584 20556
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 15930 20544 15936 20596
rect 15988 20584 15994 20596
rect 16301 20587 16359 20593
rect 16301 20584 16313 20587
rect 15988 20556 16313 20584
rect 15988 20544 15994 20556
rect 16301 20553 16313 20556
rect 16347 20553 16359 20587
rect 16301 20547 16359 20553
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18049 20587 18107 20593
rect 18049 20584 18061 20587
rect 18012 20556 18061 20584
rect 18012 20544 18018 20556
rect 18049 20553 18061 20556
rect 18095 20553 18107 20587
rect 18049 20547 18107 20553
rect 20622 20544 20628 20596
rect 20680 20584 20686 20596
rect 21453 20587 21511 20593
rect 21453 20584 21465 20587
rect 20680 20556 21465 20584
rect 20680 20544 20686 20556
rect 21453 20553 21465 20556
rect 21499 20584 21511 20587
rect 23658 20584 23664 20596
rect 21499 20556 23664 20584
rect 21499 20553 21511 20556
rect 21453 20547 21511 20553
rect 23658 20544 23664 20556
rect 23716 20544 23722 20596
rect 25866 20544 25872 20596
rect 25924 20584 25930 20596
rect 26345 20587 26403 20593
rect 26345 20584 26357 20587
rect 25924 20556 26357 20584
rect 25924 20544 25930 20556
rect 26345 20553 26357 20556
rect 26391 20553 26403 20587
rect 26510 20584 26516 20596
rect 26471 20556 26516 20584
rect 26345 20547 26403 20553
rect 26510 20544 26516 20556
rect 26568 20544 26574 20596
rect 13357 20519 13415 20525
rect 13357 20485 13369 20519
rect 13403 20485 13415 20519
rect 13538 20516 13544 20528
rect 13499 20488 13544 20516
rect 13357 20479 13415 20485
rect 13538 20476 13544 20488
rect 13596 20476 13602 20528
rect 14090 20525 14096 20528
rect 14084 20516 14096 20525
rect 14051 20488 14096 20516
rect 14084 20479 14096 20488
rect 14090 20476 14096 20479
rect 14148 20476 14154 20528
rect 18690 20516 18696 20528
rect 17328 20488 18696 20516
rect 9309 20451 9367 20457
rect 9309 20417 9321 20451
rect 9355 20448 9367 20451
rect 9674 20448 9680 20460
rect 9355 20420 9680 20448
rect 9355 20417 9367 20420
rect 9309 20411 9367 20417
rect 9674 20408 9680 20420
rect 9732 20408 9738 20460
rect 11790 20457 11796 20460
rect 11784 20411 11796 20457
rect 11848 20448 11854 20460
rect 13814 20448 13820 20460
rect 11848 20420 11884 20448
rect 13775 20420 13820 20448
rect 11790 20408 11796 20411
rect 11848 20408 11854 20420
rect 13814 20408 13820 20420
rect 13872 20408 13878 20460
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20448 15991 20451
rect 16390 20448 16396 20460
rect 15979 20420 16396 20448
rect 15979 20417 15991 20420
rect 15933 20411 15991 20417
rect 16390 20408 16396 20420
rect 16448 20408 16454 20460
rect 16942 20408 16948 20460
rect 17000 20448 17006 20460
rect 17328 20457 17356 20488
rect 18690 20476 18696 20488
rect 18748 20476 18754 20528
rect 19334 20476 19340 20528
rect 19392 20516 19398 20528
rect 19797 20519 19855 20525
rect 19797 20516 19809 20519
rect 19392 20488 19809 20516
rect 19392 20476 19398 20488
rect 19797 20485 19809 20488
rect 19843 20516 19855 20519
rect 20530 20516 20536 20528
rect 19843 20488 20536 20516
rect 19843 20485 19855 20488
rect 19797 20479 19855 20485
rect 20530 20476 20536 20488
rect 20588 20476 20594 20528
rect 25498 20516 25504 20528
rect 23400 20488 25504 20516
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 17000 20420 17325 20448
rect 17000 20408 17006 20420
rect 17313 20417 17325 20420
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20417 17463 20451
rect 18233 20451 18291 20457
rect 18233 20448 18245 20451
rect 17405 20411 17463 20417
rect 17788 20420 18245 20448
rect 8846 20340 8852 20392
rect 8904 20380 8910 20392
rect 9493 20383 9551 20389
rect 9493 20380 9505 20383
rect 8904 20352 9505 20380
rect 8904 20340 8910 20352
rect 9493 20349 9505 20352
rect 9539 20349 9551 20383
rect 11514 20380 11520 20392
rect 11475 20352 11520 20380
rect 9493 20343 9551 20349
rect 11514 20340 11520 20352
rect 11572 20340 11578 20392
rect 15749 20383 15807 20389
rect 15749 20349 15761 20383
rect 15795 20349 15807 20383
rect 15749 20343 15807 20349
rect 15841 20383 15899 20389
rect 15841 20349 15853 20383
rect 15887 20380 15899 20383
rect 16482 20380 16488 20392
rect 15887 20352 16488 20380
rect 15887 20349 15899 20352
rect 15841 20343 15899 20349
rect 15764 20312 15792 20343
rect 16482 20340 16488 20352
rect 16540 20340 16546 20392
rect 17129 20383 17187 20389
rect 17129 20349 17141 20383
rect 17175 20349 17187 20383
rect 17129 20343 17187 20349
rect 16206 20312 16212 20324
rect 15764 20284 16212 20312
rect 16206 20272 16212 20284
rect 16264 20312 16270 20324
rect 17144 20312 17172 20343
rect 17218 20340 17224 20392
rect 17276 20380 17282 20392
rect 17420 20380 17448 20411
rect 17276 20352 17448 20380
rect 17276 20340 17282 20352
rect 17788 20321 17816 20420
rect 18233 20417 18245 20420
rect 18279 20417 18291 20451
rect 18233 20411 18291 20417
rect 18322 20408 18328 20460
rect 18380 20448 18386 20460
rect 18380 20420 18425 20448
rect 18380 20408 18386 20420
rect 19058 20408 19064 20460
rect 19116 20448 19122 20460
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 19116 20420 19257 20448
rect 19116 20408 19122 20420
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 19613 20451 19671 20457
rect 19613 20417 19625 20451
rect 19659 20448 19671 20451
rect 20162 20448 20168 20460
rect 19659 20420 20168 20448
rect 19659 20417 19671 20420
rect 19613 20411 19671 20417
rect 20162 20408 20168 20420
rect 20220 20408 20226 20460
rect 20346 20457 20352 20460
rect 20340 20448 20352 20457
rect 20307 20420 20352 20448
rect 20340 20411 20352 20420
rect 20346 20408 20352 20411
rect 20404 20408 20410 20460
rect 23106 20448 23112 20460
rect 23067 20420 23112 20448
rect 23106 20408 23112 20420
rect 23164 20408 23170 20460
rect 23400 20457 23428 20488
rect 25498 20476 25504 20488
rect 25556 20476 25562 20528
rect 25682 20476 25688 20528
rect 25740 20516 25746 20528
rect 26145 20519 26203 20525
rect 26145 20516 26157 20519
rect 25740 20488 26157 20516
rect 25740 20476 25746 20488
rect 26145 20485 26157 20488
rect 26191 20485 26203 20519
rect 26145 20479 26203 20485
rect 23385 20451 23443 20457
rect 23385 20417 23397 20451
rect 23431 20448 23443 20451
rect 23474 20448 23480 20460
rect 23431 20420 23480 20448
rect 23431 20417 23443 20420
rect 23385 20411 23443 20417
rect 23474 20408 23480 20420
rect 23532 20408 23538 20460
rect 23842 20408 23848 20460
rect 23900 20448 23906 20460
rect 24581 20451 24639 20457
rect 24581 20448 24593 20451
rect 23900 20420 24593 20448
rect 23900 20408 23906 20420
rect 24581 20417 24593 20420
rect 24627 20417 24639 20451
rect 25314 20448 25320 20460
rect 25275 20420 25320 20448
rect 24581 20411 24639 20417
rect 25314 20408 25320 20420
rect 25372 20408 25378 20460
rect 25590 20448 25596 20460
rect 25551 20420 25596 20448
rect 25590 20408 25596 20420
rect 25648 20408 25654 20460
rect 26786 20408 26792 20460
rect 26844 20448 26850 20460
rect 27229 20451 27287 20457
rect 27229 20448 27241 20451
rect 26844 20420 27241 20448
rect 26844 20408 26850 20420
rect 27229 20417 27241 20420
rect 27275 20417 27287 20451
rect 27229 20411 27287 20417
rect 20073 20383 20131 20389
rect 20073 20349 20085 20383
rect 20119 20349 20131 20383
rect 20073 20343 20131 20349
rect 16264 20284 17172 20312
rect 17773 20315 17831 20321
rect 16264 20272 16270 20284
rect 17773 20281 17785 20315
rect 17819 20281 17831 20315
rect 17773 20275 17831 20281
rect 19242 20272 19248 20324
rect 19300 20312 19306 20324
rect 20088 20312 20116 20343
rect 21082 20340 21088 20392
rect 21140 20380 21146 20392
rect 23198 20380 23204 20392
rect 21140 20352 23204 20380
rect 21140 20340 21146 20352
rect 23198 20340 23204 20352
rect 23256 20380 23262 20392
rect 23661 20383 23719 20389
rect 23661 20380 23673 20383
rect 23256 20352 23673 20380
rect 23256 20340 23262 20352
rect 23661 20349 23673 20352
rect 23707 20349 23719 20383
rect 23661 20343 23719 20349
rect 24762 20340 24768 20392
rect 24820 20380 24826 20392
rect 24857 20383 24915 20389
rect 24857 20380 24869 20383
rect 24820 20352 24869 20380
rect 24820 20340 24826 20352
rect 24857 20349 24869 20352
rect 24903 20380 24915 20383
rect 25409 20383 25467 20389
rect 24903 20352 25176 20380
rect 24903 20349 24915 20352
rect 24857 20343 24915 20349
rect 19300 20284 20116 20312
rect 19300 20272 19306 20284
rect 21910 20272 21916 20324
rect 21968 20312 21974 20324
rect 24578 20312 24584 20324
rect 21968 20284 24584 20312
rect 21968 20272 21974 20284
rect 24578 20272 24584 20284
rect 24636 20272 24642 20324
rect 25148 20321 25176 20352
rect 25409 20349 25421 20383
rect 25455 20349 25467 20383
rect 25409 20343 25467 20349
rect 25133 20315 25191 20321
rect 25133 20281 25145 20315
rect 25179 20281 25191 20315
rect 25424 20312 25452 20343
rect 25498 20340 25504 20392
rect 25556 20380 25562 20392
rect 26050 20380 26056 20392
rect 25556 20352 26056 20380
rect 25556 20340 25562 20352
rect 26050 20340 26056 20352
rect 26108 20340 26114 20392
rect 26878 20340 26884 20392
rect 26936 20380 26942 20392
rect 26973 20383 27031 20389
rect 26973 20380 26985 20383
rect 26936 20352 26985 20380
rect 26936 20340 26942 20352
rect 26973 20349 26985 20352
rect 27019 20349 27031 20383
rect 26973 20343 27031 20349
rect 26418 20312 26424 20324
rect 25133 20275 25191 20281
rect 25240 20284 25452 20312
rect 25608 20284 26424 20312
rect 8386 20204 8392 20256
rect 8444 20244 8450 20256
rect 9125 20247 9183 20253
rect 9125 20244 9137 20247
rect 8444 20216 9137 20244
rect 8444 20204 8450 20216
rect 9125 20213 9137 20216
rect 9171 20213 9183 20247
rect 9125 20207 9183 20213
rect 12618 20204 12624 20256
rect 12676 20244 12682 20256
rect 13173 20247 13231 20253
rect 13173 20244 13185 20247
rect 12676 20216 13185 20244
rect 12676 20204 12682 20216
rect 13173 20213 13185 20216
rect 13219 20213 13231 20247
rect 15194 20244 15200 20256
rect 15155 20216 15200 20244
rect 13173 20207 13231 20213
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 16666 20244 16672 20256
rect 16627 20216 16672 20244
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 18414 20204 18420 20256
rect 18472 20244 18478 20256
rect 18693 20247 18751 20253
rect 18693 20244 18705 20247
rect 18472 20216 18705 20244
rect 18472 20204 18478 20216
rect 18693 20213 18705 20216
rect 18739 20213 18751 20247
rect 18693 20207 18751 20213
rect 18782 20204 18788 20256
rect 18840 20244 18846 20256
rect 19150 20244 19156 20256
rect 18840 20216 19156 20244
rect 18840 20204 18846 20216
rect 19150 20204 19156 20216
rect 19208 20204 19214 20256
rect 24026 20204 24032 20256
rect 24084 20244 24090 20256
rect 25240 20244 25268 20284
rect 25608 20253 25636 20284
rect 26418 20272 26424 20284
rect 26476 20272 26482 20324
rect 24084 20216 25268 20244
rect 25593 20247 25651 20253
rect 24084 20204 24090 20216
rect 25593 20213 25605 20247
rect 25639 20213 25651 20247
rect 26326 20244 26332 20256
rect 26287 20216 26332 20244
rect 25593 20207 25651 20213
rect 26326 20204 26332 20216
rect 26384 20204 26390 20256
rect 26436 20244 26464 20272
rect 28353 20247 28411 20253
rect 28353 20244 28365 20247
rect 26436 20216 28365 20244
rect 28353 20213 28365 20216
rect 28399 20213 28411 20247
rect 28353 20207 28411 20213
rect 1104 20154 28888 20176
rect 1104 20102 5582 20154
rect 5634 20102 5646 20154
rect 5698 20102 5710 20154
rect 5762 20102 5774 20154
rect 5826 20102 5838 20154
rect 5890 20102 14846 20154
rect 14898 20102 14910 20154
rect 14962 20102 14974 20154
rect 15026 20102 15038 20154
rect 15090 20102 15102 20154
rect 15154 20102 24110 20154
rect 24162 20102 24174 20154
rect 24226 20102 24238 20154
rect 24290 20102 24302 20154
rect 24354 20102 24366 20154
rect 24418 20102 28888 20154
rect 1104 20080 28888 20102
rect 11790 20040 11796 20052
rect 11751 20012 11796 20040
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 12250 20040 12256 20052
rect 12176 20012 12256 20040
rect 8386 19836 8392 19848
rect 8347 19808 8392 19836
rect 8386 19796 8392 19808
rect 8444 19796 8450 19848
rect 8938 19836 8944 19848
rect 8899 19808 8944 19836
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 12066 19845 12072 19848
rect 12049 19839 12072 19845
rect 12049 19805 12061 19839
rect 12049 19799 12072 19805
rect 12066 19796 12072 19799
rect 12124 19796 12130 19848
rect 12176 19842 12204 20012
rect 12250 20000 12256 20012
rect 12308 20000 12314 20052
rect 17126 20040 17132 20052
rect 15120 20012 17132 20040
rect 15120 19984 15148 20012
rect 17126 20000 17132 20012
rect 17184 20000 17190 20052
rect 17770 20040 17776 20052
rect 17731 20012 17776 20040
rect 17770 20000 17776 20012
rect 17828 20040 17834 20052
rect 20162 20040 20168 20052
rect 17828 20012 20168 20040
rect 17828 20000 17834 20012
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20346 20000 20352 20052
rect 20404 20040 20410 20052
rect 21082 20040 21088 20052
rect 20404 20012 21088 20040
rect 20404 20000 20410 20012
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 22925 20043 22983 20049
rect 22925 20009 22937 20043
rect 22971 20040 22983 20043
rect 23290 20040 23296 20052
rect 22971 20012 23296 20040
rect 22971 20009 22983 20012
rect 22925 20003 22983 20009
rect 23290 20000 23296 20012
rect 23348 20000 23354 20052
rect 23385 20043 23443 20049
rect 23385 20009 23397 20043
rect 23431 20040 23443 20043
rect 23842 20040 23848 20052
rect 23431 20012 23848 20040
rect 23431 20009 23443 20012
rect 23385 20003 23443 20009
rect 23842 20000 23848 20012
rect 23900 20000 23906 20052
rect 26786 20040 26792 20052
rect 26747 20012 26792 20040
rect 26786 20000 26792 20012
rect 26844 20000 26850 20052
rect 14274 19972 14280 19984
rect 13280 19944 14280 19972
rect 12618 19904 12624 19916
rect 12360 19876 12624 19904
rect 12174 19836 12232 19842
rect 12174 19802 12186 19836
rect 12220 19802 12232 19836
rect 12174 19796 12232 19802
rect 12274 19839 12332 19845
rect 12274 19805 12286 19839
rect 12320 19836 12332 19839
rect 12360 19836 12388 19876
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 13078 19904 13084 19916
rect 13039 19876 13084 19904
rect 13078 19864 13084 19876
rect 13136 19864 13142 19916
rect 12320 19808 12388 19836
rect 12437 19839 12495 19845
rect 12320 19805 12332 19808
rect 12274 19799 12332 19805
rect 12437 19805 12449 19839
rect 12483 19805 12495 19839
rect 12710 19836 12716 19848
rect 12671 19808 12716 19836
rect 12437 19799 12495 19805
rect 9186 19771 9244 19777
rect 9186 19768 9198 19771
rect 8588 19740 9198 19768
rect 8588 19709 8616 19740
rect 9186 19737 9198 19740
rect 9232 19737 9244 19771
rect 11333 19771 11391 19777
rect 11333 19768 11345 19771
rect 9186 19731 9244 19737
rect 9324 19740 11345 19768
rect 8573 19703 8631 19709
rect 8573 19669 8585 19703
rect 8619 19669 8631 19703
rect 8573 19663 8631 19669
rect 8846 19660 8852 19712
rect 8904 19700 8910 19712
rect 9324 19700 9352 19740
rect 11333 19737 11345 19740
rect 11379 19737 11391 19771
rect 11333 19731 11391 19737
rect 11517 19771 11575 19777
rect 11517 19737 11529 19771
rect 11563 19737 11575 19771
rect 11517 19731 11575 19737
rect 8904 19672 9352 19700
rect 8904 19660 8910 19672
rect 9858 19660 9864 19712
rect 9916 19700 9922 19712
rect 10321 19703 10379 19709
rect 10321 19700 10333 19703
rect 9916 19672 10333 19700
rect 9916 19660 9922 19672
rect 10321 19669 10333 19672
rect 10367 19669 10379 19703
rect 11532 19700 11560 19731
rect 12066 19700 12072 19712
rect 11532 19672 12072 19700
rect 10321 19663 10379 19669
rect 12066 19660 12072 19672
rect 12124 19700 12130 19712
rect 12452 19700 12480 19799
rect 12710 19796 12716 19808
rect 12768 19796 12774 19848
rect 13280 19845 13308 19944
rect 14274 19932 14280 19944
rect 14332 19972 14338 19984
rect 14918 19972 14924 19984
rect 14332 19944 14924 19972
rect 14332 19932 14338 19944
rect 14918 19932 14924 19944
rect 14976 19932 14982 19984
rect 15102 19932 15108 19984
rect 15160 19932 15166 19984
rect 15212 19944 15516 19972
rect 15212 19904 15240 19944
rect 14752 19876 15240 19904
rect 15488 19904 15516 19944
rect 23658 19932 23664 19984
rect 23716 19972 23722 19984
rect 25590 19972 25596 19984
rect 23716 19944 25596 19972
rect 23716 19932 23722 19944
rect 19242 19904 19248 19916
rect 15488 19876 15608 19904
rect 14752 19848 14780 19876
rect 13265 19839 13323 19845
rect 13265 19805 13277 19839
rect 13311 19805 13323 19839
rect 13265 19799 13323 19805
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19836 14703 19839
rect 14734 19836 14740 19848
rect 14691 19808 14740 19836
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 14918 19836 14924 19848
rect 14879 19808 14924 19836
rect 14918 19796 14924 19808
rect 14976 19796 14982 19848
rect 15102 19796 15108 19848
rect 15160 19836 15166 19848
rect 15580 19845 15608 19876
rect 17604 19876 19104 19904
rect 19203 19876 19248 19904
rect 15197 19839 15255 19845
rect 15197 19836 15209 19839
rect 15160 19808 15209 19836
rect 15160 19796 15166 19808
rect 15197 19805 15209 19808
rect 15243 19805 15255 19839
rect 15197 19799 15255 19805
rect 15381 19839 15439 19845
rect 15381 19805 15393 19839
rect 15427 19805 15439 19839
rect 15381 19799 15439 19805
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 15565 19839 15623 19845
rect 15565 19805 15577 19839
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 16393 19839 16451 19845
rect 16393 19805 16405 19839
rect 16439 19836 16451 19839
rect 17494 19836 17500 19848
rect 16439 19808 17500 19836
rect 16439 19805 16451 19808
rect 16393 19799 16451 19805
rect 14550 19728 14556 19780
rect 14608 19768 14614 19780
rect 15396 19768 15424 19799
rect 14608 19740 15424 19768
rect 15488 19768 15516 19799
rect 17494 19796 17500 19808
rect 17552 19796 17558 19848
rect 15654 19768 15660 19780
rect 15488 19740 15660 19768
rect 14608 19728 14614 19740
rect 15654 19728 15660 19740
rect 15712 19728 15718 19780
rect 15838 19768 15844 19780
rect 15799 19740 15844 19768
rect 15838 19728 15844 19740
rect 15896 19728 15902 19780
rect 16660 19771 16718 19777
rect 16660 19737 16672 19771
rect 16706 19768 16718 19771
rect 17034 19768 17040 19780
rect 16706 19740 17040 19768
rect 16706 19737 16718 19740
rect 16660 19731 16718 19737
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 12894 19700 12900 19712
rect 12124 19672 12900 19700
rect 12124 19660 12130 19672
rect 12894 19660 12900 19672
rect 12952 19660 12958 19712
rect 13449 19703 13507 19709
rect 13449 19669 13461 19703
rect 13495 19700 13507 19703
rect 13722 19700 13728 19712
rect 13495 19672 13728 19700
rect 13495 19669 13507 19672
rect 13449 19663 13507 19669
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 17604 19700 17632 19876
rect 18414 19836 18420 19848
rect 18375 19808 18420 19836
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 18509 19839 18567 19845
rect 18509 19805 18521 19839
rect 18555 19836 18567 19839
rect 18598 19836 18604 19848
rect 18555 19808 18604 19836
rect 18555 19805 18567 19808
rect 18509 19799 18567 19805
rect 18598 19796 18604 19808
rect 18656 19796 18662 19848
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 18966 19836 18972 19848
rect 18739 19808 18972 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 18966 19796 18972 19808
rect 19024 19796 19030 19848
rect 19076 19836 19104 19876
rect 19242 19864 19248 19876
rect 19300 19864 19306 19916
rect 21729 19907 21787 19913
rect 21729 19873 21741 19907
rect 21775 19904 21787 19907
rect 23201 19907 23259 19913
rect 23201 19904 23213 19907
rect 21775 19876 23213 19904
rect 21775 19873 21787 19876
rect 21729 19867 21787 19873
rect 23201 19873 23213 19876
rect 23247 19873 23259 19907
rect 24762 19904 24768 19916
rect 23201 19867 23259 19873
rect 23308 19876 24164 19904
rect 19886 19836 19892 19848
rect 19076 19808 19892 19836
rect 19886 19796 19892 19808
rect 19944 19796 19950 19848
rect 21450 19836 21456 19848
rect 21411 19808 21456 19836
rect 21450 19796 21456 19808
rect 21508 19796 21514 19848
rect 21542 19796 21548 19848
rect 21600 19836 21606 19848
rect 22189 19839 22247 19845
rect 21600 19808 21645 19836
rect 21600 19796 21606 19808
rect 22189 19805 22201 19839
rect 22235 19805 22247 19839
rect 22370 19836 22376 19848
rect 22331 19808 22376 19836
rect 22189 19799 22247 19805
rect 18877 19771 18935 19777
rect 18877 19737 18889 19771
rect 18923 19768 18935 19771
rect 19490 19771 19548 19777
rect 19490 19768 19502 19771
rect 18923 19740 19502 19768
rect 18923 19737 18935 19740
rect 18877 19731 18935 19737
rect 19490 19737 19502 19740
rect 19536 19737 19548 19771
rect 19490 19731 19548 19737
rect 22005 19771 22063 19777
rect 22005 19737 22017 19771
rect 22051 19737 22063 19771
rect 22204 19768 22232 19799
rect 22370 19796 22376 19808
rect 22428 19796 22434 19848
rect 22278 19768 22284 19780
rect 22191 19740 22284 19768
rect 22005 19731 22063 19737
rect 13872 19672 17632 19700
rect 18141 19703 18199 19709
rect 13872 19660 13878 19672
rect 18141 19669 18153 19703
rect 18187 19700 18199 19703
rect 18690 19700 18696 19712
rect 18187 19672 18696 19700
rect 18187 19669 18199 19672
rect 18141 19663 18199 19669
rect 18690 19660 18696 19672
rect 18748 19700 18754 19712
rect 19150 19700 19156 19712
rect 18748 19672 19156 19700
rect 18748 19660 18754 19672
rect 19150 19660 19156 19672
rect 19208 19660 19214 19712
rect 20622 19700 20628 19712
rect 20583 19672 20628 19700
rect 20622 19660 20628 19672
rect 20680 19660 20686 19712
rect 22020 19700 22048 19731
rect 22278 19728 22284 19740
rect 22336 19768 22342 19780
rect 23308 19768 23336 19876
rect 23474 19836 23480 19848
rect 23435 19808 23480 19836
rect 23474 19796 23480 19808
rect 23532 19796 23538 19848
rect 23658 19796 23664 19848
rect 23716 19836 23722 19848
rect 23845 19839 23903 19845
rect 23845 19836 23857 19839
rect 23716 19808 23857 19836
rect 23716 19796 23722 19808
rect 23845 19805 23857 19808
rect 23891 19805 23903 19839
rect 24026 19836 24032 19848
rect 23987 19808 24032 19836
rect 23845 19799 23903 19805
rect 24026 19796 24032 19808
rect 24084 19796 24090 19848
rect 22336 19740 23336 19768
rect 24136 19768 24164 19876
rect 24504 19876 24768 19904
rect 24504 19845 24532 19876
rect 24762 19864 24768 19876
rect 24820 19864 24826 19916
rect 24489 19839 24547 19845
rect 24489 19805 24501 19839
rect 24535 19805 24547 19839
rect 24670 19836 24676 19848
rect 24631 19808 24676 19836
rect 24489 19799 24547 19805
rect 24670 19796 24676 19808
rect 24728 19796 24734 19848
rect 24854 19836 24860 19848
rect 24815 19808 24860 19836
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 25332 19845 25360 19944
rect 25590 19932 25596 19944
rect 25648 19932 25654 19984
rect 26326 19904 26332 19916
rect 26068 19876 26332 19904
rect 25317 19839 25375 19845
rect 25317 19805 25329 19839
rect 25363 19805 25375 19839
rect 25317 19799 25375 19805
rect 25406 19796 25412 19848
rect 25464 19836 25470 19848
rect 26068 19845 26096 19876
rect 26326 19864 26332 19876
rect 26384 19864 26390 19916
rect 25777 19839 25835 19845
rect 25777 19836 25789 19839
rect 25464 19808 25789 19836
rect 25464 19796 25470 19808
rect 25777 19805 25789 19808
rect 25823 19805 25835 19839
rect 25777 19799 25835 19805
rect 26053 19839 26111 19845
rect 26053 19805 26065 19839
rect 26099 19805 26111 19839
rect 26053 19799 26111 19805
rect 26237 19839 26295 19845
rect 26237 19805 26249 19839
rect 26283 19836 26295 19839
rect 26513 19839 26571 19845
rect 26513 19836 26525 19839
rect 26283 19808 26525 19836
rect 26283 19805 26295 19808
rect 26237 19799 26295 19805
rect 26513 19805 26525 19808
rect 26559 19805 26571 19839
rect 26513 19799 26571 19805
rect 26602 19796 26608 19848
rect 26660 19796 26666 19848
rect 28350 19836 28356 19848
rect 28311 19808 28356 19836
rect 28350 19796 28356 19808
rect 28408 19796 28414 19848
rect 24136 19740 24532 19768
rect 22336 19728 22342 19740
rect 22186 19700 22192 19712
rect 22020 19672 22192 19700
rect 22186 19660 22192 19672
rect 22244 19660 22250 19712
rect 23934 19660 23940 19712
rect 23992 19700 23998 19712
rect 24504 19709 24532 19740
rect 26418 19728 26424 19780
rect 26476 19768 26482 19780
rect 26620 19768 26648 19796
rect 26789 19771 26847 19777
rect 26789 19768 26801 19771
rect 26476 19740 26801 19768
rect 26476 19728 26482 19740
rect 26789 19737 26801 19740
rect 26835 19737 26847 19771
rect 26789 19731 26847 19737
rect 24489 19703 24547 19709
rect 23992 19672 24037 19700
rect 23992 19660 23998 19672
rect 24489 19669 24501 19703
rect 24535 19669 24547 19703
rect 25406 19700 25412 19712
rect 25367 19672 25412 19700
rect 24489 19663 24547 19669
rect 25406 19660 25412 19672
rect 25464 19660 25470 19712
rect 25498 19660 25504 19712
rect 25556 19700 25562 19712
rect 25866 19700 25872 19712
rect 25556 19672 25872 19700
rect 25556 19660 25562 19672
rect 25866 19660 25872 19672
rect 25924 19660 25930 19712
rect 26234 19660 26240 19712
rect 26292 19700 26298 19712
rect 26605 19703 26663 19709
rect 26605 19700 26617 19703
rect 26292 19672 26617 19700
rect 26292 19660 26298 19672
rect 26605 19669 26617 19672
rect 26651 19669 26663 19703
rect 26605 19663 26663 19669
rect 1104 19610 28888 19632
rect 1104 19558 10214 19610
rect 10266 19558 10278 19610
rect 10330 19558 10342 19610
rect 10394 19558 10406 19610
rect 10458 19558 10470 19610
rect 10522 19558 19478 19610
rect 19530 19558 19542 19610
rect 19594 19558 19606 19610
rect 19658 19558 19670 19610
rect 19722 19558 19734 19610
rect 19786 19558 28888 19610
rect 1104 19536 28888 19558
rect 9674 19496 9680 19508
rect 9635 19468 9680 19496
rect 9674 19456 9680 19468
rect 9732 19456 9738 19508
rect 10045 19499 10103 19505
rect 10045 19465 10057 19499
rect 10091 19496 10103 19499
rect 10781 19499 10839 19505
rect 10781 19496 10793 19499
rect 10091 19468 10793 19496
rect 10091 19465 10103 19468
rect 10045 19459 10103 19465
rect 10781 19465 10793 19468
rect 10827 19496 10839 19499
rect 13814 19496 13820 19508
rect 10827 19468 13820 19496
rect 10827 19465 10839 19468
rect 10781 19459 10839 19465
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 14918 19456 14924 19508
rect 14976 19496 14982 19508
rect 15286 19496 15292 19508
rect 14976 19468 15292 19496
rect 14976 19456 14982 19468
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 15378 19456 15384 19508
rect 15436 19496 15442 19508
rect 15473 19499 15531 19505
rect 15473 19496 15485 19499
rect 15436 19468 15485 19496
rect 15436 19456 15442 19468
rect 15473 19465 15485 19468
rect 15519 19465 15531 19499
rect 15473 19459 15531 19465
rect 17494 19456 17500 19508
rect 17552 19496 17558 19508
rect 18141 19499 18199 19505
rect 18141 19496 18153 19499
rect 17552 19468 18153 19496
rect 17552 19456 17558 19468
rect 18141 19465 18153 19468
rect 18187 19496 18199 19499
rect 19242 19496 19248 19508
rect 18187 19468 19248 19496
rect 18187 19465 18199 19468
rect 18141 19459 18199 19465
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21361 19499 21419 19505
rect 21361 19496 21373 19499
rect 20864 19468 21373 19496
rect 20864 19456 20870 19468
rect 21361 19465 21373 19468
rect 21407 19465 21419 19499
rect 21361 19459 21419 19465
rect 23934 19456 23940 19508
rect 23992 19496 23998 19508
rect 25038 19496 25044 19508
rect 23992 19468 25044 19496
rect 23992 19456 23998 19468
rect 25038 19456 25044 19468
rect 25096 19496 25102 19508
rect 25409 19499 25467 19505
rect 25409 19496 25421 19499
rect 25096 19468 25421 19496
rect 25096 19456 25102 19468
rect 25409 19465 25421 19468
rect 25455 19496 25467 19499
rect 25498 19496 25504 19508
rect 25455 19468 25504 19496
rect 25455 19465 25467 19468
rect 25409 19459 25467 19465
rect 25498 19456 25504 19468
rect 25556 19456 25562 19508
rect 25593 19499 25651 19505
rect 25593 19465 25605 19499
rect 25639 19496 25651 19499
rect 26234 19496 26240 19508
rect 25639 19468 26240 19496
rect 25639 19465 25651 19468
rect 25593 19459 25651 19465
rect 26234 19456 26240 19468
rect 26292 19456 26298 19508
rect 27062 19496 27068 19508
rect 26528 19468 27068 19496
rect 11974 19428 11980 19440
rect 8496 19400 11980 19428
rect 8496 19372 8524 19400
rect 11974 19388 11980 19400
rect 12032 19388 12038 19440
rect 14369 19431 14427 19437
rect 14369 19428 14381 19431
rect 12084 19400 14381 19428
rect 8478 19360 8484 19372
rect 8439 19332 8484 19360
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 9030 19360 9036 19372
rect 8991 19332 9036 19360
rect 9030 19320 9036 19332
rect 9088 19320 9094 19372
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 10137 19363 10195 19369
rect 10137 19360 10149 19363
rect 9916 19332 10149 19360
rect 9916 19320 9922 19332
rect 10137 19329 10149 19332
rect 10183 19329 10195 19363
rect 10137 19323 10195 19329
rect 11330 19320 11336 19372
rect 11388 19360 11394 19372
rect 11517 19363 11575 19369
rect 11517 19360 11529 19363
rect 11388 19332 11529 19360
rect 11388 19320 11394 19332
rect 11517 19329 11529 19332
rect 11563 19360 11575 19363
rect 11701 19363 11759 19369
rect 11563 19332 11652 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 8021 19295 8079 19301
rect 8021 19261 8033 19295
rect 8067 19292 8079 19295
rect 8496 19292 8524 19320
rect 8846 19292 8852 19304
rect 8067 19264 8524 19292
rect 8807 19264 8852 19292
rect 8067 19261 8079 19264
rect 8021 19255 8079 19261
rect 8846 19252 8852 19264
rect 8904 19252 8910 19304
rect 10318 19292 10324 19304
rect 10279 19264 10324 19292
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 11624 19292 11652 19332
rect 11701 19329 11713 19363
rect 11747 19360 11759 19363
rect 11882 19360 11888 19372
rect 11747 19332 11888 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 11882 19320 11888 19332
rect 11940 19360 11946 19372
rect 12084 19360 12112 19400
rect 14369 19397 14381 19400
rect 14415 19397 14427 19431
rect 14369 19391 14427 19397
rect 14458 19388 14464 19440
rect 14516 19428 14522 19440
rect 16301 19431 16359 19437
rect 14516 19400 15148 19428
rect 14516 19388 14522 19400
rect 11940 19332 12112 19360
rect 12437 19363 12495 19369
rect 11940 19320 11946 19332
rect 12437 19329 12449 19363
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 12621 19363 12679 19369
rect 12621 19329 12633 19363
rect 12667 19360 12679 19363
rect 13630 19360 13636 19372
rect 12667 19332 13636 19360
rect 12667 19329 12679 19332
rect 12621 19323 12679 19329
rect 12452 19292 12480 19323
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 14182 19360 14188 19372
rect 14143 19332 14188 19360
rect 14182 19320 14188 19332
rect 14240 19320 14246 19372
rect 14829 19363 14887 19369
rect 14829 19360 14841 19363
rect 14476 19332 14841 19360
rect 11624 19264 12480 19292
rect 13909 19295 13967 19301
rect 13909 19261 13921 19295
rect 13955 19292 13967 19295
rect 14476 19292 14504 19332
rect 14829 19329 14841 19332
rect 14875 19360 14887 19363
rect 14918 19360 14924 19372
rect 14875 19332 14924 19360
rect 14875 19329 14887 19332
rect 14829 19323 14887 19329
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 15120 19369 15148 19400
rect 16301 19397 16313 19431
rect 16347 19428 16359 19431
rect 17218 19428 17224 19440
rect 16347 19400 17224 19428
rect 16347 19397 16359 19400
rect 16301 19391 16359 19397
rect 17218 19388 17224 19400
rect 17276 19388 17282 19440
rect 18233 19431 18291 19437
rect 18233 19397 18245 19431
rect 18279 19428 18291 19431
rect 19334 19428 19340 19440
rect 18279 19400 19340 19428
rect 18279 19397 18291 19400
rect 18233 19391 18291 19397
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 20162 19428 20168 19440
rect 20123 19400 20168 19428
rect 20162 19388 20168 19400
rect 20220 19388 20226 19440
rect 21913 19431 21971 19437
rect 20548 19400 21404 19428
rect 15013 19363 15071 19369
rect 15013 19329 15025 19363
rect 15059 19329 15071 19363
rect 15013 19323 15071 19329
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 15197 19363 15255 19369
rect 15197 19329 15209 19363
rect 15243 19329 15255 19363
rect 16114 19360 16120 19372
rect 16075 19332 16120 19360
rect 15197 19323 15255 19329
rect 13955 19264 14504 19292
rect 14553 19295 14611 19301
rect 13955 19261 13967 19264
rect 13909 19255 13967 19261
rect 14553 19261 14565 19295
rect 14599 19292 14611 19295
rect 15028 19292 15056 19323
rect 15212 19292 15240 19323
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19360 16727 19363
rect 17129 19363 17187 19369
rect 17129 19360 17141 19363
rect 16715 19332 17141 19360
rect 16715 19329 16727 19332
rect 16669 19323 16727 19329
rect 17129 19329 17141 19332
rect 17175 19329 17187 19363
rect 17310 19360 17316 19372
rect 17271 19332 17316 19360
rect 17129 19323 17187 19329
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 17862 19320 17868 19372
rect 17920 19360 17926 19372
rect 18598 19360 18604 19372
rect 17920 19332 18604 19360
rect 17920 19320 17926 19332
rect 18598 19320 18604 19332
rect 18656 19360 18662 19372
rect 18693 19363 18751 19369
rect 18693 19360 18705 19363
rect 18656 19332 18705 19360
rect 18656 19320 18662 19332
rect 18693 19329 18705 19332
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 18782 19320 18788 19372
rect 18840 19360 18846 19372
rect 18969 19363 19027 19369
rect 18840 19332 18885 19360
rect 18840 19320 18846 19332
rect 18969 19329 18981 19363
rect 19015 19360 19027 19363
rect 19150 19360 19156 19372
rect 19015 19332 19156 19360
rect 19015 19329 19027 19332
rect 18969 19323 19027 19329
rect 19150 19320 19156 19332
rect 19208 19320 19214 19372
rect 19518 19360 19524 19372
rect 19479 19332 19524 19360
rect 19518 19320 19524 19332
rect 19576 19320 19582 19372
rect 20548 19369 20576 19400
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 20625 19363 20683 19369
rect 20625 19329 20637 19363
rect 20671 19329 20683 19363
rect 20625 19323 20683 19329
rect 14599 19264 15056 19292
rect 15120 19264 15240 19292
rect 14599 19261 14611 19264
rect 14553 19255 14611 19261
rect 8294 19224 8300 19236
rect 8255 19196 8300 19224
rect 8294 19184 8300 19196
rect 8352 19184 8358 19236
rect 14734 19184 14740 19236
rect 14792 19224 14798 19236
rect 15120 19224 15148 19264
rect 15746 19252 15752 19304
rect 15804 19292 15810 19304
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15804 19264 15945 19292
rect 15804 19252 15810 19264
rect 15933 19261 15945 19264
rect 15979 19292 15991 19295
rect 17497 19295 17555 19301
rect 17497 19292 17509 19295
rect 15979 19264 17509 19292
rect 15979 19261 15991 19264
rect 15933 19255 15991 19261
rect 17497 19261 17509 19264
rect 17543 19292 17555 19295
rect 18322 19292 18328 19304
rect 17543 19264 18328 19292
rect 17543 19261 17555 19264
rect 17497 19255 17555 19261
rect 18322 19252 18328 19264
rect 18380 19252 18386 19304
rect 19978 19292 19984 19304
rect 18708 19264 19984 19292
rect 14792 19196 15148 19224
rect 14792 19184 14798 19196
rect 16298 19184 16304 19236
rect 16356 19224 16362 19236
rect 18708 19224 18736 19264
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 18966 19224 18972 19236
rect 16356 19196 18736 19224
rect 18927 19196 18972 19224
rect 16356 19184 16362 19196
rect 18966 19184 18972 19196
rect 19024 19184 19030 19236
rect 20640 19168 20668 19323
rect 20714 19320 20720 19372
rect 20772 19360 20778 19372
rect 20809 19363 20867 19369
rect 20809 19360 20821 19363
rect 20772 19332 20821 19360
rect 20772 19320 20778 19332
rect 20809 19329 20821 19332
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19360 21051 19363
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 21039 19332 21281 19360
rect 21039 19329 21051 19332
rect 20993 19323 21051 19329
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 21269 19323 21327 19329
rect 21376 19292 21404 19400
rect 21913 19397 21925 19431
rect 21959 19428 21971 19431
rect 21959 19400 24072 19428
rect 21959 19397 21971 19400
rect 21913 19391 21971 19397
rect 21450 19320 21456 19372
rect 21508 19360 21514 19372
rect 21818 19360 21824 19372
rect 21508 19332 21553 19360
rect 21779 19332 21824 19360
rect 21508 19320 21514 19332
rect 21818 19320 21824 19332
rect 21876 19320 21882 19372
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21928 19332 22017 19360
rect 21928 19292 21956 19332
rect 22005 19329 22017 19332
rect 22051 19360 22063 19363
rect 22051 19332 22232 19360
rect 22051 19329 22063 19332
rect 22005 19323 22063 19329
rect 21376 19264 21956 19292
rect 22204 19292 22232 19332
rect 22278 19320 22284 19372
rect 22336 19360 22342 19372
rect 22373 19363 22431 19369
rect 22373 19360 22385 19363
rect 22336 19332 22385 19360
rect 22336 19320 22342 19332
rect 22373 19329 22385 19332
rect 22419 19329 22431 19363
rect 22649 19363 22707 19369
rect 22649 19360 22661 19363
rect 22373 19323 22431 19329
rect 22480 19332 22661 19360
rect 22480 19292 22508 19332
rect 22649 19329 22661 19332
rect 22695 19360 22707 19363
rect 23658 19360 23664 19372
rect 22695 19332 23664 19360
rect 22695 19329 22707 19332
rect 22649 19323 22707 19329
rect 23658 19320 23664 19332
rect 23716 19320 23722 19372
rect 23934 19360 23940 19372
rect 23895 19332 23940 19360
rect 23934 19320 23940 19332
rect 23992 19320 23998 19372
rect 24044 19360 24072 19400
rect 24486 19388 24492 19440
rect 24544 19428 24550 19440
rect 24581 19431 24639 19437
rect 24581 19428 24593 19431
rect 24544 19400 24593 19428
rect 24544 19388 24550 19400
rect 24581 19397 24593 19400
rect 24627 19397 24639 19431
rect 24581 19391 24639 19397
rect 25130 19388 25136 19440
rect 25188 19428 25194 19440
rect 25317 19431 25375 19437
rect 25317 19428 25329 19431
rect 25188 19400 25329 19428
rect 25188 19388 25194 19400
rect 25317 19397 25329 19400
rect 25363 19397 25375 19431
rect 25317 19391 25375 19397
rect 26528 19372 26556 19468
rect 27062 19456 27068 19468
rect 27120 19456 27126 19508
rect 26605 19431 26663 19437
rect 26605 19397 26617 19431
rect 26651 19428 26663 19431
rect 27218 19431 27276 19437
rect 27218 19428 27230 19431
rect 26651 19400 27230 19428
rect 26651 19397 26663 19400
rect 26605 19391 26663 19397
rect 27218 19397 27230 19400
rect 27264 19397 27276 19431
rect 27218 19391 27276 19397
rect 25225 19363 25283 19369
rect 25225 19360 25237 19363
rect 24044 19332 25237 19360
rect 25225 19329 25237 19332
rect 25271 19329 25283 19363
rect 25225 19323 25283 19329
rect 25593 19363 25651 19369
rect 25593 19329 25605 19363
rect 25639 19360 25651 19363
rect 26326 19360 26332 19372
rect 25639 19332 26332 19360
rect 25639 19329 25651 19332
rect 25593 19323 25651 19329
rect 26326 19320 26332 19332
rect 26384 19320 26390 19372
rect 26421 19363 26479 19369
rect 26421 19329 26433 19363
rect 26467 19360 26479 19363
rect 26510 19360 26516 19372
rect 26467 19332 26516 19360
rect 26467 19329 26479 19332
rect 26421 19323 26479 19329
rect 26510 19320 26516 19332
rect 26568 19360 26574 19372
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 26568 19332 26661 19360
rect 26896 19332 26985 19360
rect 26568 19320 26574 19332
rect 22204 19264 22508 19292
rect 24213 19295 24271 19301
rect 24213 19261 24225 19295
rect 24259 19292 24271 19295
rect 24486 19292 24492 19304
rect 24259 19264 24492 19292
rect 24259 19261 24271 19264
rect 24213 19255 24271 19261
rect 24486 19252 24492 19264
rect 24544 19252 24550 19304
rect 25958 19252 25964 19304
rect 26016 19292 26022 19304
rect 26145 19295 26203 19301
rect 26145 19292 26157 19295
rect 26016 19264 26157 19292
rect 26016 19252 26022 19264
rect 26145 19261 26157 19264
rect 26191 19261 26203 19295
rect 26145 19255 26203 19261
rect 26896 19236 26924 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 22646 19184 22652 19236
rect 22704 19224 22710 19236
rect 24765 19227 24823 19233
rect 24765 19224 24777 19227
rect 22704 19196 24777 19224
rect 22704 19184 22710 19196
rect 24765 19193 24777 19196
rect 24811 19224 24823 19227
rect 26878 19224 26884 19236
rect 24811 19196 26884 19224
rect 24811 19193 24823 19196
rect 24765 19187 24823 19193
rect 26878 19184 26884 19196
rect 26936 19184 26942 19236
rect 9217 19159 9275 19165
rect 9217 19125 9229 19159
rect 9263 19156 9275 19159
rect 9490 19156 9496 19168
rect 9263 19128 9496 19156
rect 9263 19125 9275 19128
rect 9217 19119 9275 19125
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 11885 19159 11943 19165
rect 11885 19125 11897 19159
rect 11931 19156 11943 19159
rect 11974 19156 11980 19168
rect 11931 19128 11980 19156
rect 11931 19125 11943 19128
rect 11885 19119 11943 19125
rect 11974 19116 11980 19128
rect 12032 19116 12038 19168
rect 12618 19116 12624 19168
rect 12676 19156 12682 19168
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 12676 19128 12817 19156
rect 12676 19116 12682 19128
rect 12805 19125 12817 19128
rect 12851 19125 12863 19159
rect 12805 19119 12863 19125
rect 12894 19116 12900 19168
rect 12952 19156 12958 19168
rect 13173 19159 13231 19165
rect 13173 19156 13185 19159
rect 12952 19128 13185 19156
rect 12952 19116 12958 19128
rect 13173 19125 13185 19128
rect 13219 19125 13231 19159
rect 13173 19119 13231 19125
rect 16853 19159 16911 19165
rect 16853 19125 16865 19159
rect 16899 19156 16911 19159
rect 17586 19156 17592 19168
rect 16899 19128 17592 19156
rect 16899 19125 16911 19128
rect 16853 19119 16911 19125
rect 17586 19116 17592 19128
rect 17644 19116 17650 19168
rect 17678 19116 17684 19168
rect 17736 19156 17742 19168
rect 19613 19159 19671 19165
rect 19613 19156 19625 19159
rect 17736 19128 19625 19156
rect 17736 19116 17742 19128
rect 19613 19125 19625 19128
rect 19659 19125 19671 19159
rect 19613 19119 19671 19125
rect 20622 19116 20628 19168
rect 20680 19116 20686 19168
rect 23750 19156 23756 19168
rect 23711 19128 23756 19156
rect 23750 19116 23756 19128
rect 23808 19116 23814 19168
rect 24121 19159 24179 19165
rect 24121 19125 24133 19159
rect 24167 19156 24179 19159
rect 24578 19156 24584 19168
rect 24167 19128 24584 19156
rect 24167 19125 24179 19128
rect 24121 19119 24179 19125
rect 24578 19116 24584 19128
rect 24636 19116 24642 19168
rect 26234 19156 26240 19168
rect 26195 19128 26240 19156
rect 26234 19116 26240 19128
rect 26292 19116 26298 19168
rect 28166 19116 28172 19168
rect 28224 19156 28230 19168
rect 28353 19159 28411 19165
rect 28353 19156 28365 19159
rect 28224 19128 28365 19156
rect 28224 19116 28230 19128
rect 28353 19125 28365 19128
rect 28399 19125 28411 19159
rect 28353 19119 28411 19125
rect 1104 19066 28888 19088
rect 1104 19014 5582 19066
rect 5634 19014 5646 19066
rect 5698 19014 5710 19066
rect 5762 19014 5774 19066
rect 5826 19014 5838 19066
rect 5890 19014 14846 19066
rect 14898 19014 14910 19066
rect 14962 19014 14974 19066
rect 15026 19014 15038 19066
rect 15090 19014 15102 19066
rect 15154 19014 24110 19066
rect 24162 19014 24174 19066
rect 24226 19014 24238 19066
rect 24290 19014 24302 19066
rect 24354 19014 24366 19066
rect 24418 19014 28888 19066
rect 1104 18992 28888 19014
rect 9030 18912 9036 18964
rect 9088 18952 9094 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 9088 18924 9229 18952
rect 9088 18912 9094 18924
rect 9217 18921 9229 18924
rect 9263 18921 9275 18955
rect 11882 18952 11888 18964
rect 11843 18924 11888 18952
rect 9217 18915 9275 18921
rect 11882 18912 11888 18924
rect 11940 18912 11946 18964
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 13725 18955 13783 18961
rect 13725 18952 13737 18955
rect 13688 18924 13737 18952
rect 13688 18912 13694 18924
rect 13725 18921 13737 18924
rect 13771 18921 13783 18955
rect 14550 18952 14556 18964
rect 14511 18924 14556 18952
rect 13725 18915 13783 18921
rect 9030 18776 9036 18828
rect 9088 18816 9094 18828
rect 9769 18819 9827 18825
rect 9769 18816 9781 18819
rect 9088 18788 9781 18816
rect 9088 18776 9094 18788
rect 9769 18785 9781 18788
rect 9815 18816 9827 18819
rect 10318 18816 10324 18828
rect 9815 18788 10324 18816
rect 9815 18785 9827 18788
rect 9769 18779 9827 18785
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 11572 18788 12357 18816
rect 11572 18776 11578 18788
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 13740 18816 13768 18915
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 15746 18952 15752 18964
rect 15707 18924 15752 18952
rect 15746 18912 15752 18924
rect 15804 18912 15810 18964
rect 16025 18955 16083 18961
rect 16025 18921 16037 18955
rect 16071 18952 16083 18955
rect 16114 18952 16120 18964
rect 16071 18924 16120 18952
rect 16071 18921 16083 18924
rect 16025 18915 16083 18921
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 17034 18952 17040 18964
rect 16995 18924 17040 18952
rect 17034 18912 17040 18924
rect 17092 18912 17098 18964
rect 18877 18955 18935 18961
rect 18877 18921 18889 18955
rect 18923 18952 18935 18955
rect 19334 18952 19340 18964
rect 18923 18924 19340 18952
rect 18923 18921 18935 18924
rect 18877 18915 18935 18921
rect 19334 18912 19340 18924
rect 19392 18952 19398 18964
rect 19518 18952 19524 18964
rect 19392 18924 19524 18952
rect 19392 18912 19398 18924
rect 19518 18912 19524 18924
rect 19576 18912 19582 18964
rect 19613 18955 19671 18961
rect 19613 18921 19625 18955
rect 19659 18952 19671 18955
rect 20530 18952 20536 18964
rect 19659 18924 20536 18952
rect 19659 18921 19671 18924
rect 19613 18915 19671 18921
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 22189 18955 22247 18961
rect 22189 18921 22201 18955
rect 22235 18952 22247 18955
rect 22278 18952 22284 18964
rect 22235 18924 22284 18952
rect 22235 18921 22247 18924
rect 22189 18915 22247 18921
rect 22278 18912 22284 18924
rect 22336 18912 22342 18964
rect 22373 18955 22431 18961
rect 22373 18921 22385 18955
rect 22419 18952 22431 18955
rect 22554 18952 22560 18964
rect 22419 18924 22560 18952
rect 22419 18921 22431 18924
rect 22373 18915 22431 18921
rect 22554 18912 22560 18924
rect 22612 18912 22618 18964
rect 24026 18952 24032 18964
rect 23987 18924 24032 18952
rect 24026 18912 24032 18924
rect 24084 18912 24090 18964
rect 24397 18955 24455 18961
rect 24397 18921 24409 18955
rect 24443 18952 24455 18955
rect 24486 18952 24492 18964
rect 24443 18924 24492 18952
rect 24443 18921 24455 18924
rect 24397 18915 24455 18921
rect 24486 18912 24492 18924
rect 24544 18912 24550 18964
rect 25958 18952 25964 18964
rect 25919 18924 25964 18952
rect 25958 18912 25964 18924
rect 26016 18912 26022 18964
rect 26234 18952 26240 18964
rect 26195 18924 26240 18952
rect 26234 18912 26240 18924
rect 26292 18912 26298 18964
rect 27798 18952 27804 18964
rect 27759 18924 27804 18952
rect 27798 18912 27804 18924
rect 27856 18912 27862 18964
rect 28166 18952 28172 18964
rect 28127 18924 28172 18952
rect 28166 18912 28172 18924
rect 28224 18912 28230 18964
rect 13814 18844 13820 18896
rect 13872 18884 13878 18896
rect 13998 18884 14004 18896
rect 13872 18856 14004 18884
rect 13872 18844 13878 18856
rect 13998 18844 14004 18856
rect 14056 18884 14062 18896
rect 14056 18856 16712 18884
rect 14056 18844 14062 18856
rect 14829 18819 14887 18825
rect 14829 18816 14841 18819
rect 13740 18788 14841 18816
rect 12345 18779 12403 18785
rect 14829 18785 14841 18788
rect 14875 18785 14887 18819
rect 15194 18816 15200 18828
rect 14829 18779 14887 18785
rect 14936 18788 15200 18816
rect 7098 18748 7104 18760
rect 7059 18720 7104 18748
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 7561 18751 7619 18757
rect 7561 18717 7573 18751
rect 7607 18748 7619 18751
rect 8294 18748 8300 18760
rect 7607 18720 8300 18748
rect 7607 18717 7619 18720
rect 7561 18711 7619 18717
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 9585 18751 9643 18757
rect 9585 18717 9597 18751
rect 9631 18748 9643 18751
rect 9858 18748 9864 18760
rect 9631 18720 9864 18748
rect 9631 18717 9643 18720
rect 9585 18711 9643 18717
rect 9858 18708 9864 18720
rect 9916 18708 9922 18760
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18717 10563 18751
rect 10505 18711 10563 18717
rect 14369 18751 14427 18757
rect 14369 18717 14381 18751
rect 14415 18748 14427 18751
rect 14936 18748 14964 18788
rect 15194 18776 15200 18788
rect 15252 18776 15258 18828
rect 16206 18776 16212 18828
rect 16264 18816 16270 18828
rect 16574 18816 16580 18828
rect 16264 18788 16580 18816
rect 16264 18776 16270 18788
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 14415 18720 14964 18748
rect 15013 18751 15071 18757
rect 14415 18717 14427 18720
rect 14369 18711 14427 18717
rect 15013 18717 15025 18751
rect 15059 18717 15071 18751
rect 15013 18711 15071 18717
rect 15565 18751 15623 18757
rect 15565 18717 15577 18751
rect 15611 18748 15623 18751
rect 16114 18748 16120 18760
rect 15611 18720 16120 18748
rect 15611 18717 15623 18720
rect 15565 18711 15623 18717
rect 6638 18640 6644 18692
rect 6696 18680 6702 18692
rect 7377 18683 7435 18689
rect 7377 18680 7389 18683
rect 6696 18652 7389 18680
rect 6696 18640 6702 18652
rect 7377 18649 7389 18652
rect 7423 18680 7435 18683
rect 8938 18680 8944 18692
rect 7423 18652 8944 18680
rect 7423 18649 7435 18652
rect 7377 18643 7435 18649
rect 8938 18640 8944 18652
rect 8996 18680 9002 18692
rect 9398 18680 9404 18692
rect 8996 18652 9404 18680
rect 8996 18640 9002 18652
rect 9398 18640 9404 18652
rect 9456 18680 9462 18692
rect 10520 18680 10548 18711
rect 9456 18652 10548 18680
rect 10772 18683 10830 18689
rect 9456 18640 9462 18652
rect 10772 18649 10784 18683
rect 10818 18680 10830 18683
rect 11514 18680 11520 18692
rect 10818 18652 11520 18680
rect 10818 18649 10830 18652
rect 10772 18643 10830 18649
rect 11514 18640 11520 18652
rect 11572 18640 11578 18692
rect 12612 18683 12670 18689
rect 12612 18649 12624 18683
rect 12658 18680 12670 18683
rect 13078 18680 13084 18692
rect 12658 18652 13084 18680
rect 12658 18649 12670 18652
rect 12612 18643 12670 18649
rect 13078 18640 13084 18652
rect 13136 18640 13142 18692
rect 14182 18680 14188 18692
rect 14095 18652 14188 18680
rect 14182 18640 14188 18652
rect 14240 18640 14246 18692
rect 14274 18640 14280 18692
rect 14332 18680 14338 18692
rect 14734 18680 14740 18692
rect 14332 18652 14740 18680
rect 14332 18640 14338 18652
rect 14734 18640 14740 18652
rect 14792 18680 14798 18692
rect 15028 18680 15056 18711
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 14792 18652 15056 18680
rect 14792 18640 14798 18652
rect 15930 18640 15936 18692
rect 15988 18680 15994 18692
rect 16298 18680 16304 18692
rect 15988 18652 16304 18680
rect 15988 18640 15994 18652
rect 16298 18640 16304 18652
rect 16356 18680 16362 18692
rect 16485 18683 16543 18689
rect 16485 18680 16497 18683
rect 16356 18652 16497 18680
rect 16356 18640 16362 18652
rect 16485 18649 16497 18652
rect 16531 18649 16543 18683
rect 16684 18680 16712 18856
rect 19978 18844 19984 18896
rect 20036 18884 20042 18896
rect 20625 18887 20683 18893
rect 20625 18884 20637 18887
rect 20036 18856 20637 18884
rect 20036 18844 20042 18856
rect 20625 18853 20637 18856
rect 20671 18853 20683 18887
rect 22462 18884 22468 18896
rect 20625 18847 20683 18853
rect 21928 18856 22468 18884
rect 17494 18816 17500 18828
rect 17455 18788 17500 18816
rect 17494 18776 17500 18788
rect 17552 18776 17558 18828
rect 20162 18776 20168 18828
rect 20220 18816 20226 18828
rect 20533 18819 20591 18825
rect 20533 18816 20545 18819
rect 20220 18788 20545 18816
rect 20220 18776 20226 18788
rect 20533 18785 20545 18788
rect 20579 18785 20591 18819
rect 20640 18816 20668 18847
rect 20640 18788 20852 18816
rect 20533 18779 20591 18785
rect 17218 18748 17224 18760
rect 17179 18720 17224 18748
rect 17218 18708 17224 18720
rect 17276 18708 17282 18760
rect 17586 18708 17592 18760
rect 17644 18748 17650 18760
rect 17753 18751 17811 18757
rect 17753 18748 17765 18751
rect 17644 18720 17765 18748
rect 17644 18708 17650 18720
rect 17753 18717 17765 18720
rect 17799 18717 17811 18751
rect 19978 18748 19984 18760
rect 17753 18711 17811 18717
rect 17880 18720 19984 18748
rect 17880 18680 17908 18720
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 20438 18748 20444 18760
rect 20399 18720 20444 18748
rect 20438 18708 20444 18720
rect 20496 18708 20502 18760
rect 20714 18748 20720 18760
rect 20675 18720 20720 18748
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 16684 18652 17908 18680
rect 16485 18643 16543 18649
rect 19242 18640 19248 18692
rect 19300 18680 19306 18692
rect 19521 18683 19579 18689
rect 19521 18680 19533 18683
rect 19300 18652 19533 18680
rect 19300 18640 19306 18652
rect 19521 18649 19533 18652
rect 19567 18649 19579 18683
rect 20824 18680 20852 18788
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18748 20959 18751
rect 21821 18751 21879 18757
rect 21821 18748 21833 18751
rect 20947 18720 21833 18748
rect 20947 18717 20959 18720
rect 20901 18711 20959 18717
rect 21821 18717 21833 18720
rect 21867 18748 21879 18751
rect 21928 18748 21956 18856
rect 22462 18844 22468 18856
rect 22520 18844 22526 18896
rect 24670 18884 24676 18896
rect 24642 18844 24676 18884
rect 24728 18844 24734 18896
rect 26881 18887 26939 18893
rect 26881 18884 26893 18887
rect 26436 18856 26893 18884
rect 22094 18816 22100 18828
rect 21867 18720 21956 18748
rect 22020 18788 22100 18816
rect 21867 18717 21879 18720
rect 21821 18711 21879 18717
rect 22020 18680 22048 18788
rect 22094 18776 22100 18788
rect 22152 18776 22158 18828
rect 22646 18816 22652 18828
rect 22607 18788 22652 18816
rect 22646 18776 22652 18788
rect 22704 18776 22710 18828
rect 22916 18751 22974 18757
rect 22916 18717 22928 18751
rect 22962 18748 22974 18751
rect 23750 18748 23756 18760
rect 22962 18720 23756 18748
rect 22962 18717 22974 18720
rect 22916 18711 22974 18717
rect 23750 18708 23756 18720
rect 23808 18708 23814 18760
rect 24642 18757 24670 18844
rect 25498 18776 25504 18828
rect 25556 18816 25562 18828
rect 26436 18816 26464 18856
rect 26881 18853 26893 18856
rect 26927 18884 26939 18887
rect 27062 18884 27068 18896
rect 26927 18856 27068 18884
rect 26927 18853 26939 18856
rect 26881 18847 26939 18853
rect 27062 18844 27068 18856
rect 27120 18844 27126 18896
rect 27433 18819 27491 18825
rect 27433 18816 27445 18819
rect 25556 18788 26464 18816
rect 26528 18788 27445 18816
rect 25556 18776 25562 18788
rect 24642 18751 24711 18757
rect 24878 18751 24936 18757
rect 24642 18720 24665 18751
rect 24653 18717 24665 18720
rect 24699 18717 24711 18751
rect 24653 18711 24711 18717
rect 24778 18745 24836 18751
rect 24878 18748 24890 18751
rect 24778 18711 24790 18745
rect 24824 18711 24836 18745
rect 24778 18705 24836 18711
rect 24872 18717 24890 18748
rect 24924 18717 24936 18751
rect 25038 18748 25044 18760
rect 24999 18720 25044 18748
rect 24872 18711 24936 18717
rect 20824 18652 22048 18680
rect 19521 18643 19579 18649
rect 6914 18612 6920 18624
rect 6875 18584 6920 18612
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 9677 18615 9735 18621
rect 9677 18581 9689 18615
rect 9723 18612 9735 18615
rect 9950 18612 9956 18624
rect 9723 18584 9956 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 14200 18612 14228 18640
rect 14366 18612 14372 18624
rect 14200 18584 14372 18612
rect 14366 18572 14372 18584
rect 14424 18572 14430 18624
rect 15194 18612 15200 18624
rect 15155 18584 15200 18612
rect 15194 18572 15200 18584
rect 15252 18572 15258 18624
rect 16390 18612 16396 18624
rect 16351 18584 16396 18612
rect 16390 18572 16396 18584
rect 16448 18612 16454 18624
rect 16666 18612 16672 18624
rect 16448 18584 16672 18612
rect 16448 18572 16454 18584
rect 16666 18572 16672 18584
rect 16724 18572 16730 18624
rect 21358 18572 21364 18624
rect 21416 18612 21422 18624
rect 22189 18615 22247 18621
rect 22189 18612 22201 18615
rect 21416 18584 22201 18612
rect 21416 18572 21422 18584
rect 22189 18581 22201 18584
rect 22235 18581 22247 18615
rect 22189 18575 22247 18581
rect 22370 18572 22376 18624
rect 22428 18612 22434 18624
rect 24780 18612 24808 18705
rect 24872 18680 24900 18711
rect 25038 18708 25044 18720
rect 25096 18708 25102 18760
rect 25685 18751 25743 18757
rect 25685 18717 25697 18751
rect 25731 18748 25743 18751
rect 25866 18748 25872 18760
rect 25731 18720 25872 18748
rect 25731 18717 25743 18720
rect 25685 18711 25743 18717
rect 25866 18708 25872 18720
rect 25924 18708 25930 18760
rect 25961 18751 26019 18757
rect 25961 18717 25973 18751
rect 26007 18748 26019 18751
rect 26326 18748 26332 18760
rect 26007 18720 26332 18748
rect 26007 18717 26019 18720
rect 25961 18711 26019 18717
rect 26326 18708 26332 18720
rect 26384 18748 26390 18760
rect 26528 18757 26556 18788
rect 27433 18785 27445 18788
rect 27479 18785 27491 18819
rect 28184 18816 28212 18912
rect 27433 18779 27491 18785
rect 27540 18788 28212 18816
rect 27540 18757 27568 18788
rect 26513 18751 26571 18757
rect 26513 18748 26525 18751
rect 26384 18720 26525 18748
rect 26384 18708 26390 18720
rect 26513 18717 26525 18720
rect 26559 18717 26571 18751
rect 26513 18711 26571 18717
rect 26973 18751 27031 18757
rect 26973 18717 26985 18751
rect 27019 18717 27031 18751
rect 26973 18711 27031 18717
rect 27525 18751 27583 18757
rect 27525 18717 27537 18751
rect 27571 18717 27583 18751
rect 28074 18748 28080 18760
rect 28035 18720 28080 18748
rect 27525 18711 27583 18717
rect 25130 18680 25136 18692
rect 24872 18652 25136 18680
rect 25130 18640 25136 18652
rect 25188 18680 25194 18692
rect 26697 18683 26755 18689
rect 26697 18680 26709 18683
rect 25188 18652 26709 18680
rect 25188 18640 25194 18652
rect 26697 18649 26709 18652
rect 26743 18649 26755 18683
rect 26988 18680 27016 18711
rect 28074 18708 28080 18720
rect 28132 18708 28138 18760
rect 28169 18751 28227 18757
rect 28169 18717 28181 18751
rect 28215 18748 28227 18751
rect 28258 18748 28264 18760
rect 28215 18720 28264 18748
rect 28215 18717 28227 18720
rect 28169 18711 28227 18717
rect 28258 18708 28264 18720
rect 28316 18708 28322 18760
rect 28092 18680 28120 18708
rect 26988 18652 28120 18680
rect 26697 18643 26755 18649
rect 22428 18584 24808 18612
rect 25777 18615 25835 18621
rect 22428 18572 22434 18584
rect 25777 18581 25789 18615
rect 25823 18612 25835 18615
rect 26418 18612 26424 18624
rect 25823 18584 26424 18612
rect 25823 18581 25835 18584
rect 25777 18575 25835 18581
rect 26418 18572 26424 18584
rect 26476 18612 26482 18624
rect 26605 18615 26663 18621
rect 26605 18612 26617 18615
rect 26476 18584 26617 18612
rect 26476 18572 26482 18584
rect 26605 18581 26617 18584
rect 26651 18581 26663 18615
rect 26605 18575 26663 18581
rect 1104 18522 28888 18544
rect 1104 18470 10214 18522
rect 10266 18470 10278 18522
rect 10330 18470 10342 18522
rect 10394 18470 10406 18522
rect 10458 18470 10470 18522
rect 10522 18470 19478 18522
rect 19530 18470 19542 18522
rect 19594 18470 19606 18522
rect 19658 18470 19670 18522
rect 19722 18470 19734 18522
rect 19786 18470 28888 18522
rect 1104 18448 28888 18470
rect 7374 18368 7380 18420
rect 7432 18408 7438 18420
rect 8021 18411 8079 18417
rect 8021 18408 8033 18411
rect 7432 18380 8033 18408
rect 7432 18368 7438 18380
rect 8021 18377 8033 18380
rect 8067 18408 8079 18411
rect 8757 18411 8815 18417
rect 8757 18408 8769 18411
rect 8067 18380 8769 18408
rect 8067 18377 8079 18380
rect 8021 18371 8079 18377
rect 8757 18377 8769 18380
rect 8803 18377 8815 18411
rect 11514 18408 11520 18420
rect 11475 18380 11520 18408
rect 8757 18371 8815 18377
rect 11514 18368 11520 18380
rect 11572 18368 11578 18420
rect 13078 18408 13084 18420
rect 13039 18380 13084 18408
rect 13078 18368 13084 18380
rect 13136 18368 13142 18420
rect 15378 18408 15384 18420
rect 14384 18380 15384 18408
rect 6914 18349 6920 18352
rect 6908 18340 6920 18349
rect 6875 18312 6920 18340
rect 6908 18303 6920 18312
rect 6914 18300 6920 18303
rect 6972 18300 6978 18352
rect 13814 18340 13820 18352
rect 7576 18312 11652 18340
rect 2521 18275 2579 18281
rect 2521 18241 2533 18275
rect 2567 18272 2579 18275
rect 7576 18272 7604 18312
rect 2567 18244 7604 18272
rect 8665 18275 8723 18281
rect 2567 18241 2579 18244
rect 2521 18235 2579 18241
rect 8665 18241 8677 18275
rect 8711 18272 8723 18275
rect 9490 18272 9496 18284
rect 8711 18244 9352 18272
rect 9451 18244 9496 18272
rect 8711 18241 8723 18244
rect 8665 18235 8723 18241
rect 2777 18207 2835 18213
rect 2777 18173 2789 18207
rect 2823 18204 2835 18207
rect 5166 18204 5172 18216
rect 2823 18176 5172 18204
rect 2823 18173 2835 18176
rect 2777 18167 2835 18173
rect 5166 18164 5172 18176
rect 5224 18204 5230 18216
rect 6638 18204 6644 18216
rect 5224 18176 6644 18204
rect 5224 18164 5230 18176
rect 6638 18164 6644 18176
rect 6696 18164 6702 18216
rect 8941 18207 8999 18213
rect 8941 18173 8953 18207
rect 8987 18204 8999 18207
rect 9030 18204 9036 18216
rect 8987 18176 9036 18204
rect 8987 18173 8999 18176
rect 8941 18167 8999 18173
rect 9030 18164 9036 18176
rect 9088 18164 9094 18216
rect 9324 18136 9352 18244
rect 9490 18232 9496 18244
rect 9548 18232 9554 18284
rect 10036 18275 10094 18281
rect 10036 18241 10048 18275
rect 10082 18272 10094 18275
rect 11514 18272 11520 18284
rect 10082 18244 11520 18272
rect 10082 18241 10094 18244
rect 10036 18235 10094 18241
rect 11514 18232 11520 18244
rect 11572 18232 11578 18284
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 9769 18207 9827 18213
rect 9769 18204 9781 18207
rect 9456 18176 9781 18204
rect 9456 18164 9462 18176
rect 9769 18173 9781 18176
rect 9815 18173 9827 18207
rect 9769 18167 9827 18173
rect 11624 18136 11652 18312
rect 13556 18312 13820 18340
rect 11698 18232 11704 18284
rect 11756 18281 11762 18284
rect 11756 18275 11805 18281
rect 11756 18241 11759 18275
rect 11793 18241 11805 18275
rect 11756 18235 11805 18241
rect 11882 18275 11940 18281
rect 11882 18241 11894 18275
rect 11928 18241 11940 18275
rect 11882 18235 11940 18241
rect 11756 18232 11762 18235
rect 11900 18204 11928 18235
rect 11974 18232 11980 18284
rect 12032 18281 12038 18284
rect 12032 18272 12040 18281
rect 12158 18272 12164 18284
rect 12032 18244 12077 18272
rect 12119 18244 12164 18272
rect 12032 18235 12040 18244
rect 12032 18232 12038 18235
rect 12158 18232 12164 18244
rect 12216 18272 12222 18284
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 12216 18244 12449 18272
rect 12216 18232 12222 18244
rect 12437 18241 12449 18244
rect 12483 18241 12495 18275
rect 12618 18272 12624 18284
rect 12579 18244 12624 18272
rect 12437 18235 12495 18241
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 12716 18275 12774 18281
rect 12716 18241 12728 18275
rect 12762 18241 12774 18275
rect 12716 18235 12774 18241
rect 12825 18275 12883 18281
rect 12825 18241 12837 18275
rect 12871 18272 12883 18275
rect 12986 18272 12992 18284
rect 12871 18244 12992 18272
rect 12871 18241 12883 18244
rect 12825 18235 12883 18241
rect 12342 18204 12348 18216
rect 11900 18176 12348 18204
rect 12342 18164 12348 18176
rect 12400 18204 12406 18216
rect 12731 18204 12759 18235
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 13556 18281 13584 18312
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18241 13599 18275
rect 13722 18272 13728 18284
rect 13683 18244 13728 18272
rect 13541 18235 13599 18241
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 14384 18281 14412 18380
rect 15378 18368 15384 18380
rect 15436 18368 15442 18420
rect 15562 18368 15568 18420
rect 15620 18408 15626 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 15620 18380 15669 18408
rect 15620 18368 15626 18380
rect 15657 18377 15669 18380
rect 15703 18377 15715 18411
rect 15657 18371 15715 18377
rect 16114 18368 16120 18420
rect 16172 18368 16178 18420
rect 16850 18408 16856 18420
rect 16811 18380 16856 18408
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 17221 18411 17279 18417
rect 17221 18377 17233 18411
rect 17267 18408 17279 18411
rect 17310 18408 17316 18420
rect 17267 18380 17316 18408
rect 17267 18377 17279 18380
rect 17221 18371 17279 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 17402 18368 17408 18420
rect 17460 18408 17466 18420
rect 17678 18408 17684 18420
rect 17460 18380 17684 18408
rect 17460 18368 17466 18380
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 19076 18380 21036 18408
rect 16022 18340 16028 18352
rect 14476 18312 16028 18340
rect 14476 18281 14504 18312
rect 14369 18275 14427 18281
rect 14369 18241 14381 18275
rect 14415 18241 14427 18275
rect 14369 18235 14427 18241
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 14734 18272 14740 18284
rect 14608 18244 14653 18272
rect 14695 18244 14740 18272
rect 14608 18232 14614 18244
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 15304 18281 15332 18312
rect 16022 18300 16028 18312
rect 16080 18300 16086 18352
rect 16132 18340 16160 18368
rect 16761 18343 16819 18349
rect 16761 18340 16773 18343
rect 16132 18312 16773 18340
rect 16761 18309 16773 18312
rect 16807 18309 16819 18343
rect 16868 18340 16896 18368
rect 19076 18340 19104 18380
rect 19242 18340 19248 18352
rect 16868 18312 19104 18340
rect 19203 18312 19248 18340
rect 16761 18303 16819 18309
rect 19242 18300 19248 18312
rect 19300 18300 19306 18352
rect 19352 18312 20944 18340
rect 15013 18275 15071 18281
rect 15013 18241 15025 18275
rect 15059 18241 15071 18275
rect 15013 18235 15071 18241
rect 15197 18275 15255 18281
rect 15197 18241 15209 18275
rect 15243 18241 15255 18275
rect 15197 18235 15255 18241
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18241 15347 18275
rect 15289 18235 15347 18241
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 12400 18176 12759 18204
rect 13817 18207 13875 18213
rect 12400 18164 12406 18176
rect 13817 18173 13829 18207
rect 13863 18204 13875 18207
rect 14093 18207 14151 18213
rect 14093 18204 14105 18207
rect 13863 18176 14105 18204
rect 13863 18173 13875 18176
rect 13817 18167 13875 18173
rect 14093 18173 14105 18176
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 13357 18139 13415 18145
rect 13357 18136 13369 18139
rect 9324 18108 9444 18136
rect 11624 18108 13369 18136
rect 1397 18071 1455 18077
rect 1397 18037 1409 18071
rect 1443 18068 1455 18071
rect 1670 18068 1676 18080
rect 1443 18040 1676 18068
rect 1443 18037 1455 18040
rect 1397 18031 1455 18037
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 8297 18071 8355 18077
rect 8297 18037 8309 18071
rect 8343 18068 8355 18071
rect 8386 18068 8392 18080
rect 8343 18040 8392 18068
rect 8343 18037 8355 18040
rect 8297 18031 8355 18037
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 9214 18028 9220 18080
rect 9272 18068 9278 18080
rect 9309 18071 9367 18077
rect 9309 18068 9321 18071
rect 9272 18040 9321 18068
rect 9272 18028 9278 18040
rect 9309 18037 9321 18040
rect 9355 18037 9367 18071
rect 9416 18068 9444 18108
rect 13357 18105 13369 18108
rect 13403 18105 13415 18139
rect 13357 18099 13415 18105
rect 13538 18096 13544 18148
rect 13596 18136 13602 18148
rect 15028 18136 15056 18235
rect 13596 18108 15056 18136
rect 13596 18096 13602 18108
rect 9950 18068 9956 18080
rect 9416 18040 9956 18068
rect 9309 18031 9367 18037
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11149 18071 11207 18077
rect 11149 18068 11161 18071
rect 11112 18040 11161 18068
rect 11112 18028 11118 18040
rect 11149 18037 11161 18040
rect 11195 18037 11207 18071
rect 11149 18031 11207 18037
rect 11882 18028 11888 18080
rect 11940 18068 11946 18080
rect 12158 18068 12164 18080
rect 11940 18040 12164 18068
rect 11940 18028 11946 18040
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 14366 18028 14372 18080
rect 14424 18068 14430 18080
rect 15212 18068 15240 18235
rect 15396 18204 15424 18235
rect 15746 18232 15752 18284
rect 15804 18272 15810 18284
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15804 18244 15945 18272
rect 15804 18232 15810 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18272 16175 18275
rect 16666 18272 16672 18284
rect 16163 18244 16672 18272
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 16666 18232 16672 18244
rect 16724 18232 16730 18284
rect 17586 18272 17592 18284
rect 17547 18244 17592 18272
rect 17586 18232 17592 18244
rect 17644 18272 17650 18284
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 17644 18244 18613 18272
rect 17644 18232 17650 18244
rect 18601 18241 18613 18244
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 18874 18232 18880 18284
rect 18932 18272 18938 18284
rect 19352 18272 19380 18312
rect 18932 18244 19380 18272
rect 19521 18275 19579 18281
rect 18932 18232 18938 18244
rect 19521 18241 19533 18275
rect 19567 18272 19579 18275
rect 19886 18272 19892 18284
rect 19567 18244 19892 18272
rect 19567 18241 19579 18244
rect 19521 18235 19579 18241
rect 19886 18232 19892 18244
rect 19944 18232 19950 18284
rect 20162 18272 20168 18284
rect 20123 18244 20168 18272
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20438 18272 20444 18284
rect 20399 18244 20444 18272
rect 20438 18232 20444 18244
rect 20496 18232 20502 18284
rect 16942 18204 16948 18216
rect 15396 18176 16948 18204
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 17862 18204 17868 18216
rect 17823 18176 17868 18204
rect 17862 18164 17868 18176
rect 17920 18164 17926 18216
rect 18506 18164 18512 18216
rect 18564 18204 18570 18216
rect 19337 18207 19395 18213
rect 19337 18204 19349 18207
rect 18564 18176 19349 18204
rect 18564 18164 18570 18176
rect 19337 18173 19349 18176
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 15378 18096 15384 18148
rect 15436 18136 15442 18148
rect 19058 18136 19064 18148
rect 15436 18108 19064 18136
rect 15436 18096 15442 18108
rect 19058 18096 19064 18108
rect 19116 18136 19122 18148
rect 19705 18139 19763 18145
rect 19116 18108 19472 18136
rect 19116 18096 19122 18108
rect 14424 18040 15240 18068
rect 16301 18071 16359 18077
rect 14424 18028 14430 18040
rect 16301 18037 16313 18071
rect 16347 18068 16359 18071
rect 16758 18068 16764 18080
rect 16347 18040 16764 18068
rect 16347 18037 16359 18040
rect 16301 18031 16359 18037
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 17126 18028 17132 18080
rect 17184 18068 17190 18080
rect 18230 18068 18236 18080
rect 17184 18040 18236 18068
rect 17184 18028 17190 18040
rect 18230 18028 18236 18040
rect 18288 18068 18294 18080
rect 18874 18068 18880 18080
rect 18288 18040 18880 18068
rect 18288 18028 18294 18040
rect 18874 18028 18880 18040
rect 18932 18028 18938 18080
rect 19334 18068 19340 18080
rect 19295 18040 19340 18068
rect 19334 18028 19340 18040
rect 19392 18028 19398 18080
rect 19444 18068 19472 18108
rect 19705 18105 19717 18139
rect 19751 18136 19763 18139
rect 20180 18136 20208 18232
rect 20254 18164 20260 18216
rect 20312 18204 20318 18216
rect 20916 18204 20944 18312
rect 21008 18281 21036 18380
rect 21634 18368 21640 18420
rect 21692 18408 21698 18420
rect 22922 18408 22928 18420
rect 21692 18380 22928 18408
rect 21692 18368 21698 18380
rect 22922 18368 22928 18380
rect 22980 18368 22986 18420
rect 24578 18408 24584 18420
rect 24539 18380 24584 18408
rect 24578 18368 24584 18380
rect 24636 18368 24642 18420
rect 24673 18411 24731 18417
rect 24673 18377 24685 18411
rect 24719 18408 24731 18411
rect 25406 18408 25412 18420
rect 24719 18380 25412 18408
rect 24719 18377 24731 18380
rect 24673 18371 24731 18377
rect 25406 18368 25412 18380
rect 25464 18368 25470 18420
rect 27338 18340 27344 18352
rect 21100 18312 27344 18340
rect 20993 18275 21051 18281
rect 20993 18241 21005 18275
rect 21039 18241 21051 18275
rect 20993 18235 21051 18241
rect 21100 18204 21128 18312
rect 27338 18300 27344 18312
rect 27396 18300 27402 18352
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 22152 18244 22197 18272
rect 22152 18232 22158 18244
rect 22922 18232 22928 18284
rect 22980 18272 22986 18284
rect 23477 18275 23535 18281
rect 23477 18272 23489 18275
rect 22980 18244 23489 18272
rect 22980 18232 22986 18244
rect 23477 18241 23489 18244
rect 23523 18241 23535 18275
rect 23477 18235 23535 18241
rect 24026 18232 24032 18284
rect 24084 18272 24090 18284
rect 24305 18275 24363 18281
rect 24305 18272 24317 18275
rect 24084 18244 24317 18272
rect 24084 18232 24090 18244
rect 24305 18241 24317 18244
rect 24351 18241 24363 18275
rect 24305 18235 24363 18241
rect 24765 18275 24823 18281
rect 24765 18241 24777 18275
rect 24811 18272 24823 18275
rect 25866 18272 25872 18284
rect 24811 18244 25872 18272
rect 24811 18241 24823 18244
rect 24765 18235 24823 18241
rect 25866 18232 25872 18244
rect 25924 18232 25930 18284
rect 26050 18232 26056 18284
rect 26108 18272 26114 18284
rect 26145 18275 26203 18281
rect 26145 18272 26157 18275
rect 26108 18244 26157 18272
rect 26108 18232 26114 18244
rect 26145 18241 26157 18244
rect 26191 18241 26203 18275
rect 26326 18272 26332 18284
rect 26287 18244 26332 18272
rect 26145 18235 26203 18241
rect 26326 18232 26332 18244
rect 26384 18232 26390 18284
rect 27157 18275 27215 18281
rect 27157 18241 27169 18275
rect 27203 18272 27215 18275
rect 28074 18272 28080 18284
rect 27203 18244 28080 18272
rect 27203 18241 27215 18244
rect 27157 18235 27215 18241
rect 28074 18232 28080 18244
rect 28132 18232 28138 18284
rect 28353 18275 28411 18281
rect 28353 18241 28365 18275
rect 28399 18272 28411 18275
rect 28442 18272 28448 18284
rect 28399 18244 28448 18272
rect 28399 18241 28411 18244
rect 28353 18235 28411 18241
rect 28442 18232 28448 18244
rect 28500 18232 28506 18284
rect 20312 18176 20357 18204
rect 20916 18176 21128 18204
rect 20312 18164 20318 18176
rect 21174 18164 21180 18216
rect 21232 18204 21238 18216
rect 22002 18204 22008 18216
rect 21232 18176 21496 18204
rect 21963 18176 22008 18204
rect 21232 18164 21238 18176
rect 19751 18108 20208 18136
rect 20625 18139 20683 18145
rect 19751 18105 19763 18108
rect 19705 18099 19763 18105
rect 20625 18105 20637 18139
rect 20671 18136 20683 18139
rect 21358 18136 21364 18148
rect 20671 18108 21364 18136
rect 20671 18105 20683 18108
rect 20625 18099 20683 18105
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 21468 18136 21496 18176
rect 22002 18164 22008 18176
rect 22060 18164 22066 18216
rect 26237 18207 26295 18213
rect 26237 18173 26249 18207
rect 26283 18173 26295 18207
rect 26237 18167 26295 18173
rect 26421 18207 26479 18213
rect 26421 18173 26433 18207
rect 26467 18204 26479 18207
rect 27065 18207 27123 18213
rect 27065 18204 27077 18207
rect 26467 18176 27077 18204
rect 26467 18173 26479 18176
rect 26421 18167 26479 18173
rect 27065 18173 27077 18176
rect 27111 18173 27123 18207
rect 27065 18167 27123 18173
rect 22922 18136 22928 18148
rect 21468 18108 22928 18136
rect 22922 18096 22928 18108
rect 22980 18096 22986 18148
rect 23290 18136 23296 18148
rect 23251 18108 23296 18136
rect 23290 18096 23296 18108
rect 23348 18096 23354 18148
rect 26252 18136 26280 18167
rect 26252 18108 26464 18136
rect 26436 18080 26464 18108
rect 20165 18071 20223 18077
rect 20165 18068 20177 18071
rect 19444 18040 20177 18068
rect 20165 18037 20177 18040
rect 20211 18068 20223 18071
rect 20714 18068 20720 18080
rect 20211 18040 20720 18068
rect 20211 18037 20223 18040
rect 20165 18031 20223 18037
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 21174 18068 21180 18080
rect 21135 18040 21180 18068
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 25958 18068 25964 18080
rect 25919 18040 25964 18068
rect 25958 18028 25964 18040
rect 26016 18028 26022 18080
rect 26418 18028 26424 18080
rect 26476 18028 26482 18080
rect 28166 18068 28172 18080
rect 28127 18040 28172 18068
rect 28166 18028 28172 18040
rect 28224 18028 28230 18080
rect 1104 17978 28888 18000
rect 1104 17926 5582 17978
rect 5634 17926 5646 17978
rect 5698 17926 5710 17978
rect 5762 17926 5774 17978
rect 5826 17926 5838 17978
rect 5890 17926 14846 17978
rect 14898 17926 14910 17978
rect 14962 17926 14974 17978
rect 15026 17926 15038 17978
rect 15090 17926 15102 17978
rect 15154 17926 24110 17978
rect 24162 17926 24174 17978
rect 24226 17926 24238 17978
rect 24290 17926 24302 17978
rect 24354 17926 24366 17978
rect 24418 17926 28888 17978
rect 1104 17904 28888 17926
rect 6917 17867 6975 17873
rect 6917 17833 6929 17867
rect 6963 17864 6975 17867
rect 7098 17864 7104 17876
rect 6963 17836 7104 17864
rect 6963 17833 6975 17836
rect 6917 17827 6975 17833
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 7190 17824 7196 17876
rect 7248 17864 7254 17876
rect 8846 17864 8852 17876
rect 7248 17836 8852 17864
rect 7248 17824 7254 17836
rect 8846 17824 8852 17836
rect 8904 17864 8910 17876
rect 8904 17836 11744 17864
rect 8904 17824 8910 17836
rect 1394 17796 1400 17808
rect 1355 17768 1400 17796
rect 1394 17756 1400 17768
rect 1452 17756 1458 17808
rect 8938 17796 8944 17808
rect 7944 17768 8944 17796
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17629 7159 17663
rect 7101 17623 7159 17629
rect 7116 17592 7144 17623
rect 7190 17620 7196 17672
rect 7248 17660 7254 17672
rect 7944 17669 7972 17768
rect 8938 17756 8944 17768
rect 8996 17756 9002 17808
rect 8386 17728 8392 17740
rect 8036 17700 8392 17728
rect 7929 17663 7987 17669
rect 7248 17632 7293 17660
rect 7248 17620 7254 17632
rect 7929 17629 7941 17663
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8036 17592 8064 17700
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 11716 17737 11744 17836
rect 11974 17824 11980 17876
rect 12032 17864 12038 17876
rect 15194 17864 15200 17876
rect 12032 17836 15056 17864
rect 15155 17836 15200 17864
rect 12032 17824 12038 17836
rect 15028 17796 15056 17836
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 15654 17824 15660 17876
rect 15712 17864 15718 17876
rect 15841 17867 15899 17873
rect 15841 17864 15853 17867
rect 15712 17836 15853 17864
rect 15712 17824 15718 17836
rect 15841 17833 15853 17836
rect 15887 17833 15899 17867
rect 17494 17864 17500 17876
rect 15841 17827 15899 17833
rect 17144 17836 17500 17864
rect 16390 17796 16396 17808
rect 15028 17768 16396 17796
rect 16390 17756 16396 17768
rect 16448 17756 16454 17808
rect 11701 17731 11759 17737
rect 11701 17697 11713 17731
rect 11747 17697 11759 17731
rect 11701 17691 11759 17697
rect 11977 17731 12035 17737
rect 11977 17697 11989 17731
rect 12023 17728 12035 17731
rect 12158 17728 12164 17740
rect 12023 17700 12164 17728
rect 12023 17697 12035 17700
rect 11977 17691 12035 17697
rect 12158 17688 12164 17700
rect 12216 17688 12222 17740
rect 14090 17688 14096 17740
rect 14148 17728 14154 17740
rect 14148 17700 14780 17728
rect 14148 17688 14154 17700
rect 8294 17620 8300 17672
rect 8352 17660 8358 17672
rect 9214 17669 9220 17672
rect 8481 17663 8539 17669
rect 8481 17660 8493 17663
rect 8352 17632 8493 17660
rect 8352 17620 8358 17632
rect 8481 17629 8493 17632
rect 8527 17629 8539 17663
rect 8481 17623 8539 17629
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17629 8999 17663
rect 9208 17660 9220 17669
rect 9175 17632 9220 17660
rect 8941 17623 8999 17629
rect 9208 17623 9220 17632
rect 8956 17592 8984 17623
rect 9214 17620 9220 17623
rect 9272 17620 9278 17672
rect 12250 17660 12256 17672
rect 12211 17632 12256 17660
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 12434 17620 12440 17672
rect 12492 17660 12498 17672
rect 12529 17663 12587 17669
rect 12529 17660 12541 17663
rect 12492 17632 12541 17660
rect 12492 17620 12498 17632
rect 12529 17629 12541 17632
rect 12575 17629 12587 17663
rect 12529 17623 12587 17629
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17629 13599 17663
rect 13722 17660 13728 17672
rect 13683 17632 13728 17660
rect 13541 17623 13599 17629
rect 7116 17564 8064 17592
rect 8404 17564 8984 17592
rect 8404 17536 8432 17564
rect 11330 17552 11336 17604
rect 11388 17592 11394 17604
rect 12618 17592 12624 17604
rect 11388 17564 12624 17592
rect 11388 17552 11394 17564
rect 12618 17552 12624 17564
rect 12676 17552 12682 17604
rect 13556 17592 13584 17623
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 14369 17663 14427 17669
rect 14369 17629 14381 17663
rect 14415 17629 14427 17663
rect 14369 17623 14427 17629
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17629 14519 17663
rect 14461 17623 14519 17629
rect 14274 17592 14280 17604
rect 13556 17564 14280 17592
rect 14274 17552 14280 17564
rect 14332 17552 14338 17604
rect 7650 17484 7656 17536
rect 7708 17524 7714 17536
rect 7837 17527 7895 17533
rect 7837 17524 7849 17527
rect 7708 17496 7849 17524
rect 7708 17484 7714 17496
rect 7837 17493 7849 17496
rect 7883 17493 7895 17527
rect 8386 17524 8392 17536
rect 8347 17496 8392 17524
rect 7837 17487 7895 17493
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 9950 17484 9956 17536
rect 10008 17524 10014 17536
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 10008 17496 10333 17524
rect 10008 17484 10014 17496
rect 10321 17493 10333 17496
rect 10367 17493 10379 17527
rect 10778 17524 10784 17536
rect 10739 17496 10784 17524
rect 10321 17487 10379 17493
rect 10778 17484 10784 17496
rect 10836 17484 10842 17536
rect 11882 17484 11888 17536
rect 11940 17524 11946 17536
rect 12342 17524 12348 17536
rect 11940 17496 12348 17524
rect 11940 17484 11946 17496
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 13354 17524 13360 17536
rect 13315 17496 13360 17524
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 13446 17484 13452 17536
rect 13504 17524 13510 17536
rect 14093 17527 14151 17533
rect 14093 17524 14105 17527
rect 13504 17496 14105 17524
rect 13504 17484 13510 17496
rect 14093 17493 14105 17496
rect 14139 17493 14151 17527
rect 14384 17524 14412 17623
rect 14476 17592 14504 17623
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 14752 17669 14780 17700
rect 14826 17688 14832 17740
rect 14884 17728 14890 17740
rect 15562 17728 15568 17740
rect 14884 17700 15424 17728
rect 15523 17700 15568 17728
rect 14884 17688 14890 17700
rect 14737 17663 14795 17669
rect 14608 17632 14653 17660
rect 14608 17620 14614 17632
rect 14737 17629 14749 17663
rect 14783 17629 14795 17663
rect 15102 17660 15108 17672
rect 15063 17632 15108 17660
rect 14737 17623 14795 17629
rect 15102 17620 15108 17632
rect 15160 17620 15166 17672
rect 15396 17669 15424 17700
rect 15562 17688 15568 17700
rect 15620 17688 15626 17740
rect 17144 17737 17172 17836
rect 17494 17824 17500 17836
rect 17552 17824 17558 17876
rect 18506 17864 18512 17876
rect 18467 17836 18512 17864
rect 18506 17824 18512 17836
rect 18564 17824 18570 17876
rect 21910 17864 21916 17876
rect 19352 17836 21916 17864
rect 17129 17731 17187 17737
rect 15672 17700 17080 17728
rect 15381 17663 15439 17669
rect 15381 17629 15393 17663
rect 15427 17660 15439 17663
rect 15672 17660 15700 17700
rect 15427 17632 15700 17660
rect 15427 17629 15439 17632
rect 15381 17623 15439 17629
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 16025 17663 16083 17669
rect 16025 17660 16037 17663
rect 15896 17632 16037 17660
rect 15896 17620 15902 17632
rect 16025 17629 16037 17632
rect 16071 17629 16083 17663
rect 16206 17660 16212 17672
rect 16167 17632 16212 17660
rect 16025 17623 16083 17629
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17629 16359 17663
rect 16301 17623 16359 17629
rect 16316 17592 16344 17623
rect 16390 17620 16396 17672
rect 16448 17660 16454 17672
rect 16577 17663 16635 17669
rect 16577 17660 16589 17663
rect 16448 17632 16589 17660
rect 16448 17620 16454 17632
rect 16577 17629 16589 17632
rect 16623 17629 16635 17663
rect 16577 17623 16635 17629
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17660 16727 17663
rect 17052 17660 17080 17700
rect 17129 17697 17141 17731
rect 17175 17697 17187 17731
rect 18524 17728 18552 17824
rect 19245 17731 19303 17737
rect 19245 17728 19257 17731
rect 18524 17700 19257 17728
rect 17129 17691 17187 17697
rect 19245 17697 19257 17700
rect 19291 17697 19303 17731
rect 19245 17691 19303 17697
rect 16715 17632 16988 17660
rect 17052 17632 19288 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 16482 17592 16488 17604
rect 14476 17564 16068 17592
rect 16316 17564 16488 17592
rect 16040 17536 16068 17564
rect 16482 17552 16488 17564
rect 16540 17592 16546 17604
rect 16850 17592 16856 17604
rect 16540 17564 16712 17592
rect 16811 17564 16856 17592
rect 16540 17552 16546 17564
rect 15930 17524 15936 17536
rect 14384 17496 15936 17524
rect 14093 17487 14151 17493
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 16022 17484 16028 17536
rect 16080 17524 16086 17536
rect 16577 17527 16635 17533
rect 16577 17524 16589 17527
rect 16080 17496 16589 17524
rect 16080 17484 16086 17496
rect 16577 17493 16589 17496
rect 16623 17493 16635 17527
rect 16684 17524 16712 17564
rect 16850 17552 16856 17564
rect 16908 17552 16914 17604
rect 16960 17592 16988 17632
rect 19260 17604 19288 17632
rect 17034 17592 17040 17604
rect 16960 17564 17040 17592
rect 17034 17552 17040 17564
rect 17092 17552 17098 17604
rect 17218 17552 17224 17604
rect 17276 17592 17282 17604
rect 17374 17595 17432 17601
rect 17374 17592 17386 17595
rect 17276 17564 17386 17592
rect 17276 17552 17282 17564
rect 17374 17561 17386 17564
rect 17420 17561 17432 17595
rect 17374 17555 17432 17561
rect 17512 17564 18920 17592
rect 17512 17524 17540 17564
rect 16684 17496 17540 17524
rect 16577 17487 16635 17493
rect 18598 17484 18604 17536
rect 18656 17524 18662 17536
rect 18785 17527 18843 17533
rect 18785 17524 18797 17527
rect 18656 17496 18797 17524
rect 18656 17484 18662 17496
rect 18785 17493 18797 17496
rect 18831 17493 18843 17527
rect 18892 17524 18920 17564
rect 19242 17552 19248 17604
rect 19300 17552 19306 17604
rect 19352 17524 19380 17836
rect 21910 17824 21916 17836
rect 21968 17824 21974 17876
rect 23842 17824 23848 17876
rect 23900 17864 23906 17876
rect 24397 17867 24455 17873
rect 24397 17864 24409 17867
rect 23900 17836 24409 17864
rect 23900 17824 23906 17836
rect 24397 17833 24409 17836
rect 24443 17833 24455 17867
rect 25498 17864 25504 17876
rect 24397 17827 24455 17833
rect 25332 17836 25504 17864
rect 22005 17799 22063 17805
rect 22005 17796 22017 17799
rect 21652 17768 22017 17796
rect 21453 17731 21511 17737
rect 21453 17697 21465 17731
rect 21499 17728 21511 17731
rect 21652 17728 21680 17768
rect 22005 17765 22017 17768
rect 22051 17765 22063 17799
rect 22005 17759 22063 17765
rect 23109 17799 23167 17805
rect 23109 17765 23121 17799
rect 23155 17796 23167 17799
rect 25332 17796 25360 17836
rect 25498 17824 25504 17836
rect 25556 17824 25562 17876
rect 28074 17824 28080 17876
rect 28132 17864 28138 17876
rect 28353 17867 28411 17873
rect 28353 17864 28365 17867
rect 28132 17836 28365 17864
rect 28132 17824 28138 17836
rect 28353 17833 28365 17836
rect 28399 17833 28411 17867
rect 28353 17827 28411 17833
rect 23155 17768 25360 17796
rect 25409 17799 25467 17805
rect 23155 17765 23167 17768
rect 23109 17759 23167 17765
rect 25409 17765 25421 17799
rect 25455 17765 25467 17799
rect 25409 17759 25467 17765
rect 26053 17799 26111 17805
rect 26053 17765 26065 17799
rect 26099 17765 26111 17799
rect 26053 17759 26111 17765
rect 21499 17700 21680 17728
rect 21499 17697 21511 17700
rect 21453 17691 21511 17697
rect 21910 17688 21916 17740
rect 21968 17728 21974 17740
rect 21968 17700 22876 17728
rect 21968 17688 21974 17700
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17660 19579 17663
rect 19886 17660 19892 17672
rect 19567 17632 19892 17660
rect 19567 17629 19579 17632
rect 19521 17623 19579 17629
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 20162 17620 20168 17672
rect 20220 17660 20226 17672
rect 20533 17663 20591 17669
rect 20533 17660 20545 17663
rect 20220 17632 20545 17660
rect 20220 17620 20226 17632
rect 20533 17629 20545 17632
rect 20579 17629 20591 17663
rect 20714 17660 20720 17672
rect 20675 17632 20720 17660
rect 20533 17623 20591 17629
rect 20548 17592 20576 17623
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 20806 17620 20812 17672
rect 20864 17660 20870 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 20864 17632 21373 17660
rect 20864 17620 20870 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 22002 17660 22008 17672
rect 21963 17632 22008 17660
rect 21361 17623 21419 17629
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 22094 17620 22100 17672
rect 22152 17660 22158 17672
rect 22848 17669 22876 17700
rect 23658 17688 23664 17740
rect 23716 17728 23722 17740
rect 24486 17728 24492 17740
rect 23716 17700 24492 17728
rect 23716 17688 23722 17700
rect 24486 17688 24492 17700
rect 24544 17728 24550 17740
rect 24765 17731 24823 17737
rect 24765 17728 24777 17731
rect 24544 17700 24777 17728
rect 24544 17688 24550 17700
rect 24765 17697 24777 17700
rect 24811 17728 24823 17731
rect 24811 17700 25268 17728
rect 24811 17697 24823 17700
rect 24765 17691 24823 17697
rect 22189 17663 22247 17669
rect 22189 17660 22201 17663
rect 22152 17632 22201 17660
rect 22152 17620 22158 17632
rect 22189 17629 22201 17632
rect 22235 17629 22247 17663
rect 22189 17623 22247 17629
rect 22833 17663 22891 17669
rect 22833 17629 22845 17663
rect 22879 17629 22891 17663
rect 23106 17660 23112 17672
rect 23067 17632 23112 17660
rect 22833 17623 22891 17629
rect 23106 17620 23112 17632
rect 23164 17620 23170 17672
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17629 24639 17663
rect 24581 17623 24639 17629
rect 24673 17663 24731 17669
rect 24673 17629 24685 17663
rect 24719 17629 24731 17663
rect 24854 17660 24860 17672
rect 24815 17632 24860 17660
rect 24673 17623 24731 17629
rect 22020 17592 22048 17620
rect 20548 17564 22048 17592
rect 18892 17496 19380 17524
rect 20901 17527 20959 17533
rect 18785 17487 18843 17493
rect 20901 17493 20913 17527
rect 20947 17524 20959 17527
rect 20990 17524 20996 17536
rect 20947 17496 20996 17524
rect 20947 17493 20959 17496
rect 20901 17487 20959 17493
rect 20990 17484 20996 17496
rect 21048 17524 21054 17536
rect 21542 17524 21548 17536
rect 21048 17496 21548 17524
rect 21048 17484 21054 17496
rect 21542 17484 21548 17496
rect 21600 17484 21606 17536
rect 21729 17527 21787 17533
rect 21729 17493 21741 17527
rect 21775 17524 21787 17527
rect 23198 17524 23204 17536
rect 21775 17496 23204 17524
rect 21775 17493 21787 17496
rect 21729 17487 21787 17493
rect 23198 17484 23204 17496
rect 23256 17524 23262 17536
rect 24596 17524 24624 17623
rect 24688 17592 24716 17623
rect 24854 17620 24860 17632
rect 24912 17620 24918 17672
rect 25240 17669 25268 17700
rect 25225 17663 25283 17669
rect 25225 17629 25237 17663
rect 25271 17629 25283 17663
rect 25424 17660 25452 17759
rect 26068 17728 26096 17759
rect 26068 17700 27108 17728
rect 25777 17663 25835 17669
rect 25777 17660 25789 17663
rect 25424 17632 25789 17660
rect 25225 17623 25283 17629
rect 25777 17629 25789 17632
rect 25823 17629 25835 17663
rect 25777 17623 25835 17629
rect 25869 17663 25927 17669
rect 25869 17629 25881 17663
rect 25915 17660 25927 17663
rect 25958 17660 25964 17672
rect 25915 17632 25964 17660
rect 25915 17629 25927 17632
rect 25869 17623 25927 17629
rect 25958 17620 25964 17632
rect 26016 17620 26022 17672
rect 26234 17660 26240 17672
rect 26068 17632 26240 17660
rect 25130 17592 25136 17604
rect 24688 17564 25136 17592
rect 25130 17552 25136 17564
rect 25188 17552 25194 17604
rect 25317 17595 25375 17601
rect 25317 17561 25329 17595
rect 25363 17561 25375 17595
rect 25498 17592 25504 17604
rect 25459 17564 25504 17592
rect 25317 17555 25375 17561
rect 23256 17496 24624 17524
rect 25332 17524 25360 17555
rect 25498 17552 25504 17564
rect 25556 17552 25562 17604
rect 25682 17552 25688 17604
rect 25740 17592 25746 17604
rect 26068 17601 26096 17632
rect 26234 17620 26240 17632
rect 26292 17620 26298 17672
rect 26329 17663 26387 17669
rect 26329 17629 26341 17663
rect 26375 17660 26387 17663
rect 26418 17660 26424 17672
rect 26375 17632 26424 17660
rect 26375 17629 26387 17632
rect 26329 17623 26387 17629
rect 26418 17620 26424 17632
rect 26476 17620 26482 17672
rect 26513 17663 26571 17669
rect 26513 17629 26525 17663
rect 26559 17629 26571 17663
rect 26513 17623 26571 17629
rect 26053 17595 26111 17601
rect 26053 17592 26065 17595
rect 25740 17564 26065 17592
rect 25740 17552 25746 17564
rect 26053 17561 26065 17564
rect 26099 17561 26111 17595
rect 26528 17592 26556 17623
rect 26878 17620 26884 17672
rect 26936 17660 26942 17672
rect 26973 17663 27031 17669
rect 26973 17660 26985 17663
rect 26936 17632 26985 17660
rect 26936 17620 26942 17632
rect 26973 17629 26985 17632
rect 27019 17629 27031 17663
rect 27080 17660 27108 17700
rect 27229 17663 27287 17669
rect 27229 17660 27241 17663
rect 27080 17632 27241 17660
rect 26973 17623 27031 17629
rect 27229 17629 27241 17632
rect 27275 17629 27287 17663
rect 27229 17623 27287 17629
rect 26053 17555 26111 17561
rect 26206 17564 26556 17592
rect 25866 17524 25872 17536
rect 25332 17496 25872 17524
rect 23256 17484 23262 17496
rect 25866 17484 25872 17496
rect 25924 17524 25930 17536
rect 26206 17524 26234 17564
rect 26326 17524 26332 17536
rect 25924 17496 26234 17524
rect 26287 17496 26332 17524
rect 25924 17484 25930 17496
rect 26326 17484 26332 17496
rect 26384 17484 26390 17536
rect 1104 17434 28888 17456
rect 1104 17382 10214 17434
rect 10266 17382 10278 17434
rect 10330 17382 10342 17434
rect 10394 17382 10406 17434
rect 10458 17382 10470 17434
rect 10522 17382 19478 17434
rect 19530 17382 19542 17434
rect 19594 17382 19606 17434
rect 19658 17382 19670 17434
rect 19722 17382 19734 17434
rect 19786 17382 28888 17434
rect 1104 17360 28888 17382
rect 7374 17320 7380 17332
rect 7335 17292 7380 17320
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 11514 17320 11520 17332
rect 11475 17292 11520 17320
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 12437 17323 12495 17329
rect 11808 17292 12020 17320
rect 10781 17255 10839 17261
rect 10781 17221 10793 17255
rect 10827 17252 10839 17255
rect 11808 17252 11836 17292
rect 10827 17224 11836 17252
rect 10827 17221 10839 17224
rect 10781 17215 10839 17221
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17184 6055 17187
rect 6365 17187 6423 17193
rect 6365 17184 6377 17187
rect 6043 17156 6377 17184
rect 6043 17153 6055 17156
rect 5997 17147 6055 17153
rect 6365 17153 6377 17156
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 7190 17184 7196 17196
rect 6779 17156 7196 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 6564 17048 6592 17147
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 8656 17187 8714 17193
rect 8656 17153 8668 17187
rect 8702 17184 8714 17187
rect 8938 17184 8944 17196
rect 8702 17156 8944 17184
rect 8702 17153 8714 17156
rect 8656 17147 8714 17153
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17184 11023 17187
rect 11054 17184 11060 17196
rect 11011 17156 11060 17184
rect 11011 17153 11023 17156
rect 10965 17147 11023 17153
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 11330 17184 11336 17196
rect 11195 17156 11336 17184
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 11992 17193 12020 17292
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12618 17320 12624 17332
rect 12483 17292 12624 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 13078 17280 13084 17332
rect 13136 17320 13142 17332
rect 14826 17320 14832 17332
rect 13136 17292 14832 17320
rect 13136 17280 13142 17292
rect 14826 17280 14832 17292
rect 14884 17280 14890 17332
rect 15102 17280 15108 17332
rect 15160 17320 15166 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 15160 17292 15577 17320
rect 15160 17280 15166 17292
rect 15565 17289 15577 17292
rect 15611 17289 15623 17323
rect 16666 17320 16672 17332
rect 16627 17292 16672 17320
rect 15565 17283 15623 17289
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 17402 17320 17408 17332
rect 16960 17292 17408 17320
rect 12636 17252 12664 17280
rect 13633 17255 13691 17261
rect 13633 17252 13645 17255
rect 12636 17224 13645 17252
rect 13633 17221 13645 17224
rect 13679 17221 13691 17255
rect 13633 17215 13691 17221
rect 14550 17212 14556 17264
rect 14608 17252 14614 17264
rect 15746 17252 15752 17264
rect 14608 17224 15148 17252
rect 14608 17212 14614 17224
rect 11773 17187 11831 17193
rect 11773 17153 11785 17187
rect 11819 17153 11831 17187
rect 11773 17147 11831 17153
rect 11882 17187 11940 17193
rect 11882 17153 11894 17187
rect 11928 17153 11940 17187
rect 11882 17147 11940 17153
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 7098 17076 7104 17128
rect 7156 17116 7162 17128
rect 7469 17119 7527 17125
rect 7469 17116 7481 17119
rect 7156 17088 7481 17116
rect 7156 17076 7162 17088
rect 7469 17085 7481 17088
rect 7515 17085 7527 17119
rect 7650 17116 7656 17128
rect 7611 17088 7656 17116
rect 7469 17079 7527 17085
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 8386 17116 8392 17128
rect 8347 17088 8392 17116
rect 8386 17076 8392 17088
rect 8444 17076 8450 17128
rect 7009 17051 7067 17057
rect 7009 17048 7021 17051
rect 6564 17020 7021 17048
rect 7009 17017 7021 17020
rect 7055 17017 7067 17051
rect 7009 17011 7067 17017
rect 5813 16983 5871 16989
rect 5813 16949 5825 16983
rect 5859 16980 5871 16983
rect 5994 16980 6000 16992
rect 5859 16952 6000 16980
rect 5859 16949 5871 16952
rect 5813 16943 5871 16949
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 6730 16940 6736 16992
rect 6788 16980 6794 16992
rect 7668 16980 7696 17076
rect 9766 16980 9772 16992
rect 6788 16952 7696 16980
rect 9727 16952 9772 16980
rect 6788 16940 6794 16952
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10505 16983 10563 16989
rect 10505 16949 10517 16983
rect 10551 16980 10563 16983
rect 11799 16980 11827 17147
rect 11900 17116 11928 17147
rect 12066 17144 12072 17196
rect 12124 17184 12130 17196
rect 12161 17187 12219 17193
rect 12161 17184 12173 17187
rect 12124 17156 12173 17184
rect 12124 17144 12130 17156
rect 12161 17153 12173 17156
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17184 12679 17187
rect 12710 17184 12716 17196
rect 12667 17156 12716 17184
rect 12667 17153 12679 17156
rect 12621 17147 12679 17153
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 13078 17184 13084 17196
rect 13039 17156 13084 17184
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 13357 17187 13415 17193
rect 13357 17153 13369 17187
rect 13403 17184 13415 17187
rect 13446 17184 13452 17196
rect 13403 17156 13452 17184
rect 13403 17153 13415 17156
rect 13357 17147 13415 17153
rect 13446 17144 13452 17156
rect 13504 17144 13510 17196
rect 13722 17144 13728 17196
rect 13780 17184 13786 17196
rect 13817 17187 13875 17193
rect 13817 17184 13829 17187
rect 13780 17156 13829 17184
rect 13780 17144 13786 17156
rect 13817 17153 13829 17156
rect 13863 17153 13875 17187
rect 13817 17147 13875 17153
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14332 17156 14473 17184
rect 14332 17144 14338 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14642 17184 14648 17196
rect 14603 17156 14648 17184
rect 14461 17147 14519 17153
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 15120 17193 15148 17224
rect 15212 17224 15752 17252
rect 15212 17193 15240 17224
rect 15746 17212 15752 17224
rect 15804 17252 15810 17264
rect 15804 17224 16252 17252
rect 15804 17212 15810 17224
rect 16224 17196 16252 17224
rect 14921 17187 14979 17193
rect 14921 17153 14933 17187
rect 14967 17153 14979 17187
rect 14921 17147 14979 17153
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15197 17187 15255 17193
rect 15197 17153 15209 17187
rect 15243 17153 15255 17187
rect 15197 17147 15255 17153
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17153 15347 17187
rect 15289 17147 15347 17153
rect 12434 17116 12440 17128
rect 11900 17088 12440 17116
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 13906 17076 13912 17128
rect 13964 17116 13970 17128
rect 14936 17116 14964 17147
rect 13964 17088 14964 17116
rect 15304 17116 15332 17147
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 16025 17187 16083 17193
rect 16025 17184 16037 17187
rect 15528 17156 16037 17184
rect 15528 17144 15534 17156
rect 16025 17153 16037 17156
rect 16071 17153 16083 17187
rect 16206 17184 16212 17196
rect 16167 17156 16212 17184
rect 16025 17147 16083 17153
rect 16206 17144 16212 17156
rect 16264 17144 16270 17196
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 16960 17184 16988 17292
rect 17402 17280 17408 17292
rect 17460 17320 17466 17332
rect 19521 17323 19579 17329
rect 17460 17292 19104 17320
rect 17460 17280 17466 17292
rect 17126 17252 17132 17264
rect 17052 17224 17132 17252
rect 17052 17193 17080 17224
rect 17126 17212 17132 17224
rect 17184 17212 17190 17264
rect 19076 17252 19104 17292
rect 19521 17289 19533 17323
rect 19567 17320 19579 17323
rect 20714 17320 20720 17332
rect 19567 17292 20720 17320
rect 19567 17289 19579 17292
rect 19521 17283 19579 17289
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 26418 17280 26424 17332
rect 26476 17320 26482 17332
rect 26973 17323 27031 17329
rect 26973 17320 26985 17323
rect 26476 17292 26985 17320
rect 26476 17280 26482 17292
rect 26973 17289 26985 17292
rect 27019 17289 27031 17323
rect 28166 17320 28172 17332
rect 28127 17292 28172 17320
rect 26973 17283 27031 17289
rect 28166 17280 28172 17292
rect 28224 17280 28230 17332
rect 19794 17252 19800 17264
rect 17236 17224 18644 17252
rect 16347 17156 16988 17184
rect 17037 17187 17095 17193
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 17037 17153 17049 17187
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 17129 17119 17187 17125
rect 17129 17116 17141 17119
rect 15304 17088 17141 17116
rect 13964 17076 13970 17088
rect 17129 17085 17141 17088
rect 17175 17116 17187 17119
rect 17236 17116 17264 17224
rect 17865 17187 17923 17193
rect 17865 17153 17877 17187
rect 17911 17153 17923 17187
rect 17865 17147 17923 17153
rect 17175 17088 17264 17116
rect 17313 17119 17371 17125
rect 17175 17085 17187 17088
rect 17129 17079 17187 17085
rect 17313 17085 17325 17119
rect 17359 17116 17371 17119
rect 17770 17116 17776 17128
rect 17359 17088 17776 17116
rect 17359 17085 17371 17088
rect 17313 17079 17371 17085
rect 17770 17076 17776 17088
rect 17828 17076 17834 17128
rect 11882 17008 11888 17060
rect 11940 17048 11946 17060
rect 12897 17051 12955 17057
rect 12897 17048 12909 17051
rect 11940 17020 12909 17048
rect 11940 17008 11946 17020
rect 12897 17017 12909 17020
rect 12943 17017 12955 17051
rect 12897 17011 12955 17017
rect 13265 17051 13323 17057
rect 13265 17017 13277 17051
rect 13311 17048 13323 17051
rect 17681 17051 17739 17057
rect 17681 17048 17693 17051
rect 13311 17020 17693 17048
rect 13311 17017 13323 17020
rect 13265 17011 13323 17017
rect 17681 17017 17693 17020
rect 17727 17017 17739 17051
rect 17681 17011 17739 17017
rect 11974 16980 11980 16992
rect 10551 16952 11980 16980
rect 10551 16949 10563 16952
rect 10505 16943 10563 16949
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 13998 16980 14004 16992
rect 13959 16952 14004 16980
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 14274 16980 14280 16992
rect 14235 16952 14280 16980
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 14458 16940 14464 16992
rect 14516 16980 14522 16992
rect 15841 16983 15899 16989
rect 15841 16980 15853 16983
rect 14516 16952 15853 16980
rect 14516 16940 14522 16952
rect 15841 16949 15853 16952
rect 15887 16949 15899 16983
rect 15841 16943 15899 16949
rect 16206 16940 16212 16992
rect 16264 16980 16270 16992
rect 17880 16980 17908 17147
rect 17954 17144 17960 17196
rect 18012 17184 18018 17196
rect 18012 17156 18057 17184
rect 18012 17144 18018 17156
rect 18616 17116 18644 17224
rect 19076 17224 19800 17252
rect 19076 17193 19104 17224
rect 19794 17212 19800 17224
rect 19852 17212 19858 17264
rect 19978 17252 19984 17264
rect 19904 17224 19984 17252
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17153 19119 17187
rect 19334 17184 19340 17196
rect 19295 17156 19340 17184
rect 19061 17147 19119 17153
rect 19334 17144 19340 17156
rect 19392 17144 19398 17196
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17184 19579 17187
rect 19702 17184 19708 17196
rect 19567 17156 19708 17184
rect 19567 17153 19579 17156
rect 19521 17147 19579 17153
rect 19702 17144 19708 17156
rect 19760 17184 19766 17196
rect 19904 17184 19932 17224
rect 19978 17212 19984 17224
rect 20036 17212 20042 17264
rect 20254 17252 20260 17264
rect 20167 17224 20260 17252
rect 20254 17212 20260 17224
rect 20312 17252 20318 17264
rect 20809 17255 20867 17261
rect 20809 17252 20821 17255
rect 20312 17224 20821 17252
rect 20312 17212 20318 17224
rect 20809 17221 20821 17224
rect 20855 17221 20867 17255
rect 20809 17215 20867 17221
rect 22462 17212 22468 17264
rect 22520 17252 22526 17264
rect 25774 17252 25780 17264
rect 22520 17224 23244 17252
rect 22520 17212 22526 17224
rect 20070 17184 20076 17196
rect 19760 17156 19932 17184
rect 20031 17156 20076 17184
rect 19760 17144 19766 17156
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 20714 17184 20720 17196
rect 20675 17156 20720 17184
rect 20714 17144 20720 17156
rect 20772 17144 20778 17196
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17153 20959 17187
rect 20901 17147 20959 17153
rect 19199 17119 19257 17125
rect 19199 17116 19211 17119
rect 18616 17088 19211 17116
rect 19199 17085 19211 17088
rect 19245 17116 19257 17119
rect 19886 17116 19892 17128
rect 19245 17088 19892 17116
rect 19245 17085 19257 17088
rect 19199 17079 19257 17085
rect 19886 17076 19892 17088
rect 19944 17116 19950 17128
rect 20916 17116 20944 17147
rect 21910 17144 21916 17196
rect 21968 17184 21974 17196
rect 22281 17187 22339 17193
rect 22281 17184 22293 17187
rect 21968 17156 22293 17184
rect 21968 17144 21974 17156
rect 22281 17153 22293 17156
rect 22327 17153 22339 17187
rect 22925 17187 22983 17193
rect 22925 17184 22937 17187
rect 22281 17147 22339 17153
rect 22572 17156 22937 17184
rect 19944 17088 20944 17116
rect 19944 17076 19950 17088
rect 21358 17076 21364 17128
rect 21416 17116 21422 17128
rect 22189 17119 22247 17125
rect 22189 17116 22201 17119
rect 21416 17088 22201 17116
rect 21416 17076 21422 17088
rect 22189 17085 22201 17088
rect 22235 17116 22247 17119
rect 22572 17116 22600 17156
rect 22925 17153 22937 17156
rect 22971 17184 22983 17187
rect 23106 17184 23112 17196
rect 22971 17156 23112 17184
rect 22971 17153 22983 17156
rect 22925 17147 22983 17153
rect 23106 17144 23112 17156
rect 23164 17144 23170 17196
rect 23216 17193 23244 17224
rect 24412 17224 25780 17252
rect 23201 17187 23259 17193
rect 23201 17153 23213 17187
rect 23247 17153 23259 17187
rect 23201 17147 23259 17153
rect 22235 17088 22600 17116
rect 22649 17119 22707 17125
rect 22235 17085 22247 17088
rect 22189 17079 22247 17085
rect 22649 17085 22661 17119
rect 22695 17116 22707 17119
rect 24412 17116 24440 17224
rect 24578 17184 24584 17196
rect 24539 17156 24584 17184
rect 24578 17144 24584 17156
rect 24636 17144 24642 17196
rect 24872 17193 24900 17224
rect 25774 17212 25780 17224
rect 25832 17212 25838 17264
rect 26605 17255 26663 17261
rect 26605 17221 26617 17255
rect 26651 17252 26663 17255
rect 27433 17255 27491 17261
rect 27433 17252 27445 17255
rect 26651 17224 27445 17252
rect 26651 17221 26663 17224
rect 26605 17215 26663 17221
rect 27433 17221 27445 17224
rect 27479 17252 27491 17255
rect 28258 17252 28264 17264
rect 27479 17224 28264 17252
rect 27479 17221 27491 17224
rect 27433 17215 27491 17221
rect 28258 17212 28264 17224
rect 28316 17212 28322 17264
rect 24857 17187 24915 17193
rect 24857 17153 24869 17187
rect 24903 17153 24915 17187
rect 24857 17147 24915 17153
rect 24946 17144 24952 17196
rect 25004 17184 25010 17196
rect 25314 17184 25320 17196
rect 25004 17156 25320 17184
rect 25004 17144 25010 17156
rect 25314 17144 25320 17156
rect 25372 17184 25378 17196
rect 25409 17187 25467 17193
rect 25409 17184 25421 17187
rect 25372 17156 25421 17184
rect 25372 17144 25378 17156
rect 25409 17153 25421 17156
rect 25455 17153 25467 17187
rect 26145 17187 26203 17193
rect 26145 17184 26157 17187
rect 25409 17147 25467 17153
rect 25516 17156 26157 17184
rect 22695 17088 24440 17116
rect 22695 17085 22707 17088
rect 22649 17079 22707 17085
rect 24486 17076 24492 17128
rect 24544 17116 24550 17128
rect 24673 17119 24731 17125
rect 24673 17116 24685 17119
rect 24544 17088 24685 17116
rect 24544 17076 24550 17088
rect 24673 17085 24685 17088
rect 24719 17085 24731 17119
rect 24673 17079 24731 17085
rect 24765 17119 24823 17125
rect 24765 17085 24777 17119
rect 24811 17085 24823 17119
rect 25130 17116 25136 17128
rect 24765 17079 24823 17085
rect 24964 17088 25136 17116
rect 20441 17051 20499 17057
rect 20441 17017 20453 17051
rect 20487 17048 20499 17051
rect 21910 17048 21916 17060
rect 20487 17020 21916 17048
rect 20487 17017 20499 17020
rect 20441 17011 20499 17017
rect 21910 17008 21916 17020
rect 21968 17048 21974 17060
rect 22370 17048 22376 17060
rect 21968 17020 22376 17048
rect 21968 17008 21974 17020
rect 22370 17008 22376 17020
rect 22428 17008 22434 17060
rect 24780 17048 24808 17079
rect 24964 17048 24992 17088
rect 25130 17076 25136 17088
rect 25188 17116 25194 17128
rect 25516 17116 25544 17156
rect 26145 17153 26157 17156
rect 26191 17153 26203 17187
rect 26145 17147 26203 17153
rect 27801 17187 27859 17193
rect 27801 17153 27813 17187
rect 27847 17184 27859 17187
rect 28350 17184 28356 17196
rect 27847 17156 28356 17184
rect 27847 17153 27859 17156
rect 27801 17147 27859 17153
rect 28350 17144 28356 17156
rect 28408 17144 28414 17196
rect 25188 17088 25544 17116
rect 25188 17076 25194 17088
rect 26050 17076 26056 17128
rect 26108 17116 26114 17128
rect 26237 17119 26295 17125
rect 26237 17116 26249 17119
rect 26108 17088 26249 17116
rect 26108 17076 26114 17088
rect 26237 17085 26249 17088
rect 26283 17116 26295 17119
rect 26283 17088 27108 17116
rect 26283 17085 26295 17088
rect 26237 17079 26295 17085
rect 24780 17020 24992 17048
rect 25041 17051 25099 17057
rect 25041 17017 25053 17051
rect 25087 17048 25099 17051
rect 26418 17048 26424 17060
rect 25087 17020 26424 17048
rect 25087 17017 25099 17020
rect 25041 17011 25099 17017
rect 26418 17008 26424 17020
rect 26476 17008 26482 17060
rect 27080 17057 27108 17088
rect 27065 17051 27123 17057
rect 27065 17017 27077 17051
rect 27111 17017 27123 17051
rect 27065 17011 27123 17017
rect 16264 16952 17908 16980
rect 18417 16983 18475 16989
rect 16264 16940 16270 16952
rect 18417 16949 18429 16983
rect 18463 16980 18475 16983
rect 18690 16980 18696 16992
rect 18463 16952 18696 16980
rect 18463 16949 18475 16952
rect 18417 16943 18475 16949
rect 18690 16940 18696 16952
rect 18748 16940 18754 16992
rect 18785 16983 18843 16989
rect 18785 16949 18797 16983
rect 18831 16980 18843 16983
rect 18874 16980 18880 16992
rect 18831 16952 18880 16980
rect 18831 16949 18843 16952
rect 18785 16943 18843 16949
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 20714 16940 20720 16992
rect 20772 16980 20778 16992
rect 21082 16980 21088 16992
rect 20772 16952 21088 16980
rect 20772 16940 20778 16952
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 23293 16983 23351 16989
rect 23293 16949 23305 16983
rect 23339 16980 23351 16983
rect 23382 16980 23388 16992
rect 23339 16952 23388 16980
rect 23339 16949 23351 16952
rect 23293 16943 23351 16949
rect 23382 16940 23388 16952
rect 23440 16940 23446 16992
rect 23477 16983 23535 16989
rect 23477 16949 23489 16983
rect 23523 16980 23535 16983
rect 24946 16980 24952 16992
rect 23523 16952 24952 16980
rect 23523 16949 23535 16952
rect 23477 16943 23535 16949
rect 24946 16940 24952 16952
rect 25004 16940 25010 16992
rect 25406 16940 25412 16992
rect 25464 16980 25470 16992
rect 25501 16983 25559 16989
rect 25501 16980 25513 16983
rect 25464 16952 25513 16980
rect 25464 16940 25470 16952
rect 25501 16949 25513 16952
rect 25547 16980 25559 16983
rect 25682 16980 25688 16992
rect 25547 16952 25688 16980
rect 25547 16949 25559 16952
rect 25501 16943 25559 16949
rect 25682 16940 25688 16952
rect 25740 16940 25746 16992
rect 25961 16983 26019 16989
rect 25961 16949 25973 16983
rect 26007 16980 26019 16983
rect 26142 16980 26148 16992
rect 26007 16952 26148 16980
rect 26007 16949 26019 16952
rect 25961 16943 26019 16949
rect 26142 16940 26148 16952
rect 26200 16940 26206 16992
rect 1104 16890 28888 16912
rect 1104 16838 5582 16890
rect 5634 16838 5646 16890
rect 5698 16838 5710 16890
rect 5762 16838 5774 16890
rect 5826 16838 5838 16890
rect 5890 16838 14846 16890
rect 14898 16838 14910 16890
rect 14962 16838 14974 16890
rect 15026 16838 15038 16890
rect 15090 16838 15102 16890
rect 15154 16838 24110 16890
rect 24162 16838 24174 16890
rect 24226 16838 24238 16890
rect 24290 16838 24302 16890
rect 24354 16838 24366 16890
rect 24418 16838 28888 16890
rect 1104 16816 28888 16838
rect 8386 16776 8392 16788
rect 5736 16748 8392 16776
rect 5736 16649 5764 16748
rect 8386 16736 8392 16748
rect 8444 16736 8450 16788
rect 8938 16776 8944 16788
rect 8899 16748 8944 16776
rect 8938 16736 8944 16748
rect 8996 16736 9002 16788
rect 11333 16779 11391 16785
rect 11333 16745 11345 16779
rect 11379 16776 11391 16779
rect 11422 16776 11428 16788
rect 11379 16748 11428 16776
rect 11379 16745 11391 16748
rect 11333 16739 11391 16745
rect 11422 16736 11428 16748
rect 11480 16736 11486 16788
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 13081 16779 13139 16785
rect 13081 16776 13093 16779
rect 12860 16748 13093 16776
rect 12860 16736 12866 16748
rect 13081 16745 13093 16748
rect 13127 16745 13139 16779
rect 13081 16739 13139 16745
rect 13354 16736 13360 16788
rect 13412 16776 13418 16788
rect 13449 16779 13507 16785
rect 13449 16776 13461 16779
rect 13412 16748 13461 16776
rect 13412 16736 13418 16748
rect 13449 16745 13461 16748
rect 13495 16745 13507 16779
rect 13449 16739 13507 16745
rect 15286 16736 15292 16788
rect 15344 16776 15350 16788
rect 16206 16776 16212 16788
rect 15344 16748 16212 16776
rect 15344 16736 15350 16748
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 20438 16776 20444 16788
rect 16316 16748 20444 16776
rect 8404 16708 8432 16736
rect 16316 16720 16344 16748
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 23842 16736 23848 16788
rect 23900 16776 23906 16788
rect 25406 16776 25412 16788
rect 23900 16748 25412 16776
rect 23900 16736 23906 16748
rect 25406 16736 25412 16748
rect 25464 16736 25470 16788
rect 28258 16776 28264 16788
rect 28219 16748 28264 16776
rect 28258 16736 28264 16748
rect 28316 16736 28322 16788
rect 8570 16708 8576 16720
rect 8404 16680 8576 16708
rect 8570 16668 8576 16680
rect 8628 16708 8634 16720
rect 8628 16680 9996 16708
rect 8628 16668 8634 16680
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 5721 16643 5779 16649
rect 5721 16640 5733 16643
rect 2823 16612 5733 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 5721 16609 5733 16612
rect 5767 16609 5779 16643
rect 5721 16603 5779 16609
rect 7374 16600 7380 16652
rect 7432 16640 7438 16652
rect 9968 16649 9996 16680
rect 11698 16668 11704 16720
rect 11756 16708 11762 16720
rect 11756 16680 12092 16708
rect 11756 16668 11762 16680
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 7432 16612 8309 16640
rect 7432 16600 7438 16612
rect 8297 16609 8309 16612
rect 8343 16609 8355 16643
rect 8297 16603 8355 16609
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16609 8447 16643
rect 8389 16603 8447 16609
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16609 10011 16643
rect 9953 16603 10011 16609
rect 5994 16581 6000 16584
rect 5988 16572 6000 16581
rect 5955 16544 6000 16572
rect 5988 16535 6000 16544
rect 5994 16532 6000 16535
rect 6052 16532 6058 16584
rect 8202 16532 8208 16584
rect 8260 16572 8266 16584
rect 8404 16572 8432 16603
rect 9122 16572 9128 16584
rect 8260 16544 8432 16572
rect 9083 16544 9128 16572
rect 8260 16532 8266 16544
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 12064 16581 12092 16680
rect 12710 16668 12716 16720
rect 12768 16708 12774 16720
rect 13630 16708 13636 16720
rect 12768 16680 13636 16708
rect 12768 16668 12774 16680
rect 13630 16668 13636 16680
rect 13688 16708 13694 16720
rect 14182 16708 14188 16720
rect 13688 16680 14188 16708
rect 13688 16668 13694 16680
rect 14182 16668 14188 16680
rect 14240 16668 14246 16720
rect 14550 16668 14556 16720
rect 14608 16668 14614 16720
rect 16298 16708 16304 16720
rect 16259 16680 16304 16708
rect 16298 16668 16304 16680
rect 16356 16668 16362 16720
rect 17218 16708 17224 16720
rect 17179 16680 17224 16708
rect 17218 16668 17224 16680
rect 17276 16668 17282 16720
rect 20349 16711 20407 16717
rect 20349 16677 20361 16711
rect 20395 16708 20407 16711
rect 20898 16708 20904 16720
rect 20395 16680 20904 16708
rect 20395 16677 20407 16680
rect 20349 16671 20407 16677
rect 20898 16668 20904 16680
rect 20956 16708 20962 16720
rect 21818 16708 21824 16720
rect 20956 16680 21824 16708
rect 20956 16668 20962 16680
rect 21818 16668 21824 16680
rect 21876 16668 21882 16720
rect 22002 16708 22008 16720
rect 21963 16680 22008 16708
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 25130 16668 25136 16720
rect 25188 16708 25194 16720
rect 25777 16711 25835 16717
rect 25777 16708 25789 16711
rect 25188 16680 25789 16708
rect 25188 16668 25194 16680
rect 25777 16677 25789 16680
rect 25823 16708 25835 16711
rect 26234 16708 26240 16720
rect 25823 16680 26240 16708
rect 25823 16677 25835 16680
rect 25777 16671 25835 16677
rect 26234 16668 26240 16680
rect 26292 16668 26298 16720
rect 26421 16711 26479 16717
rect 26421 16677 26433 16711
rect 26467 16677 26479 16711
rect 26421 16671 26479 16677
rect 12802 16640 12808 16652
rect 12715 16612 12808 16640
rect 12802 16600 12808 16612
rect 12860 16640 12866 16652
rect 12986 16640 12992 16652
rect 12860 16612 12992 16640
rect 12860 16600 12866 16612
rect 12986 16600 12992 16612
rect 13044 16600 13050 16652
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13587 16612 14105 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14568 16640 14596 16668
rect 17494 16640 17500 16652
rect 14568 16612 14780 16640
rect 17455 16612 17500 16640
rect 14093 16603 14151 16609
rect 11839 16575 11897 16581
rect 11839 16541 11851 16575
rect 11885 16572 11897 16575
rect 11974 16572 12032 16578
rect 11885 16541 11908 16572
rect 11839 16535 11908 16541
rect 11880 16516 11908 16535
rect 11974 16538 11986 16572
rect 12020 16538 12032 16572
rect 12064 16575 12127 16581
rect 12064 16546 12081 16575
rect 11974 16532 12032 16538
rect 12069 16541 12081 16546
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12253 16575 12311 16581
rect 12253 16541 12265 16575
rect 12299 16572 12311 16575
rect 12342 16572 12348 16584
rect 12299 16544 12348 16572
rect 12299 16541 12311 16544
rect 12253 16535 12311 16541
rect 12342 16532 12348 16544
rect 12400 16532 12406 16584
rect 13078 16532 13084 16584
rect 13136 16572 13142 16584
rect 13265 16575 13323 16581
rect 13265 16572 13277 16575
rect 13136 16544 13277 16572
rect 13136 16532 13142 16544
rect 13265 16541 13277 16544
rect 13311 16541 13323 16575
rect 13265 16535 13323 16541
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 14461 16575 14519 16581
rect 14461 16541 14473 16575
rect 14507 16541 14519 16575
rect 14461 16535 14519 16541
rect 2532 16507 2590 16513
rect 2532 16473 2544 16507
rect 2578 16504 2590 16507
rect 10220 16507 10278 16513
rect 2578 16476 9904 16504
rect 2578 16473 2590 16476
rect 2532 16467 2590 16473
rect 1397 16439 1455 16445
rect 1397 16405 1409 16439
rect 1443 16436 1455 16439
rect 1486 16436 1492 16448
rect 1443 16408 1492 16436
rect 1443 16405 1455 16408
rect 1397 16399 1455 16405
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 7098 16436 7104 16448
rect 7059 16408 7104 16436
rect 7098 16396 7104 16408
rect 7156 16396 7162 16448
rect 7834 16436 7840 16448
rect 7795 16408 7840 16436
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 8205 16439 8263 16445
rect 8205 16405 8217 16439
rect 8251 16436 8263 16439
rect 9766 16436 9772 16448
rect 8251 16408 9772 16436
rect 8251 16405 8263 16408
rect 8205 16399 8263 16405
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 9876 16436 9904 16476
rect 10220 16473 10232 16507
rect 10266 16504 10278 16507
rect 11609 16507 11667 16513
rect 11609 16504 11621 16507
rect 10266 16476 11621 16504
rect 10266 16473 10278 16476
rect 10220 16467 10278 16473
rect 11609 16473 11621 16476
rect 11655 16473 11667 16507
rect 11880 16476 11888 16516
rect 11609 16467 11667 16473
rect 11882 16464 11888 16476
rect 11940 16464 11946 16516
rect 11790 16436 11796 16448
rect 9876 16408 11796 16436
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 11989 16436 12017 16532
rect 12434 16504 12440 16516
rect 12064 16476 12440 16504
rect 12064 16436 12092 16476
rect 12434 16464 12440 16476
rect 12492 16464 12498 16516
rect 11989 16408 12092 16436
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 14384 16436 14412 16535
rect 14476 16504 14504 16535
rect 14550 16532 14556 16584
rect 14608 16572 14614 16584
rect 14752 16581 14780 16612
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 19242 16640 19248 16652
rect 19203 16612 19248 16640
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 19702 16600 19708 16652
rect 19760 16640 19766 16652
rect 19886 16640 19892 16652
rect 19760 16612 19892 16640
rect 19760 16600 19766 16612
rect 19886 16600 19892 16612
rect 19944 16600 19950 16652
rect 20073 16643 20131 16649
rect 20073 16609 20085 16643
rect 20119 16640 20131 16643
rect 20254 16640 20260 16652
rect 20119 16612 20260 16640
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 24504 16612 24716 16640
rect 14737 16575 14795 16581
rect 14608 16544 14653 16572
rect 14608 16532 14614 16544
rect 14737 16541 14749 16575
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 16758 16532 16764 16584
rect 16816 16572 16822 16584
rect 17037 16575 17095 16581
rect 17037 16572 17049 16575
rect 16816 16544 17049 16572
rect 16816 16532 16822 16544
rect 17037 16541 17049 16544
rect 17083 16541 17095 16575
rect 17037 16535 17095 16541
rect 19334 16532 19340 16584
rect 19392 16532 19398 16584
rect 19794 16532 19800 16584
rect 19852 16572 19858 16584
rect 19981 16575 20039 16581
rect 19981 16572 19993 16575
rect 19852 16544 19993 16572
rect 19852 16532 19858 16544
rect 19981 16541 19993 16544
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 21634 16532 21640 16584
rect 21692 16572 21698 16584
rect 21729 16575 21787 16581
rect 21729 16572 21741 16575
rect 21692 16544 21741 16572
rect 21692 16532 21698 16544
rect 21729 16541 21741 16544
rect 21775 16541 21787 16575
rect 21729 16535 21787 16541
rect 24397 16575 24455 16581
rect 24397 16541 24409 16575
rect 24443 16572 24455 16575
rect 24504 16572 24532 16612
rect 24443 16544 24532 16572
rect 24581 16575 24639 16581
rect 24443 16541 24455 16544
rect 24397 16535 24455 16541
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24688 16572 24716 16612
rect 25038 16572 25044 16584
rect 24688 16544 25044 16572
rect 24581 16535 24639 16541
rect 15010 16504 15016 16516
rect 14476 16476 14596 16504
rect 14971 16476 15016 16504
rect 13872 16408 14412 16436
rect 14568 16436 14596 16476
rect 15010 16464 15016 16476
rect 15068 16464 15074 16516
rect 17764 16507 17822 16513
rect 17764 16473 17776 16507
rect 17810 16504 17822 16507
rect 18782 16504 18788 16516
rect 17810 16476 18788 16504
rect 17810 16473 17822 16476
rect 17764 16467 17822 16473
rect 18782 16464 18788 16476
rect 18840 16464 18846 16516
rect 19352 16504 19380 16532
rect 18892 16476 19380 16504
rect 19429 16507 19487 16513
rect 15194 16436 15200 16448
rect 14568 16408 15200 16436
rect 13872 16396 13878 16408
rect 15194 16396 15200 16408
rect 15252 16436 15258 16448
rect 15746 16436 15752 16448
rect 15252 16408 15752 16436
rect 15252 16396 15258 16408
rect 15746 16396 15752 16408
rect 15804 16396 15810 16448
rect 18892 16445 18920 16476
rect 19429 16473 19441 16507
rect 19475 16504 19487 16507
rect 21174 16504 21180 16516
rect 19475 16476 21180 16504
rect 19475 16473 19487 16476
rect 19429 16467 19487 16473
rect 21174 16464 21180 16476
rect 21232 16464 21238 16516
rect 22005 16507 22063 16513
rect 22005 16504 22017 16507
rect 21284 16476 22017 16504
rect 18877 16439 18935 16445
rect 18877 16405 18889 16439
rect 18923 16405 18935 16439
rect 18877 16399 18935 16405
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 21284 16436 21312 16476
rect 22005 16473 22017 16476
rect 22051 16473 22063 16507
rect 22005 16467 22063 16473
rect 20772 16408 21312 16436
rect 20772 16396 20778 16408
rect 21450 16396 21456 16448
rect 21508 16436 21514 16448
rect 21821 16439 21879 16445
rect 21821 16436 21833 16439
rect 21508 16408 21833 16436
rect 21508 16396 21514 16408
rect 21821 16405 21833 16408
rect 21867 16405 21879 16439
rect 21821 16399 21879 16405
rect 23474 16396 23480 16448
rect 23532 16436 23538 16448
rect 24489 16439 24547 16445
rect 24489 16436 24501 16439
rect 23532 16408 24501 16436
rect 23532 16396 23538 16408
rect 24489 16405 24501 16408
rect 24535 16405 24547 16439
rect 24596 16436 24624 16535
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 25222 16572 25228 16584
rect 25183 16544 25228 16572
rect 25222 16532 25228 16544
rect 25280 16532 25286 16584
rect 26142 16572 26148 16584
rect 26103 16544 26148 16572
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 26237 16575 26295 16581
rect 26237 16541 26249 16575
rect 26283 16572 26295 16575
rect 26326 16572 26332 16584
rect 26283 16544 26332 16572
rect 26283 16541 26295 16544
rect 26237 16535 26295 16541
rect 26326 16532 26332 16544
rect 26384 16532 26390 16584
rect 26436 16572 26464 16671
rect 26878 16572 26884 16584
rect 26436 16544 26740 16572
rect 26839 16544 26884 16572
rect 26418 16504 26424 16516
rect 26379 16476 26424 16504
rect 26418 16464 26424 16476
rect 26476 16464 26482 16516
rect 26712 16504 26740 16544
rect 26878 16532 26884 16544
rect 26936 16532 26942 16584
rect 27126 16507 27184 16513
rect 27126 16504 27138 16507
rect 26712 16476 27138 16504
rect 27126 16473 27138 16476
rect 27172 16473 27184 16507
rect 27126 16467 27184 16473
rect 25409 16439 25467 16445
rect 25409 16436 25421 16439
rect 24596 16408 25421 16436
rect 24489 16399 24547 16405
rect 25409 16405 25421 16408
rect 25455 16436 25467 16439
rect 25498 16436 25504 16448
rect 25455 16408 25504 16436
rect 25455 16405 25467 16408
rect 25409 16399 25467 16405
rect 25498 16396 25504 16408
rect 25556 16396 25562 16448
rect 1104 16346 28888 16368
rect 1104 16294 10214 16346
rect 10266 16294 10278 16346
rect 10330 16294 10342 16346
rect 10394 16294 10406 16346
rect 10458 16294 10470 16346
rect 10522 16294 19478 16346
rect 19530 16294 19542 16346
rect 19594 16294 19606 16346
rect 19658 16294 19670 16346
rect 19722 16294 19734 16346
rect 19786 16294 28888 16346
rect 1104 16272 28888 16294
rect 8389 16235 8447 16241
rect 8389 16201 8401 16235
rect 8435 16232 8447 16235
rect 9122 16232 9128 16244
rect 8435 16204 9128 16232
rect 8435 16201 8447 16204
rect 8389 16195 8447 16201
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 9950 16232 9956 16244
rect 9911 16204 9956 16232
rect 9950 16192 9956 16204
rect 10008 16192 10014 16244
rect 11146 16232 11152 16244
rect 11107 16204 11152 16232
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 12897 16235 12955 16241
rect 12897 16201 12909 16235
rect 12943 16232 12955 16235
rect 13722 16232 13728 16244
rect 12943 16204 13728 16232
rect 12943 16201 12955 16204
rect 12897 16195 12955 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 16945 16235 17003 16241
rect 16945 16232 16957 16235
rect 13872 16204 16957 16232
rect 13872 16192 13878 16204
rect 16945 16201 16957 16204
rect 16991 16232 17003 16235
rect 16991 16204 17816 16232
rect 16991 16201 17003 16204
rect 16945 16195 17003 16201
rect 10686 16124 10692 16176
rect 10744 16164 10750 16176
rect 15010 16164 15016 16176
rect 10744 16136 15016 16164
rect 10744 16124 10750 16136
rect 15010 16124 15016 16136
rect 15068 16124 15074 16176
rect 17678 16164 17684 16176
rect 16868 16136 17684 16164
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 5629 16099 5687 16105
rect 5629 16065 5641 16099
rect 5675 16096 5687 16099
rect 5902 16096 5908 16108
rect 5675 16068 5908 16096
rect 5675 16065 5687 16068
rect 5629 16059 5687 16065
rect 5902 16056 5908 16068
rect 5960 16056 5966 16108
rect 7558 16096 7564 16108
rect 7519 16068 7564 16096
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 8205 16099 8263 16105
rect 8205 16096 8217 16099
rect 7892 16068 8217 16096
rect 7892 16056 7898 16068
rect 8205 16065 8217 16068
rect 8251 16065 8263 16099
rect 8205 16059 8263 16065
rect 9033 16099 9091 16105
rect 9033 16065 9045 16099
rect 9079 16096 9091 16099
rect 9861 16099 9919 16105
rect 9079 16068 9536 16096
rect 9079 16065 9091 16068
rect 9033 16059 9091 16065
rect 7377 16031 7435 16037
rect 7377 15997 7389 16031
rect 7423 16028 7435 16031
rect 8021 16031 8079 16037
rect 8021 16028 8033 16031
rect 7423 16000 8033 16028
rect 7423 15997 7435 16000
rect 7377 15991 7435 15997
rect 8021 15997 8033 16000
rect 8067 16028 8079 16031
rect 8849 16031 8907 16037
rect 8849 16028 8861 16031
rect 8067 16000 8861 16028
rect 8067 15997 8079 16000
rect 8021 15991 8079 15997
rect 8849 15997 8861 16000
rect 8895 16028 8907 16031
rect 9214 16028 9220 16040
rect 8895 16000 9220 16028
rect 8895 15997 8907 16000
rect 8849 15991 8907 15997
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 9508 15969 9536 16068
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 11054 16096 11060 16108
rect 9907 16068 11060 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 11790 16105 11796 16108
rect 11784 16059 11796 16105
rect 11848 16096 11854 16108
rect 11848 16068 11884 16096
rect 11790 16056 11796 16059
rect 11848 16056 11854 16068
rect 13078 16056 13084 16108
rect 13136 16096 13142 16108
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 13136 16068 13369 16096
rect 13136 16056 13142 16068
rect 13357 16065 13369 16068
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16096 13599 16099
rect 14274 16096 14280 16108
rect 13587 16068 14280 16096
rect 13587 16065 13599 16068
rect 13541 16059 13599 16065
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 14458 16056 14464 16108
rect 14516 16096 14522 16108
rect 14642 16096 14648 16108
rect 14516 16068 14648 16096
rect 14516 16056 14522 16068
rect 14642 16056 14648 16068
rect 14700 16056 14706 16108
rect 15746 16096 15752 16108
rect 15707 16068 15752 16096
rect 15746 16056 15752 16068
rect 15804 16056 15810 16108
rect 16022 16096 16028 16108
rect 15983 16068 16028 16096
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 9950 15988 9956 16040
rect 10008 16028 10014 16040
rect 10045 16031 10103 16037
rect 10045 16028 10057 16031
rect 10008 16000 10057 16028
rect 10008 15988 10014 16000
rect 10045 15997 10057 16000
rect 10091 15997 10103 16031
rect 10045 15991 10103 15997
rect 11517 16031 11575 16037
rect 11517 15997 11529 16031
rect 11563 15997 11575 16031
rect 13630 16028 13636 16040
rect 13591 16000 13636 16028
rect 11517 15991 11575 15997
rect 9493 15963 9551 15969
rect 9493 15929 9505 15963
rect 9539 15929 9551 15963
rect 9493 15923 9551 15929
rect 9582 15920 9588 15972
rect 9640 15960 9646 15972
rect 11532 15960 11560 15991
rect 13630 15988 13636 16000
rect 13688 15988 13694 16040
rect 16868 16037 16896 16136
rect 17678 16124 17684 16136
rect 17736 16124 17742 16176
rect 17788 16164 17816 16204
rect 17862 16192 17868 16244
rect 17920 16232 17926 16244
rect 18509 16235 18567 16241
rect 18509 16232 18521 16235
rect 17920 16204 18521 16232
rect 17920 16192 17926 16204
rect 18509 16201 18521 16204
rect 18555 16201 18567 16235
rect 18509 16195 18567 16201
rect 18782 16192 18788 16244
rect 18840 16232 18846 16244
rect 18877 16235 18935 16241
rect 18877 16232 18889 16235
rect 18840 16204 18889 16232
rect 18840 16192 18846 16204
rect 18877 16201 18889 16204
rect 18923 16201 18935 16235
rect 18877 16195 18935 16201
rect 19797 16235 19855 16241
rect 19797 16201 19809 16235
rect 19843 16232 19855 16235
rect 20070 16232 20076 16244
rect 19843 16204 20076 16232
rect 19843 16201 19855 16204
rect 19797 16195 19855 16201
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 21450 16232 21456 16244
rect 21411 16204 21456 16232
rect 21450 16192 21456 16204
rect 21508 16192 21514 16244
rect 26237 16235 26295 16241
rect 26237 16201 26249 16235
rect 26283 16232 26295 16235
rect 26283 16204 27108 16232
rect 26283 16201 26295 16204
rect 26237 16195 26295 16201
rect 21082 16164 21088 16176
rect 17788 16136 21088 16164
rect 21082 16124 21088 16136
rect 21140 16124 21146 16176
rect 22002 16124 22008 16176
rect 22060 16164 22066 16176
rect 22934 16167 22992 16173
rect 22934 16164 22946 16167
rect 22060 16136 22946 16164
rect 22060 16124 22066 16136
rect 22934 16133 22946 16136
rect 22980 16133 22992 16167
rect 26878 16164 26884 16176
rect 22934 16127 22992 16133
rect 24044 16136 26884 16164
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16096 17095 16099
rect 17126 16096 17132 16108
rect 17083 16068 17132 16096
rect 17083 16065 17095 16068
rect 17037 16059 17095 16065
rect 17126 16056 17132 16068
rect 17184 16056 17190 16108
rect 17865 16099 17923 16105
rect 17865 16096 17877 16099
rect 17420 16068 17877 16096
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 16853 16031 16911 16037
rect 16853 15997 16865 16031
rect 16899 15997 16911 16031
rect 16853 15991 16911 15997
rect 9640 15932 11560 15960
rect 9640 15920 9646 15932
rect 14366 15920 14372 15972
rect 14424 15960 14430 15972
rect 14642 15960 14648 15972
rect 14424 15932 14648 15960
rect 14424 15920 14430 15932
rect 14642 15920 14648 15932
rect 14700 15960 14706 15972
rect 14936 15960 14964 15991
rect 17420 15969 17448 16068
rect 17865 16065 17877 16068
rect 17911 16065 17923 16099
rect 18417 16099 18475 16105
rect 18417 16096 18429 16099
rect 17865 16059 17923 16065
rect 17972 16068 18429 16096
rect 17678 16028 17684 16040
rect 17639 16000 17684 16028
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 14700 15932 14964 15960
rect 17405 15963 17463 15969
rect 14700 15920 14706 15932
rect 17405 15929 17417 15963
rect 17451 15929 17463 15963
rect 17405 15923 17463 15929
rect 17862 15920 17868 15972
rect 17920 15960 17926 15972
rect 17972 15960 18000 16068
rect 18417 16065 18429 16068
rect 18463 16065 18475 16099
rect 18417 16059 18475 16065
rect 19061 16099 19119 16105
rect 19061 16065 19073 16099
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 19076 16028 19104 16059
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19613 16099 19671 16105
rect 19613 16096 19625 16099
rect 19392 16068 19625 16096
rect 19392 16056 19398 16068
rect 19613 16065 19625 16068
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 20806 16096 20812 16108
rect 20767 16068 20812 16096
rect 20625 16059 20683 16065
rect 18095 16000 19104 16028
rect 19429 16031 19487 16037
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 19429 15997 19441 16031
rect 19475 16028 19487 16031
rect 19978 16028 19984 16040
rect 19475 16000 19984 16028
rect 19475 15997 19487 16000
rect 19429 15991 19487 15997
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 20640 16028 20668 16059
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21266 16096 21272 16108
rect 20956 16068 21001 16096
rect 21179 16068 21272 16096
rect 20956 16056 20962 16068
rect 21201 16028 21229 16068
rect 21266 16056 21272 16068
rect 21324 16056 21330 16108
rect 21453 16099 21511 16105
rect 21453 16065 21465 16099
rect 21499 16065 21511 16099
rect 23474 16096 23480 16108
rect 23435 16068 23480 16096
rect 21453 16059 21511 16065
rect 20640 16000 21229 16028
rect 17920 15932 18000 15960
rect 21468 15960 21496 16059
rect 23474 16056 23480 16068
rect 23532 16056 23538 16108
rect 23566 16056 23572 16108
rect 23624 16096 23630 16108
rect 23753 16099 23811 16105
rect 23624 16068 23669 16096
rect 23624 16056 23630 16068
rect 23753 16065 23765 16099
rect 23799 16096 23811 16099
rect 23842 16096 23848 16108
rect 23799 16068 23848 16096
rect 23799 16065 23811 16068
rect 23753 16059 23811 16065
rect 23842 16056 23848 16068
rect 23900 16056 23906 16108
rect 24044 16105 24072 16136
rect 26878 16124 26884 16136
rect 26936 16164 26942 16176
rect 27080 16164 27108 16204
rect 27218 16167 27276 16173
rect 27218 16164 27230 16167
rect 26936 16136 27016 16164
rect 27080 16136 27230 16164
rect 26936 16124 26942 16136
rect 24029 16099 24087 16105
rect 24029 16096 24041 16099
rect 23952 16068 24041 16096
rect 23201 16031 23259 16037
rect 23201 15997 23213 16031
rect 23247 16028 23259 16031
rect 23952 16028 23980 16068
rect 24029 16065 24041 16068
rect 24075 16065 24087 16099
rect 24285 16099 24343 16105
rect 24285 16096 24297 16099
rect 24029 16059 24087 16065
rect 24136 16068 24297 16096
rect 24136 16028 24164 16068
rect 24285 16065 24297 16068
rect 24331 16065 24343 16099
rect 25774 16096 25780 16108
rect 25735 16068 25780 16096
rect 24285 16059 24343 16065
rect 25774 16056 25780 16068
rect 25832 16056 25838 16108
rect 25869 16099 25927 16105
rect 25869 16065 25881 16099
rect 25915 16065 25927 16099
rect 25869 16059 25927 16065
rect 25961 16099 26019 16105
rect 25961 16065 25973 16099
rect 26007 16065 26019 16099
rect 26142 16096 26148 16108
rect 26103 16068 26148 16096
rect 25961 16059 26019 16065
rect 23247 16000 23980 16028
rect 24044 16000 24164 16028
rect 23247 15997 23259 16000
rect 23201 15991 23259 15997
rect 21821 15963 21879 15969
rect 21821 15960 21833 15963
rect 21468 15932 21833 15960
rect 17920 15920 17926 15932
rect 21821 15929 21833 15932
rect 21867 15960 21879 15963
rect 23753 15963 23811 15969
rect 21867 15932 22094 15960
rect 21867 15929 21879 15932
rect 21821 15923 21879 15929
rect 5442 15892 5448 15904
rect 5403 15864 5448 15892
rect 5442 15852 5448 15864
rect 5500 15852 5506 15904
rect 7742 15892 7748 15904
rect 7703 15864 7748 15892
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 9217 15895 9275 15901
rect 9217 15861 9229 15895
rect 9263 15892 9275 15895
rect 10134 15892 10140 15904
rect 9263 15864 10140 15892
rect 9263 15861 9275 15864
rect 9217 15855 9275 15861
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 10686 15892 10692 15904
rect 10647 15864 10692 15892
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 12250 15852 12256 15904
rect 12308 15892 12314 15904
rect 12986 15892 12992 15904
rect 12308 15864 12992 15892
rect 12308 15852 12314 15864
rect 12986 15852 12992 15864
rect 13044 15852 13050 15904
rect 13170 15892 13176 15904
rect 13131 15864 13176 15892
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 16942 15892 16948 15904
rect 15344 15864 16948 15892
rect 15344 15852 15350 15864
rect 16942 15852 16948 15864
rect 17000 15852 17006 15904
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 20073 15895 20131 15901
rect 20073 15892 20085 15895
rect 17368 15864 20085 15892
rect 17368 15852 17374 15864
rect 20073 15861 20085 15864
rect 20119 15861 20131 15895
rect 20438 15892 20444 15904
rect 20399 15864 20444 15892
rect 20073 15855 20131 15861
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 22066 15892 22094 15932
rect 23753 15929 23765 15963
rect 23799 15960 23811 15963
rect 24044 15960 24072 16000
rect 25406 15988 25412 16040
rect 25464 16028 25470 16040
rect 25884 16028 25912 16059
rect 25464 16000 25912 16028
rect 25976 16028 26004 16059
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 26234 16056 26240 16108
rect 26292 16096 26298 16108
rect 26988 16105 27016 16136
rect 27218 16133 27230 16136
rect 27264 16133 27276 16167
rect 27218 16127 27276 16133
rect 26973 16099 27031 16105
rect 26292 16068 26337 16096
rect 26292 16056 26298 16068
rect 26973 16065 26985 16099
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 26878 16028 26884 16040
rect 25976 16000 26884 16028
rect 25464 15988 25470 16000
rect 26878 15988 26884 16000
rect 26936 15988 26942 16040
rect 23799 15932 24072 15960
rect 23799 15929 23811 15932
rect 23753 15923 23811 15929
rect 22278 15892 22284 15904
rect 22066 15864 22284 15892
rect 22278 15852 22284 15864
rect 22336 15852 22342 15904
rect 25222 15852 25228 15904
rect 25280 15892 25286 15904
rect 25409 15895 25467 15901
rect 25409 15892 25421 15895
rect 25280 15864 25421 15892
rect 25280 15852 25286 15864
rect 25409 15861 25421 15864
rect 25455 15861 25467 15895
rect 28350 15892 28356 15904
rect 28311 15864 28356 15892
rect 25409 15855 25467 15861
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 1104 15802 28888 15824
rect 1104 15750 5582 15802
rect 5634 15750 5646 15802
rect 5698 15750 5710 15802
rect 5762 15750 5774 15802
rect 5826 15750 5838 15802
rect 5890 15750 14846 15802
rect 14898 15750 14910 15802
rect 14962 15750 14974 15802
rect 15026 15750 15038 15802
rect 15090 15750 15102 15802
rect 15154 15750 24110 15802
rect 24162 15750 24174 15802
rect 24226 15750 24238 15802
rect 24290 15750 24302 15802
rect 24354 15750 24366 15802
rect 24418 15750 28888 15802
rect 1104 15728 28888 15750
rect 11054 15688 11060 15700
rect 11015 15660 11060 15688
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 11790 15648 11796 15700
rect 11848 15688 11854 15700
rect 11977 15691 12035 15697
rect 11977 15688 11989 15691
rect 11848 15660 11989 15688
rect 11848 15648 11854 15660
rect 11977 15657 11989 15660
rect 12023 15657 12035 15691
rect 12434 15688 12440 15700
rect 11977 15651 12035 15657
rect 12189 15660 12440 15688
rect 5166 15552 5172 15564
rect 5127 15524 5172 15552
rect 5166 15512 5172 15524
rect 5224 15512 5230 15564
rect 8570 15552 8576 15564
rect 8531 15524 8576 15552
rect 8570 15512 8576 15524
rect 8628 15552 8634 15564
rect 9582 15552 9588 15564
rect 8628 15524 9588 15552
rect 8628 15512 8634 15524
rect 9582 15512 9588 15524
rect 9640 15552 9646 15564
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9640 15524 9689 15552
rect 9640 15512 9646 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9677 15515 9735 15521
rect 5442 15493 5448 15496
rect 5436 15484 5448 15493
rect 5403 15456 5448 15484
rect 5436 15447 5448 15456
rect 5442 15444 5448 15447
rect 5500 15444 5506 15496
rect 7742 15444 7748 15496
rect 7800 15484 7806 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 7800 15456 9137 15484
rect 7800 15444 7806 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 8328 15419 8386 15425
rect 8328 15385 8340 15419
rect 8374 15416 8386 15419
rect 9944 15419 10002 15425
rect 8374 15388 8984 15416
rect 8374 15385 8386 15388
rect 8328 15379 8386 15385
rect 6549 15351 6607 15357
rect 6549 15317 6561 15351
rect 6595 15348 6607 15351
rect 6822 15348 6828 15360
rect 6595 15320 6828 15348
rect 6595 15317 6607 15320
rect 6549 15311 6607 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 7190 15348 7196 15360
rect 7151 15320 7196 15348
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 8956 15357 8984 15388
rect 9944 15385 9956 15419
rect 9990 15416 10002 15419
rect 10042 15416 10048 15428
rect 9990 15388 10048 15416
rect 9990 15385 10002 15388
rect 9944 15379 10002 15385
rect 10042 15376 10048 15388
rect 10100 15376 10106 15428
rect 8941 15351 8999 15357
rect 8941 15317 8953 15351
rect 8987 15317 8999 15351
rect 11072 15348 11100 15648
rect 11698 15620 11704 15632
rect 11659 15592 11704 15620
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 12189 15552 12217 15660
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 13630 15648 13636 15700
rect 13688 15688 13694 15700
rect 15013 15691 15071 15697
rect 15013 15688 15025 15691
rect 13688 15660 15025 15688
rect 13688 15648 13694 15660
rect 15013 15657 15025 15660
rect 15059 15657 15071 15691
rect 15013 15651 15071 15657
rect 16025 15691 16083 15697
rect 16025 15657 16037 15691
rect 16071 15688 16083 15691
rect 16206 15688 16212 15700
rect 16071 15660 16212 15688
rect 16071 15657 16083 15660
rect 16025 15651 16083 15657
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 16761 15691 16819 15697
rect 16761 15657 16773 15691
rect 16807 15688 16819 15691
rect 17770 15688 17776 15700
rect 16807 15660 17776 15688
rect 16807 15657 16819 15660
rect 16761 15651 16819 15657
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 21634 15688 21640 15700
rect 21595 15660 21640 15688
rect 21634 15648 21640 15660
rect 21692 15648 21698 15700
rect 23566 15648 23572 15700
rect 23624 15688 23630 15700
rect 24397 15691 24455 15697
rect 24397 15688 24409 15691
rect 23624 15660 24409 15688
rect 23624 15648 23630 15660
rect 24397 15657 24409 15660
rect 24443 15657 24455 15691
rect 24854 15688 24860 15700
rect 24815 15660 24860 15688
rect 24397 15651 24455 15657
rect 24854 15648 24860 15660
rect 24912 15688 24918 15700
rect 25038 15688 25044 15700
rect 24912 15660 25044 15688
rect 24912 15648 24918 15660
rect 25038 15648 25044 15660
rect 25096 15648 25102 15700
rect 25498 15688 25504 15700
rect 25459 15660 25504 15688
rect 25498 15648 25504 15660
rect 25556 15688 25562 15700
rect 25556 15660 26648 15688
rect 25556 15648 25562 15660
rect 12250 15580 12256 15632
rect 12308 15620 12314 15632
rect 12802 15620 12808 15632
rect 12308 15592 12808 15620
rect 12308 15580 12314 15592
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 12986 15580 12992 15632
rect 13044 15620 13050 15632
rect 16393 15623 16451 15629
rect 16393 15620 16405 15623
rect 13044 15592 16405 15620
rect 13044 15580 13050 15592
rect 16393 15589 16405 15592
rect 16439 15589 16451 15623
rect 16850 15620 16856 15632
rect 16393 15583 16451 15589
rect 16500 15592 16856 15620
rect 13998 15552 14004 15564
rect 12189 15524 12388 15552
rect 11330 15484 11336 15496
rect 11291 15456 11336 15484
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 11422 15444 11428 15496
rect 11480 15484 11486 15496
rect 11517 15487 11575 15493
rect 11517 15484 11529 15487
rect 11480 15456 11529 15484
rect 11480 15444 11486 15456
rect 11517 15453 11529 15456
rect 11563 15453 11575 15487
rect 12250 15484 12256 15496
rect 12211 15456 12256 15484
rect 11517 15447 11575 15453
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 12360 15493 12388 15524
rect 12452 15524 14004 15552
rect 12452 15493 12480 15524
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 15194 15552 15200 15564
rect 14660 15524 15200 15552
rect 12345 15487 12403 15493
rect 12345 15453 12357 15487
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 12437 15487 12495 15493
rect 12437 15453 12449 15487
rect 12483 15453 12495 15487
rect 12437 15447 12495 15453
rect 12526 15444 12532 15496
rect 12584 15484 12590 15496
rect 12621 15487 12679 15493
rect 12621 15484 12633 15487
rect 12584 15456 12633 15484
rect 12584 15444 12590 15456
rect 12621 15453 12633 15456
rect 12667 15453 12679 15487
rect 13078 15484 13084 15496
rect 13039 15456 13084 15484
rect 12621 15447 12679 15453
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 13174 15487 13232 15493
rect 13174 15453 13186 15487
rect 13220 15453 13232 15487
rect 13446 15484 13452 15496
rect 13407 15456 13452 15484
rect 13174 15447 13232 15453
rect 13188 15416 13216 15447
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 13587 15487 13645 15493
rect 13587 15453 13599 15487
rect 13633 15484 13645 15487
rect 13722 15484 13728 15496
rect 13633 15456 13728 15484
rect 13633 15453 13645 15456
rect 13587 15447 13645 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14366 15484 14372 15496
rect 14327 15456 14372 15484
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 14458 15444 14464 15496
rect 14516 15484 14522 15496
rect 14660 15493 14688 15524
rect 15194 15512 15200 15524
rect 15252 15512 15258 15564
rect 15930 15552 15936 15564
rect 15843 15524 15936 15552
rect 14553 15487 14611 15493
rect 14553 15484 14565 15487
rect 14516 15456 14565 15484
rect 14516 15444 14522 15456
rect 14553 15453 14565 15456
rect 14599 15453 14611 15487
rect 14553 15447 14611 15453
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 15286 15484 15292 15496
rect 14783 15456 15292 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15856 15493 15884 15524
rect 15930 15512 15936 15524
rect 15988 15552 15994 15564
rect 16500 15552 16528 15592
rect 16850 15580 16856 15592
rect 16908 15580 16914 15632
rect 16942 15580 16948 15632
rect 17000 15620 17006 15632
rect 17000 15592 17632 15620
rect 17000 15580 17006 15592
rect 17221 15555 17279 15561
rect 17221 15552 17233 15555
rect 15988 15524 16528 15552
rect 16592 15524 17233 15552
rect 15988 15512 15994 15524
rect 16592 15496 16620 15524
rect 17221 15521 17233 15524
rect 17267 15521 17279 15555
rect 17221 15515 17279 15521
rect 15749 15487 15807 15493
rect 15749 15484 15761 15487
rect 15436 15456 15761 15484
rect 15436 15444 15442 15456
rect 15749 15453 15761 15456
rect 15795 15453 15807 15487
rect 15749 15447 15807 15453
rect 15841 15487 15899 15493
rect 15841 15453 15853 15487
rect 15887 15453 15899 15487
rect 16574 15484 16580 15496
rect 16487 15456 16580 15484
rect 15841 15447 15899 15453
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 16669 15487 16727 15493
rect 16669 15453 16681 15487
rect 16715 15484 16727 15487
rect 16715 15456 17264 15484
rect 16715 15453 16727 15456
rect 16669 15447 16727 15453
rect 17236 15428 17264 15456
rect 17310 15444 17316 15496
rect 17368 15484 17374 15496
rect 17604 15484 17632 15592
rect 17862 15512 17868 15564
rect 17920 15552 17926 15564
rect 18141 15555 18199 15561
rect 18141 15552 18153 15555
rect 17920 15524 18153 15552
rect 17920 15512 17926 15524
rect 18141 15521 18153 15524
rect 18187 15521 18199 15555
rect 19886 15552 19892 15564
rect 18141 15515 18199 15521
rect 18616 15524 19892 15552
rect 18049 15487 18107 15493
rect 18049 15484 18061 15487
rect 17368 15456 17461 15484
rect 17604 15456 18061 15484
rect 17368 15444 17374 15456
rect 18049 15453 18061 15456
rect 18095 15484 18107 15487
rect 18616 15484 18644 15524
rect 19886 15512 19892 15524
rect 19944 15512 19950 15564
rect 21266 15512 21272 15564
rect 21324 15552 21330 15564
rect 21726 15552 21732 15564
rect 21324 15524 21732 15552
rect 21324 15512 21330 15524
rect 21726 15512 21732 15524
rect 21784 15552 21790 15564
rect 24673 15555 24731 15561
rect 21784 15524 22140 15552
rect 21784 15512 21790 15524
rect 18782 15484 18788 15496
rect 18095 15456 18644 15484
rect 18743 15456 18788 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 18782 15444 18788 15456
rect 18840 15444 18846 15496
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19978 15484 19984 15496
rect 19939 15456 19984 15484
rect 19521 15447 19579 15453
rect 12406 15388 13216 15416
rect 13357 15419 13415 15425
rect 12406 15348 12434 15388
rect 13357 15385 13369 15419
rect 13403 15385 13415 15419
rect 13357 15379 13415 15385
rect 11072 15320 12434 15348
rect 8941 15311 8999 15317
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 13372 15348 13400 15379
rect 15194 15376 15200 15428
rect 15252 15416 15258 15428
rect 15473 15419 15531 15425
rect 15473 15416 15485 15419
rect 15252 15388 15485 15416
rect 15252 15376 15258 15388
rect 15473 15385 15485 15388
rect 15519 15385 15531 15419
rect 15473 15379 15531 15385
rect 15654 15376 15660 15428
rect 15712 15416 15718 15428
rect 16390 15416 16396 15428
rect 15712 15388 16396 15416
rect 15712 15376 15718 15388
rect 16390 15376 16396 15388
rect 16448 15376 16454 15428
rect 16850 15416 16856 15428
rect 16811 15388 16856 15416
rect 16850 15376 16856 15388
rect 16908 15376 16914 15428
rect 17218 15376 17224 15428
rect 17276 15376 17282 15428
rect 13446 15348 13452 15360
rect 12768 15320 13452 15348
rect 12768 15308 12774 15320
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 13538 15308 13544 15360
rect 13596 15348 13602 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13596 15320 13737 15348
rect 13596 15308 13602 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 16758 15308 16764 15360
rect 16816 15348 16822 15360
rect 17328 15348 17356 15444
rect 17402 15376 17408 15428
rect 17460 15416 17466 15428
rect 17954 15416 17960 15428
rect 17460 15388 17724 15416
rect 17915 15388 17960 15416
rect 17460 15376 17466 15388
rect 17586 15348 17592 15360
rect 16816 15320 17356 15348
rect 17547 15320 17592 15348
rect 16816 15308 16822 15320
rect 17586 15308 17592 15320
rect 17644 15308 17650 15360
rect 17696 15348 17724 15388
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 19536 15416 19564 15447
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 20990 15444 20996 15496
rect 21048 15484 21054 15496
rect 22112 15493 22140 15524
rect 24673 15521 24685 15555
rect 24719 15552 24731 15555
rect 25516 15552 25544 15648
rect 25869 15623 25927 15629
rect 25869 15589 25881 15623
rect 25915 15589 25927 15623
rect 25869 15583 25927 15589
rect 24719 15524 25544 15552
rect 25884 15552 25912 15583
rect 26142 15552 26148 15564
rect 25884 15524 26148 15552
rect 24719 15521 24731 15524
rect 24673 15515 24731 15521
rect 26142 15512 26148 15524
rect 26200 15552 26206 15564
rect 26421 15555 26479 15561
rect 26421 15552 26433 15555
rect 26200 15524 26433 15552
rect 26200 15512 26206 15524
rect 26421 15521 26433 15524
rect 26467 15521 26479 15555
rect 26421 15515 26479 15521
rect 21821 15487 21879 15493
rect 21821 15484 21833 15487
rect 21048 15456 21833 15484
rect 21048 15444 21054 15456
rect 21821 15453 21833 15456
rect 21867 15453 21879 15487
rect 21821 15447 21879 15453
rect 21913 15487 21971 15493
rect 21913 15453 21925 15487
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 22097 15487 22155 15493
rect 22097 15453 22109 15487
rect 22143 15453 22155 15487
rect 22097 15447 22155 15453
rect 22189 15487 22247 15493
rect 22189 15453 22201 15487
rect 22235 15484 22247 15487
rect 22278 15484 22284 15496
rect 22235 15456 22284 15484
rect 22235 15453 22247 15456
rect 22189 15447 22247 15453
rect 19886 15416 19892 15428
rect 18064 15388 19380 15416
rect 19536 15388 19892 15416
rect 18064 15348 18092 15388
rect 18598 15348 18604 15360
rect 17696 15320 18092 15348
rect 18559 15320 18604 15348
rect 18598 15308 18604 15320
rect 18656 15308 18662 15360
rect 19352 15357 19380 15388
rect 19886 15376 19892 15388
rect 19944 15376 19950 15428
rect 20254 15425 20260 15428
rect 20248 15379 20260 15425
rect 20312 15416 20318 15428
rect 20312 15388 20348 15416
rect 20254 15376 20260 15379
rect 20312 15376 20318 15388
rect 20806 15376 20812 15428
rect 20864 15416 20870 15428
rect 21928 15416 21956 15447
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 24946 15484 24952 15496
rect 24907 15456 24952 15484
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 25501 15487 25559 15493
rect 25501 15453 25513 15487
rect 25547 15453 25559 15487
rect 25501 15447 25559 15453
rect 25685 15487 25743 15493
rect 25685 15453 25697 15487
rect 25731 15453 25743 15487
rect 26510 15484 26516 15496
rect 26471 15456 26516 15484
rect 25685 15447 25743 15453
rect 22554 15416 22560 15428
rect 20864 15388 22560 15416
rect 20864 15376 20870 15388
rect 22554 15376 22560 15388
rect 22612 15376 22618 15428
rect 24854 15376 24860 15428
rect 24912 15416 24918 15428
rect 25516 15416 25544 15447
rect 25590 15416 25596 15428
rect 24912 15388 25596 15416
rect 24912 15376 24918 15388
rect 25590 15376 25596 15388
rect 25648 15376 25654 15428
rect 25700 15416 25728 15447
rect 26510 15444 26516 15456
rect 26568 15444 26574 15496
rect 26620 15484 26648 15660
rect 26878 15648 26884 15700
rect 26936 15688 26942 15700
rect 27341 15691 27399 15697
rect 27341 15688 27353 15691
rect 26936 15660 27353 15688
rect 26936 15648 26942 15660
rect 27341 15657 27353 15660
rect 27387 15657 27399 15691
rect 27341 15651 27399 15657
rect 26786 15580 26792 15632
rect 26844 15620 26850 15632
rect 27249 15623 27307 15629
rect 27249 15620 27261 15623
rect 26844 15592 27261 15620
rect 26844 15580 26850 15592
rect 27249 15589 27261 15592
rect 27295 15589 27307 15623
rect 27249 15583 27307 15589
rect 27433 15555 27491 15561
rect 27433 15521 27445 15555
rect 27479 15552 27491 15555
rect 28350 15552 28356 15564
rect 27479 15524 28356 15552
rect 27479 15521 27491 15524
rect 27433 15515 27491 15521
rect 27157 15487 27215 15493
rect 27157 15484 27169 15487
rect 26620 15456 27169 15484
rect 27157 15453 27169 15456
rect 27203 15453 27215 15487
rect 27157 15447 27215 15453
rect 26050 15416 26056 15428
rect 25700 15388 26056 15416
rect 26050 15376 26056 15388
rect 26108 15416 26114 15428
rect 27448 15416 27476 15515
rect 28350 15512 28356 15524
rect 28408 15512 28414 15564
rect 26108 15388 27476 15416
rect 26108 15376 26114 15388
rect 19337 15351 19395 15357
rect 19337 15317 19349 15351
rect 19383 15348 19395 15351
rect 20530 15348 20536 15360
rect 19383 15320 20536 15348
rect 19383 15317 19395 15320
rect 19337 15311 19395 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 21358 15348 21364 15360
rect 21319 15320 21364 15348
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 25608 15348 25636 15376
rect 26786 15348 26792 15360
rect 25608 15320 26792 15348
rect 26786 15308 26792 15320
rect 26844 15308 26850 15360
rect 26881 15351 26939 15357
rect 26881 15317 26893 15351
rect 26927 15348 26939 15351
rect 26970 15348 26976 15360
rect 26927 15320 26976 15348
rect 26927 15317 26939 15320
rect 26881 15311 26939 15317
rect 26970 15308 26976 15320
rect 27028 15308 27034 15360
rect 28258 15348 28264 15360
rect 28219 15320 28264 15348
rect 28258 15308 28264 15320
rect 28316 15308 28322 15360
rect 1104 15258 28888 15280
rect 1104 15206 10214 15258
rect 10266 15206 10278 15258
rect 10330 15206 10342 15258
rect 10394 15206 10406 15258
rect 10458 15206 10470 15258
rect 10522 15206 19478 15258
rect 19530 15206 19542 15258
rect 19594 15206 19606 15258
rect 19658 15206 19670 15258
rect 19722 15206 19734 15258
rect 19786 15206 28888 15258
rect 1104 15184 28888 15206
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 10686 15144 10692 15156
rect 4120 15116 10692 15144
rect 4120 15104 4126 15116
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 11149 15147 11207 15153
rect 11149 15113 11161 15147
rect 11195 15144 11207 15147
rect 12250 15144 12256 15156
rect 11195 15116 12256 15144
rect 11195 15113 11207 15116
rect 11149 15107 11207 15113
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 13722 15104 13728 15156
rect 13780 15104 13786 15156
rect 14001 15147 14059 15153
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 14366 15144 14372 15156
rect 14047 15116 14372 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 14366 15104 14372 15116
rect 14424 15104 14430 15156
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 14792 15116 14933 15144
rect 14792 15104 14798 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 15473 15147 15531 15153
rect 15473 15113 15485 15147
rect 15519 15144 15531 15147
rect 15654 15144 15660 15156
rect 15519 15116 15660 15144
rect 15519 15113 15531 15116
rect 15473 15107 15531 15113
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 16666 15104 16672 15156
rect 16724 15144 16730 15156
rect 17221 15147 17279 15153
rect 17221 15144 17233 15147
rect 16724 15116 17233 15144
rect 16724 15104 16730 15116
rect 17221 15113 17233 15116
rect 17267 15144 17279 15147
rect 17862 15144 17868 15156
rect 17267 15116 17868 15144
rect 17267 15113 17279 15116
rect 17221 15107 17279 15113
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 19886 15144 19892 15156
rect 18156 15116 19892 15144
rect 5537 15079 5595 15085
rect 5537 15045 5549 15079
rect 5583 15076 5595 15079
rect 5902 15076 5908 15088
rect 5583 15048 5908 15076
rect 5583 15045 5595 15048
rect 5537 15039 5595 15045
rect 5902 15036 5908 15048
rect 5960 15036 5966 15088
rect 7190 15036 7196 15088
rect 7248 15076 7254 15088
rect 7929 15079 7987 15085
rect 7929 15076 7941 15079
rect 7248 15048 7941 15076
rect 7248 15036 7254 15048
rect 7929 15045 7941 15048
rect 7975 15076 7987 15079
rect 7975 15048 12572 15076
rect 7975 15045 7987 15048
rect 7929 15039 7987 15045
rect 5721 15011 5779 15017
rect 5721 14977 5733 15011
rect 5767 15008 5779 15011
rect 6733 15011 6791 15017
rect 5767 14980 6408 15008
rect 5767 14977 5779 14980
rect 5721 14971 5779 14977
rect 5261 14943 5319 14949
rect 5261 14909 5273 14943
rect 5307 14940 5319 14943
rect 5902 14940 5908 14952
rect 5307 14912 5908 14940
rect 5307 14909 5319 14912
rect 5261 14903 5319 14909
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 6380 14881 6408 14980
rect 6733 14977 6745 15011
rect 6779 15008 6791 15011
rect 7098 15008 7104 15020
rect 6779 14980 7104 15008
rect 6779 14977 6791 14980
rect 6733 14971 6791 14977
rect 7098 14968 7104 14980
rect 7156 15008 7162 15020
rect 8021 15011 8079 15017
rect 8021 15008 8033 15011
rect 7156 14980 8033 15008
rect 7156 14968 7162 14980
rect 8021 14977 8033 14980
rect 8067 14977 8079 15011
rect 9398 15008 9404 15020
rect 9359 14980 9404 15008
rect 8021 14971 8079 14977
rect 9398 14968 9404 14980
rect 9456 14968 9462 15020
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 9953 15011 10011 15017
rect 9953 15008 9965 15011
rect 9631 14980 9965 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 9953 14977 9965 14980
rect 9999 14977 10011 15011
rect 9953 14971 10011 14977
rect 10134 14968 10140 15020
rect 10192 15008 10198 15020
rect 10597 15011 10655 15017
rect 10597 15008 10609 15011
rect 10192 14980 10609 15008
rect 10192 14968 10198 14980
rect 10597 14977 10609 14980
rect 10643 14977 10655 15011
rect 12066 15008 12072 15020
rect 12027 14980 12072 15008
rect 10597 14971 10655 14977
rect 12066 14968 12072 14980
rect 12124 14968 12130 15020
rect 12544 15017 12572 15048
rect 12618 15036 12624 15088
rect 12676 15076 12682 15088
rect 12805 15079 12863 15085
rect 12805 15076 12817 15079
rect 12676 15048 12817 15076
rect 12676 15036 12682 15048
rect 12805 15045 12817 15048
rect 12851 15045 12863 15079
rect 13740 15076 13768 15104
rect 15933 15079 15991 15085
rect 12805 15039 12863 15045
rect 12917 15048 14785 15076
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12530 15011 12588 15017
rect 12530 14977 12542 15011
rect 12576 14977 12588 15011
rect 12710 15008 12716 15020
rect 12671 14980 12716 15008
rect 12530 14971 12588 14977
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14909 6975 14943
rect 8202 14940 8208 14952
rect 8163 14912 8208 14940
rect 6917 14903 6975 14909
rect 6365 14875 6423 14881
rect 6365 14841 6377 14875
rect 6411 14841 6423 14875
rect 6365 14835 6423 14841
rect 6730 14832 6736 14884
rect 6788 14872 6794 14884
rect 6932 14872 6960 14903
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 9214 14940 9220 14952
rect 9175 14912 9220 14940
rect 9214 14900 9220 14912
rect 9272 14900 9278 14952
rect 11790 14900 11796 14952
rect 11848 14940 11854 14952
rect 12342 14940 12348 14952
rect 11848 14912 12348 14940
rect 11848 14900 11854 14912
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 12452 14940 12480 14971
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 12917 15017 12945 15048
rect 12902 15011 12960 15017
rect 12902 14977 12914 15011
rect 12948 14977 12960 15011
rect 12902 14971 12960 14977
rect 13078 14968 13084 15020
rect 13136 15008 13142 15020
rect 13354 15008 13360 15020
rect 13136 14980 13360 15008
rect 13136 14968 13142 14980
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 13630 15008 13636 15020
rect 13504 14980 13549 15008
rect 13591 14980 13636 15008
rect 13504 14968 13510 14980
rect 13630 14968 13636 14980
rect 13688 14968 13694 15020
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 14977 13783 15011
rect 13725 14971 13783 14977
rect 13096 14940 13124 14968
rect 12452 14912 13124 14940
rect 13740 14940 13768 14971
rect 13814 14968 13820 15020
rect 13872 15017 13878 15020
rect 13872 15008 13880 15017
rect 13872 14980 13917 15008
rect 13872 14971 13880 14980
rect 13872 14968 13878 14971
rect 14182 14968 14188 15020
rect 14240 15008 14246 15020
rect 14277 15011 14335 15017
rect 14277 15008 14289 15011
rect 14240 14980 14289 15008
rect 14240 14968 14246 14980
rect 14277 14977 14289 14980
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14757 15017 14785 15048
rect 15933 15045 15945 15079
rect 15979 15076 15991 15079
rect 15979 15048 17724 15076
rect 15979 15045 15991 15048
rect 15933 15039 15991 15045
rect 14553 15011 14611 15017
rect 14424 14980 14469 15008
rect 14424 14968 14430 14980
rect 14553 14977 14565 15011
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 14645 15011 14703 15017
rect 14645 14977 14657 15011
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 14742 15011 14800 15017
rect 14742 14977 14754 15011
rect 14788 14977 14800 15011
rect 14742 14971 14800 14977
rect 13998 14940 14004 14952
rect 13740 14912 14004 14940
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 14568 14940 14596 14971
rect 14200 14912 14596 14940
rect 7558 14872 7564 14884
rect 6788 14844 6960 14872
rect 7519 14844 7564 14872
rect 6788 14832 6794 14844
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 10042 14832 10048 14884
rect 10100 14872 10106 14884
rect 10413 14875 10471 14881
rect 10413 14872 10425 14875
rect 10100 14844 10425 14872
rect 10100 14832 10106 14844
rect 10413 14841 10425 14844
rect 10459 14841 10471 14875
rect 10413 14835 10471 14841
rect 11609 14875 11667 14881
rect 11609 14841 11621 14875
rect 11655 14872 11667 14875
rect 13078 14872 13084 14884
rect 11655 14844 12434 14872
rect 13039 14844 13084 14872
rect 11655 14841 11667 14844
rect 11609 14835 11667 14841
rect 10134 14804 10140 14816
rect 10095 14776 10140 14804
rect 10134 14764 10140 14776
rect 10192 14764 10198 14816
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 11977 14807 12035 14813
rect 11977 14804 11989 14807
rect 11848 14776 11989 14804
rect 11848 14764 11854 14776
rect 11977 14773 11989 14776
rect 12023 14773 12035 14807
rect 12406 14804 12434 14844
rect 13078 14832 13084 14844
rect 13136 14832 13142 14884
rect 12894 14804 12900 14816
rect 12406 14776 12900 14804
rect 11977 14767 12035 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 13630 14764 13636 14816
rect 13688 14804 13694 14816
rect 14200 14804 14228 14912
rect 14660 14872 14688 14971
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 15252 14980 16681 15008
rect 15252 14968 15258 14980
rect 16669 14977 16681 14980
rect 16715 15008 16727 15011
rect 16758 15008 16764 15020
rect 16715 14980 16764 15008
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 16758 14968 16764 14980
rect 16816 14968 16822 15020
rect 17034 15008 17040 15020
rect 16995 14980 17040 15008
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 17589 15011 17647 15017
rect 17589 15008 17601 15011
rect 17368 14980 17601 15008
rect 17368 14968 17374 14980
rect 17589 14977 17601 14980
rect 17635 14977 17647 15011
rect 17589 14971 17647 14977
rect 15378 14940 15384 14952
rect 15339 14912 15384 14940
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 17497 14943 17555 14949
rect 17497 14909 17509 14943
rect 17543 14940 17555 14943
rect 17696 14940 17724 15048
rect 17770 14940 17776 14952
rect 17543 14912 17776 14940
rect 17543 14909 17555 14912
rect 17497 14903 17555 14909
rect 17770 14900 17776 14912
rect 17828 14900 17834 14952
rect 14292 14844 14688 14872
rect 15933 14875 15991 14881
rect 14292 14816 14320 14844
rect 15933 14841 15945 14875
rect 15979 14872 15991 14875
rect 16574 14872 16580 14884
rect 15979 14844 16580 14872
rect 15979 14841 15991 14844
rect 15933 14835 15991 14841
rect 16574 14832 16580 14844
rect 16632 14832 16638 14884
rect 13688 14776 14228 14804
rect 13688 14764 13694 14776
rect 14274 14764 14280 14816
rect 14332 14764 14338 14816
rect 14366 14764 14372 14816
rect 14424 14804 14430 14816
rect 15197 14807 15255 14813
rect 15197 14804 15209 14807
rect 14424 14776 15209 14804
rect 14424 14764 14430 14776
rect 15197 14773 15209 14776
rect 15243 14773 15255 14807
rect 15197 14767 15255 14773
rect 15286 14764 15292 14816
rect 15344 14804 15350 14816
rect 18156 14804 18184 15116
rect 19886 15104 19892 15116
rect 19944 15104 19950 15156
rect 20349 15147 20407 15153
rect 20349 15113 20361 15147
rect 20395 15144 20407 15147
rect 21269 15147 21327 15153
rect 21269 15144 21281 15147
rect 20395 15116 21281 15144
rect 20395 15113 20407 15116
rect 20349 15107 20407 15113
rect 21269 15113 21281 15116
rect 21315 15113 21327 15147
rect 21269 15107 21327 15113
rect 21726 15104 21732 15156
rect 21784 15144 21790 15156
rect 21821 15147 21879 15153
rect 21821 15144 21833 15147
rect 21784 15116 21833 15144
rect 21784 15104 21790 15116
rect 21821 15113 21833 15116
rect 21867 15113 21879 15147
rect 22554 15144 22560 15156
rect 22515 15116 22560 15144
rect 21821 15107 21879 15113
rect 22554 15104 22560 15116
rect 22612 15104 22618 15156
rect 19978 15076 19984 15088
rect 18340 15048 19984 15076
rect 18340 14952 18368 15048
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 20165 15079 20223 15085
rect 20165 15045 20177 15079
rect 20211 15076 20223 15079
rect 20622 15076 20628 15088
rect 20211 15048 20628 15076
rect 20211 15045 20223 15048
rect 20165 15039 20223 15045
rect 20364 15020 20392 15048
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 21358 15076 21364 15088
rect 21271 15048 21364 15076
rect 18598 15017 18604 15020
rect 18592 15008 18604 15017
rect 18559 14980 18604 15008
rect 18592 14971 18604 14980
rect 18598 14968 18604 14971
rect 18656 14968 18662 15020
rect 20346 14968 20352 15020
rect 20404 14968 20410 15020
rect 20438 14968 20444 15020
rect 20496 15008 20502 15020
rect 21284 15017 21312 15048
rect 21358 15036 21364 15048
rect 21416 15076 21422 15088
rect 21416 15048 21772 15076
rect 21416 15036 21422 15048
rect 21744 15020 21772 15048
rect 22094 15036 22100 15088
rect 22152 15076 22158 15088
rect 26786 15076 26792 15088
rect 22152 15048 22692 15076
rect 22152 15036 22158 15048
rect 21269 15011 21327 15017
rect 20496 14980 20541 15008
rect 20496 14968 20502 14980
rect 21269 14977 21281 15011
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 21453 15011 21511 15017
rect 21453 14977 21465 15011
rect 21499 14977 21511 15011
rect 21453 14971 21511 14977
rect 18322 14940 18328 14952
rect 18283 14912 18328 14940
rect 18322 14900 18328 14912
rect 18380 14900 18386 14952
rect 19702 14900 19708 14952
rect 19760 14940 19766 14952
rect 20070 14940 20076 14952
rect 19760 14912 20076 14940
rect 19760 14900 19766 14912
rect 20070 14900 20076 14912
rect 20128 14900 20134 14952
rect 21468 14940 21496 14971
rect 21726 14968 21732 15020
rect 21784 15008 21790 15020
rect 22664 15017 22692 15048
rect 22940 15048 26792 15076
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21784 14980 22017 15008
rect 21784 14968 21790 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22189 15011 22247 15017
rect 22189 14977 22201 15011
rect 22235 15008 22247 15011
rect 22649 15011 22707 15017
rect 22235 14980 22269 15008
rect 22235 14977 22247 14980
rect 22189 14971 22247 14977
rect 22649 14977 22661 15011
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 22204 14940 22232 14971
rect 22554 14940 22560 14952
rect 21468 14912 22560 14940
rect 22554 14900 22560 14912
rect 22612 14900 22618 14952
rect 20165 14875 20223 14881
rect 19260 14844 19840 14872
rect 15344 14776 18184 14804
rect 15344 14764 15350 14776
rect 18506 14764 18512 14816
rect 18564 14804 18570 14816
rect 19260 14804 19288 14844
rect 19702 14804 19708 14816
rect 18564 14776 19288 14804
rect 19663 14776 19708 14804
rect 18564 14764 18570 14776
rect 19702 14764 19708 14776
rect 19760 14764 19766 14816
rect 19812 14804 19840 14844
rect 20165 14841 20177 14875
rect 20211 14872 20223 14875
rect 20254 14872 20260 14884
rect 20211 14844 20260 14872
rect 20211 14841 20223 14844
rect 20165 14835 20223 14841
rect 20254 14832 20260 14844
rect 20312 14832 20318 14884
rect 20530 14832 20536 14884
rect 20588 14872 20594 14884
rect 22940 14872 22968 15048
rect 26786 15036 26792 15048
rect 26844 15036 26850 15088
rect 23273 15011 23331 15017
rect 23273 14977 23285 15011
rect 23319 15008 23331 15011
rect 23658 15008 23664 15020
rect 23319 14980 23664 15008
rect 23319 14977 23331 14980
rect 23273 14971 23331 14977
rect 23658 14968 23664 14980
rect 23716 14968 23722 15020
rect 24673 15011 24731 15017
rect 24673 15008 24685 15011
rect 24412 14980 24685 15008
rect 23017 14943 23075 14949
rect 23017 14909 23029 14943
rect 23063 14909 23075 14943
rect 23017 14903 23075 14909
rect 20588 14844 21036 14872
rect 20588 14832 20594 14844
rect 20809 14807 20867 14813
rect 20809 14804 20821 14807
rect 19812 14776 20821 14804
rect 20809 14773 20821 14776
rect 20855 14804 20867 14807
rect 20898 14804 20904 14816
rect 20855 14776 20904 14804
rect 20855 14773 20867 14776
rect 20809 14767 20867 14773
rect 20898 14764 20904 14776
rect 20956 14764 20962 14816
rect 21008 14804 21036 14844
rect 22066 14844 22968 14872
rect 22066 14804 22094 14844
rect 21008 14776 22094 14804
rect 23032 14804 23060 14903
rect 23382 14804 23388 14816
rect 23032 14776 23388 14804
rect 23382 14764 23388 14776
rect 23440 14764 23446 14816
rect 24026 14764 24032 14816
rect 24084 14804 24090 14816
rect 24412 14813 24440 14980
rect 24673 14977 24685 14980
rect 24719 14977 24731 15011
rect 24673 14971 24731 14977
rect 24857 15011 24915 15017
rect 24857 14977 24869 15011
rect 24903 15008 24915 15011
rect 26050 15008 26056 15020
rect 24903 14980 26056 15008
rect 24903 14977 24915 14980
rect 24857 14971 24915 14977
rect 26050 14968 26056 14980
rect 26108 14968 26114 15020
rect 27246 15017 27252 15020
rect 27240 14971 27252 15017
rect 27304 15008 27310 15020
rect 27304 14980 27340 15008
rect 27246 14968 27252 14971
rect 27304 14968 27310 14980
rect 25317 14943 25375 14949
rect 25317 14909 25329 14943
rect 25363 14909 25375 14943
rect 25590 14940 25596 14952
rect 25551 14912 25596 14940
rect 25317 14903 25375 14909
rect 25222 14872 25228 14884
rect 24872 14844 25228 14872
rect 24872 14813 24900 14844
rect 25222 14832 25228 14844
rect 25280 14832 25286 14884
rect 25332 14872 25360 14903
rect 25590 14900 25596 14912
rect 25648 14900 25654 14952
rect 26142 14900 26148 14952
rect 26200 14940 26206 14952
rect 26973 14943 27031 14949
rect 26973 14940 26985 14943
rect 26200 14912 26985 14940
rect 26200 14900 26206 14912
rect 26973 14909 26985 14912
rect 27019 14909 27031 14943
rect 26973 14903 27031 14909
rect 25866 14872 25872 14884
rect 25332 14844 25872 14872
rect 25866 14832 25872 14844
rect 25924 14832 25930 14884
rect 24397 14807 24455 14813
rect 24397 14804 24409 14807
rect 24084 14776 24409 14804
rect 24084 14764 24090 14776
rect 24397 14773 24409 14776
rect 24443 14773 24455 14807
rect 24397 14767 24455 14773
rect 24857 14807 24915 14813
rect 24857 14773 24869 14807
rect 24903 14773 24915 14807
rect 25038 14804 25044 14816
rect 24999 14776 25044 14804
rect 24857 14767 24915 14773
rect 25038 14764 25044 14776
rect 25096 14764 25102 14816
rect 28350 14804 28356 14816
rect 28311 14776 28356 14804
rect 28350 14764 28356 14776
rect 28408 14764 28414 14816
rect 1104 14714 28888 14736
rect 1104 14662 5582 14714
rect 5634 14662 5646 14714
rect 5698 14662 5710 14714
rect 5762 14662 5774 14714
rect 5826 14662 5838 14714
rect 5890 14662 14846 14714
rect 14898 14662 14910 14714
rect 14962 14662 14974 14714
rect 15026 14662 15038 14714
rect 15090 14662 15102 14714
rect 15154 14662 24110 14714
rect 24162 14662 24174 14714
rect 24226 14662 24238 14714
rect 24290 14662 24302 14714
rect 24354 14662 24366 14714
rect 24418 14662 28888 14714
rect 1104 14640 28888 14662
rect 11606 14560 11612 14612
rect 11664 14600 11670 14612
rect 13446 14600 13452 14612
rect 11664 14572 13452 14600
rect 11664 14560 11670 14572
rect 13446 14560 13452 14572
rect 13504 14560 13510 14612
rect 16393 14603 16451 14609
rect 16393 14569 16405 14603
rect 16439 14600 16451 14603
rect 17218 14600 17224 14612
rect 16439 14572 17224 14600
rect 16439 14569 16451 14572
rect 16393 14563 16451 14569
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 18233 14603 18291 14609
rect 18233 14569 18245 14603
rect 18279 14600 18291 14603
rect 18782 14600 18788 14612
rect 18279 14572 18788 14600
rect 18279 14569 18291 14572
rect 18233 14563 18291 14569
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 24026 14600 24032 14612
rect 22848 14572 24032 14600
rect 12158 14532 12164 14544
rect 11992 14504 12164 14532
rect 7377 14467 7435 14473
rect 7377 14433 7389 14467
rect 7423 14464 7435 14467
rect 9214 14464 9220 14476
rect 7423 14436 9220 14464
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 9214 14424 9220 14436
rect 9272 14464 9278 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9272 14436 9689 14464
rect 9272 14424 9278 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 9766 14424 9772 14476
rect 9824 14464 9830 14476
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 9824 14436 10241 14464
rect 9824 14424 9830 14436
rect 10229 14433 10241 14436
rect 10275 14433 10287 14467
rect 10229 14427 10287 14433
rect 7558 14396 7564 14408
rect 7519 14368 7564 14396
rect 7558 14356 7564 14368
rect 7616 14356 7622 14408
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14396 7803 14399
rect 8205 14399 8263 14405
rect 8205 14396 8217 14399
rect 7791 14368 8217 14396
rect 7791 14365 7803 14368
rect 7745 14359 7803 14365
rect 8205 14365 8217 14368
rect 8251 14365 8263 14399
rect 9950 14396 9956 14408
rect 9911 14368 9956 14396
rect 8205 14359 8263 14365
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 10134 14356 10140 14408
rect 10192 14396 10198 14408
rect 10485 14399 10543 14405
rect 10485 14396 10497 14399
rect 10192 14368 10497 14396
rect 10192 14356 10198 14368
rect 10485 14365 10497 14368
rect 10531 14365 10543 14399
rect 11992 14396 12020 14504
rect 12158 14492 12164 14504
rect 12216 14532 12222 14544
rect 13265 14535 13323 14541
rect 13265 14532 13277 14535
rect 12216 14504 13277 14532
rect 12216 14492 12222 14504
rect 13265 14501 13277 14504
rect 13311 14532 13323 14535
rect 13814 14532 13820 14544
rect 13311 14504 13820 14532
rect 13311 14501 13323 14504
rect 13265 14495 13323 14501
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 15286 14532 15292 14544
rect 14113 14504 15292 14532
rect 12066 14424 12072 14476
rect 12124 14464 12130 14476
rect 12437 14467 12495 14473
rect 12437 14464 12449 14467
rect 12124 14436 12449 14464
rect 12124 14424 12130 14436
rect 12437 14433 12449 14436
rect 12483 14464 12495 14467
rect 14113 14464 14141 14504
rect 15286 14492 15292 14504
rect 15344 14492 15350 14544
rect 15378 14492 15384 14544
rect 15436 14532 15442 14544
rect 16945 14535 17003 14541
rect 16945 14532 16957 14535
rect 15436 14504 16957 14532
rect 15436 14492 15442 14504
rect 16945 14501 16957 14504
rect 16991 14501 17003 14535
rect 16945 14495 17003 14501
rect 18414 14492 18420 14544
rect 18472 14532 18478 14544
rect 19150 14532 19156 14544
rect 18472 14504 19156 14532
rect 18472 14492 18478 14504
rect 19150 14492 19156 14504
rect 19208 14532 19214 14544
rect 20349 14535 20407 14541
rect 19208 14504 19555 14532
rect 19208 14492 19214 14504
rect 12483 14436 14141 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 14182 14424 14188 14476
rect 14240 14464 14246 14476
rect 14369 14467 14427 14473
rect 14369 14464 14381 14467
rect 14240 14436 14381 14464
rect 14240 14424 14246 14436
rect 14369 14433 14381 14436
rect 14415 14433 14427 14467
rect 14369 14427 14427 14433
rect 14458 14424 14464 14476
rect 14516 14464 14522 14476
rect 16114 14464 16120 14476
rect 14516 14436 16120 14464
rect 14516 14424 14522 14436
rect 12161 14399 12219 14405
rect 12161 14396 12173 14399
rect 11992 14368 12173 14396
rect 10485 14359 10543 14365
rect 12161 14365 12173 14368
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 13354 14356 13360 14408
rect 13412 14396 13418 14408
rect 14090 14396 14096 14408
rect 13412 14368 13584 14396
rect 14051 14368 14096 14396
rect 13412 14356 13418 14368
rect 9306 14288 9312 14340
rect 9364 14328 9370 14340
rect 9364 14300 12434 14328
rect 9364 14288 9370 14300
rect 5902 14220 5908 14272
rect 5960 14260 5966 14272
rect 6089 14263 6147 14269
rect 6089 14260 6101 14263
rect 5960 14232 6101 14260
rect 5960 14220 5966 14232
rect 6089 14229 6101 14232
rect 6135 14260 6147 14263
rect 6546 14260 6552 14272
rect 6135 14232 6552 14260
rect 6135 14229 6147 14232
rect 6089 14223 6147 14229
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 8018 14260 8024 14272
rect 7979 14232 8024 14260
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 11606 14260 11612 14272
rect 11567 14232 11612 14260
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 12406 14260 12434 14300
rect 12894 14288 12900 14340
rect 12952 14328 12958 14340
rect 13446 14328 13452 14340
rect 12952 14300 13308 14328
rect 13407 14300 13452 14328
rect 12952 14288 12958 14300
rect 13078 14260 13084 14272
rect 12406 14232 13084 14260
rect 13078 14220 13084 14232
rect 13136 14220 13142 14272
rect 13280 14260 13308 14300
rect 13446 14288 13452 14300
rect 13504 14288 13510 14340
rect 13556 14328 13584 14368
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 14200 14328 14228 14424
rect 15194 14396 15200 14408
rect 13556 14300 14228 14328
rect 14568 14368 15200 14396
rect 14568 14260 14596 14368
rect 15194 14356 15200 14368
rect 15252 14356 15258 14408
rect 15488 14405 15516 14436
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 16574 14464 16580 14476
rect 16316 14436 16580 14464
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14365 15531 14399
rect 15930 14396 15936 14408
rect 15891 14368 15936 14396
rect 15473 14359 15531 14365
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16316 14405 16344 14436
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 18601 14467 18659 14473
rect 18601 14464 18613 14467
rect 16960 14436 18613 14464
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14365 16359 14399
rect 16301 14359 16359 14365
rect 16485 14399 16543 14405
rect 16485 14365 16497 14399
rect 16531 14396 16543 14399
rect 16850 14396 16856 14408
rect 16531 14368 16856 14396
rect 16531 14365 16543 14368
rect 16485 14359 16543 14365
rect 16850 14356 16856 14368
rect 16908 14396 16914 14408
rect 16960 14396 16988 14436
rect 18601 14433 18613 14436
rect 18647 14433 18659 14467
rect 18601 14427 18659 14433
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 19392 14436 19472 14464
rect 19392 14424 19398 14436
rect 17221 14399 17279 14405
rect 16908 14368 16988 14396
rect 17126 14393 17184 14399
rect 17126 14390 17138 14393
rect 16908 14356 16914 14368
rect 17052 14362 17138 14390
rect 14642 14288 14648 14340
rect 14700 14328 14706 14340
rect 14700 14300 16160 14328
rect 14700 14288 14706 14300
rect 15286 14260 15292 14272
rect 13280 14232 14596 14260
rect 15247 14232 15292 14260
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 16132 14269 16160 14300
rect 16117 14263 16175 14269
rect 16117 14229 16129 14263
rect 16163 14229 16175 14263
rect 17052 14260 17080 14362
rect 17126 14359 17138 14362
rect 17172 14359 17184 14393
rect 17221 14365 17233 14399
rect 17267 14396 17279 14399
rect 17328 14396 17417 14398
rect 17267 14370 17540 14396
rect 17267 14368 17356 14370
rect 17389 14368 17540 14370
rect 17267 14365 17279 14368
rect 17221 14359 17279 14365
rect 17126 14353 17184 14359
rect 17512 14340 17540 14368
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 17865 14399 17923 14405
rect 17865 14396 17877 14399
rect 17644 14368 17877 14396
rect 17644 14356 17650 14368
rect 17865 14365 17877 14368
rect 17911 14365 17923 14399
rect 18506 14396 18512 14408
rect 17865 14359 17923 14365
rect 17972 14368 18512 14396
rect 17494 14288 17500 14340
rect 17552 14328 17558 14340
rect 17972 14328 18000 14368
rect 18506 14356 18512 14368
rect 18564 14356 18570 14408
rect 18690 14396 18696 14408
rect 18651 14368 18696 14396
rect 18690 14356 18696 14368
rect 18748 14356 18754 14408
rect 19444 14405 19472 14436
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 17552 14300 18000 14328
rect 18049 14331 18107 14337
rect 17552 14288 17558 14300
rect 18049 14297 18061 14331
rect 18095 14328 18107 14331
rect 19334 14328 19340 14340
rect 18095 14300 19340 14328
rect 18095 14297 18107 14300
rect 18049 14291 18107 14297
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 19527 14328 19555 14504
rect 20349 14501 20361 14535
rect 20395 14532 20407 14535
rect 21910 14532 21916 14544
rect 20395 14504 21916 14532
rect 20395 14501 20407 14504
rect 20349 14495 20407 14501
rect 21910 14492 21916 14504
rect 21968 14492 21974 14544
rect 22848 14473 22876 14572
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 25130 14560 25136 14612
rect 25188 14560 25194 14612
rect 25317 14603 25375 14609
rect 25317 14569 25329 14603
rect 25363 14569 25375 14603
rect 26050 14600 26056 14612
rect 26011 14572 26056 14600
rect 25317 14563 25375 14569
rect 23658 14492 23664 14544
rect 23716 14532 23722 14544
rect 23937 14535 23995 14541
rect 23716 14504 23761 14532
rect 23716 14492 23722 14504
rect 23937 14501 23949 14535
rect 23983 14532 23995 14535
rect 25148 14532 25176 14560
rect 23983 14504 25176 14532
rect 25332 14532 25360 14563
rect 26050 14560 26056 14572
rect 26108 14560 26114 14612
rect 27246 14560 27252 14612
rect 27304 14600 27310 14612
rect 27433 14603 27491 14609
rect 27433 14600 27445 14603
rect 27304 14572 27445 14600
rect 27304 14560 27310 14572
rect 27433 14569 27445 14572
rect 27479 14569 27491 14603
rect 27433 14563 27491 14569
rect 25332 14504 27261 14532
rect 23983 14501 23995 14504
rect 23937 14495 23995 14501
rect 19613 14467 19671 14473
rect 19613 14433 19625 14467
rect 19659 14464 19671 14467
rect 21545 14467 21603 14473
rect 21545 14464 21557 14467
rect 19659 14436 21557 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 21545 14433 21557 14436
rect 21591 14433 21603 14467
rect 22833 14467 22891 14473
rect 21545 14427 21603 14433
rect 21652 14436 22787 14464
rect 19705 14399 19763 14405
rect 19705 14365 19717 14399
rect 19751 14396 19763 14399
rect 19981 14399 20039 14405
rect 19981 14396 19993 14399
rect 19751 14368 19993 14396
rect 19751 14365 19763 14368
rect 19705 14359 19763 14365
rect 19981 14365 19993 14368
rect 20027 14365 20039 14399
rect 19981 14359 20039 14365
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14396 20223 14399
rect 20254 14396 20260 14408
rect 20211 14368 20260 14396
rect 20211 14365 20223 14368
rect 20165 14359 20223 14365
rect 20254 14356 20260 14368
rect 20312 14356 20318 14408
rect 20438 14396 20444 14408
rect 20399 14368 20444 14396
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 20990 14356 20996 14408
rect 21048 14396 21054 14408
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 21048 14368 21097 14396
rect 21048 14356 21054 14368
rect 21085 14365 21097 14368
rect 21131 14365 21143 14399
rect 21085 14359 21143 14365
rect 21652 14328 21680 14436
rect 21729 14399 21787 14405
rect 21729 14365 21741 14399
rect 21775 14365 21787 14399
rect 22002 14396 22008 14408
rect 21963 14368 22008 14396
rect 21729 14359 21787 14365
rect 19527 14300 21680 14328
rect 21744 14328 21772 14359
rect 22002 14356 22008 14368
rect 22060 14356 22066 14408
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 22189 14399 22247 14405
rect 22189 14396 22201 14399
rect 22152 14368 22201 14396
rect 22152 14356 22158 14368
rect 22189 14365 22201 14368
rect 22235 14365 22247 14399
rect 22189 14359 22247 14365
rect 22462 14356 22468 14408
rect 22520 14396 22526 14408
rect 22557 14399 22615 14405
rect 22557 14396 22569 14399
rect 22520 14368 22569 14396
rect 22520 14356 22526 14368
rect 22557 14365 22569 14368
rect 22603 14365 22615 14399
rect 22557 14359 22615 14365
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14365 22707 14399
rect 22759 14396 22787 14436
rect 22833 14433 22845 14467
rect 22879 14433 22891 14467
rect 22833 14427 22891 14433
rect 23124 14436 23704 14464
rect 23124 14396 23152 14436
rect 22759 14368 23152 14396
rect 23196 14377 23254 14383
rect 22649 14359 22707 14365
rect 22664 14328 22692 14359
rect 23196 14343 23208 14377
rect 23242 14343 23254 14377
rect 23290 14356 23296 14408
rect 23348 14396 23354 14408
rect 23676 14405 23704 14436
rect 23569 14399 23627 14405
rect 23348 14368 23393 14396
rect 23348 14356 23354 14368
rect 23569 14365 23581 14399
rect 23615 14365 23627 14399
rect 23569 14359 23627 14365
rect 23661 14399 23719 14405
rect 23661 14365 23673 14399
rect 23707 14396 23719 14399
rect 23952 14396 23980 14495
rect 24578 14424 24584 14476
rect 24636 14464 24642 14476
rect 25133 14467 25191 14473
rect 25133 14464 25145 14467
rect 24636 14436 25145 14464
rect 24636 14424 24642 14436
rect 25133 14433 25145 14436
rect 25179 14433 25191 14467
rect 25133 14427 25191 14433
rect 25498 14424 25504 14476
rect 25556 14464 25562 14476
rect 25961 14467 26019 14473
rect 25961 14464 25973 14467
rect 25556 14436 25973 14464
rect 25556 14424 25562 14436
rect 25961 14433 25973 14436
rect 26007 14433 26019 14467
rect 25961 14427 26019 14433
rect 25038 14396 25044 14408
rect 23707 14368 23980 14396
rect 24999 14368 25044 14396
rect 23707 14365 23719 14368
rect 23661 14359 23719 14365
rect 23196 14340 23254 14343
rect 23014 14328 23020 14340
rect 21744 14300 22600 14328
rect 22664 14300 23020 14328
rect 22572 14272 22600 14300
rect 23014 14288 23020 14300
rect 23072 14288 23078 14340
rect 23196 14337 23204 14340
rect 23198 14288 23204 14337
rect 23256 14288 23262 14340
rect 23385 14331 23443 14337
rect 23385 14297 23397 14331
rect 23431 14297 23443 14331
rect 23584 14328 23612 14359
rect 25038 14356 25044 14368
rect 25096 14356 25102 14408
rect 25317 14399 25375 14405
rect 25317 14365 25329 14399
rect 25363 14365 25375 14399
rect 25317 14359 25375 14365
rect 26145 14399 26203 14405
rect 26145 14365 26157 14399
rect 26191 14396 26203 14399
rect 26510 14396 26516 14408
rect 26191 14368 26516 14396
rect 26191 14365 26203 14368
rect 26145 14359 26203 14365
rect 24854 14328 24860 14340
rect 23584 14300 24860 14328
rect 23385 14291 23443 14297
rect 17126 14260 17132 14272
rect 17052 14232 17132 14260
rect 16117 14223 16175 14229
rect 17126 14220 17132 14232
rect 17184 14220 17190 14272
rect 19242 14260 19248 14272
rect 19203 14232 19248 14260
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 20809 14263 20867 14269
rect 20809 14229 20821 14263
rect 20855 14260 20867 14263
rect 20898 14260 20904 14272
rect 20855 14232 20904 14260
rect 20855 14229 20867 14232
rect 20809 14223 20867 14229
rect 20898 14220 20904 14232
rect 20956 14220 20962 14272
rect 21634 14220 21640 14272
rect 21692 14260 21698 14272
rect 22094 14260 22100 14272
rect 21692 14232 22100 14260
rect 21692 14220 21698 14232
rect 22094 14220 22100 14232
rect 22152 14220 22158 14272
rect 22554 14220 22560 14272
rect 22612 14220 22618 14272
rect 22833 14263 22891 14269
rect 22833 14229 22845 14263
rect 22879 14260 22891 14263
rect 23400 14260 23428 14291
rect 24854 14288 24860 14300
rect 24912 14288 24918 14340
rect 25332 14328 25360 14359
rect 26510 14356 26516 14368
rect 26568 14356 26574 14408
rect 26786 14396 26792 14408
rect 26747 14368 26792 14396
rect 26786 14356 26792 14368
rect 26844 14356 26850 14408
rect 26970 14396 26976 14408
rect 26931 14368 26976 14396
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27062 14356 27068 14408
rect 27120 14396 27126 14408
rect 27233 14405 27261 14504
rect 27203 14399 27261 14405
rect 27120 14368 27165 14396
rect 27120 14356 27126 14368
rect 27203 14365 27215 14399
rect 27249 14396 27261 14399
rect 27709 14399 27767 14405
rect 27709 14396 27721 14399
rect 27249 14368 27721 14396
rect 27249 14365 27261 14368
rect 27203 14359 27261 14365
rect 27709 14365 27721 14368
rect 27755 14365 27767 14399
rect 28077 14399 28135 14405
rect 28077 14396 28089 14399
rect 27709 14359 27767 14365
rect 27816 14368 28089 14396
rect 25866 14328 25872 14340
rect 25056 14300 25360 14328
rect 25827 14300 25872 14328
rect 25056 14272 25084 14300
rect 25866 14288 25872 14300
rect 25924 14288 25930 14340
rect 26528 14328 26556 14356
rect 27816 14328 27844 14368
rect 28077 14365 28089 14368
rect 28123 14396 28135 14399
rect 28350 14396 28356 14408
rect 28123 14368 28356 14396
rect 28123 14365 28135 14368
rect 28077 14359 28135 14365
rect 28350 14356 28356 14368
rect 28408 14356 28414 14408
rect 26528 14300 27844 14328
rect 27890 14288 27896 14340
rect 27948 14328 27954 14340
rect 27948 14300 27993 14328
rect 27948 14288 27954 14300
rect 22879 14232 23428 14260
rect 22879 14229 22891 14232
rect 22833 14223 22891 14229
rect 23842 14220 23848 14272
rect 23900 14260 23906 14272
rect 24210 14260 24216 14272
rect 23900 14232 24216 14260
rect 23900 14220 23906 14232
rect 24210 14220 24216 14232
rect 24268 14220 24274 14272
rect 25038 14220 25044 14272
rect 25096 14220 25102 14272
rect 25498 14260 25504 14272
rect 25459 14232 25504 14260
rect 25498 14220 25504 14232
rect 25556 14220 25562 14272
rect 26326 14260 26332 14272
rect 26287 14232 26332 14260
rect 26326 14220 26332 14232
rect 26384 14220 26390 14272
rect 1104 14170 28888 14192
rect 1104 14118 10214 14170
rect 10266 14118 10278 14170
rect 10330 14118 10342 14170
rect 10394 14118 10406 14170
rect 10458 14118 10470 14170
rect 10522 14118 19478 14170
rect 19530 14118 19542 14170
rect 19594 14118 19606 14170
rect 19658 14118 19670 14170
rect 19722 14118 19734 14170
rect 19786 14118 28888 14170
rect 1104 14096 28888 14118
rect 5261 14059 5319 14065
rect 5261 14025 5273 14059
rect 5307 14056 5319 14059
rect 5902 14056 5908 14068
rect 5307 14028 5908 14056
rect 5307 14025 5319 14028
rect 5261 14019 5319 14025
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 6365 14059 6423 14065
rect 6365 14025 6377 14059
rect 6411 14025 6423 14059
rect 8938 14056 8944 14068
rect 8899 14028 8944 14056
rect 6365 14019 6423 14025
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13920 5135 13923
rect 5537 13923 5595 13929
rect 5537 13920 5549 13923
rect 5123 13892 5549 13920
rect 5123 13889 5135 13892
rect 5077 13883 5135 13889
rect 5537 13889 5549 13892
rect 5583 13889 5595 13923
rect 5537 13883 5595 13889
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13920 5779 13923
rect 6380 13920 6408 14019
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9217 14059 9275 14065
rect 9217 14025 9229 14059
rect 9263 14056 9275 14059
rect 9398 14056 9404 14068
rect 9263 14028 9404 14056
rect 9263 14025 9275 14028
rect 9217 14019 9275 14025
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9585 14059 9643 14065
rect 9585 14025 9597 14059
rect 9631 14056 9643 14059
rect 11606 14056 11612 14068
rect 9631 14028 11612 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 12526 14056 12532 14068
rect 12406 14028 12532 14056
rect 6822 13948 6828 14000
rect 6880 13948 6886 14000
rect 7828 13991 7886 13997
rect 7828 13957 7840 13991
rect 7874 13988 7886 13991
rect 8018 13988 8024 14000
rect 7874 13960 8024 13988
rect 7874 13957 7886 13960
rect 7828 13951 7886 13957
rect 8018 13948 8024 13960
rect 8076 13948 8082 14000
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 10042 13988 10048 14000
rect 8260 13960 10048 13988
rect 8260 13948 8266 13960
rect 5767 13892 6408 13920
rect 6733 13923 6791 13929
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 6840 13920 6868 13948
rect 9677 13923 9735 13929
rect 9677 13920 9689 13923
rect 6779 13892 9689 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 9677 13889 9689 13892
rect 9723 13889 9735 13923
rect 9677 13883 9735 13889
rect 5905 13855 5963 13861
rect 5905 13821 5917 13855
rect 5951 13852 5963 13855
rect 6546 13852 6552 13864
rect 5951 13824 6552 13852
rect 5951 13821 5963 13824
rect 5905 13815 5963 13821
rect 6546 13812 6552 13824
rect 6604 13812 6610 13864
rect 9784 13861 9812 13960
rect 10042 13948 10048 13960
rect 10100 13988 10106 14000
rect 10321 13991 10379 13997
rect 10321 13988 10333 13991
rect 10100 13960 10333 13988
rect 10100 13948 10106 13960
rect 10321 13957 10333 13960
rect 10367 13957 10379 13991
rect 10321 13951 10379 13957
rect 10505 13991 10563 13997
rect 10505 13957 10517 13991
rect 10551 13988 10563 13991
rect 10594 13988 10600 14000
rect 10551 13960 10600 13988
rect 10551 13957 10563 13960
rect 10505 13951 10563 13957
rect 10594 13948 10600 13960
rect 10652 13988 10658 14000
rect 12406 13988 12434 14028
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 12986 14016 12992 14068
rect 13044 14056 13050 14068
rect 13354 14056 13360 14068
rect 13044 14028 13360 14056
rect 13044 14016 13050 14028
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 13446 14016 13452 14068
rect 13504 14056 13510 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 13504 14028 17785 14056
rect 13504 14016 13510 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 18233 14059 18291 14065
rect 18233 14025 18245 14059
rect 18279 14056 18291 14059
rect 18414 14056 18420 14068
rect 18279 14028 18420 14056
rect 18279 14025 18291 14028
rect 18233 14019 18291 14025
rect 18414 14016 18420 14028
rect 18472 14016 18478 14068
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14056 20131 14059
rect 20254 14056 20260 14068
rect 20119 14028 20260 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 20254 14016 20260 14028
rect 20312 14056 20318 14068
rect 21634 14056 21640 14068
rect 20312 14028 21229 14056
rect 20312 14016 20318 14028
rect 13464 13988 13492 14016
rect 10652 13960 11100 13988
rect 10652 13948 10658 13960
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13889 11023 13923
rect 11072 13920 11100 13960
rect 11256 13960 12434 13988
rect 12728 13960 13492 13988
rect 11256 13920 11284 13960
rect 11072 13892 11284 13920
rect 11609 13923 11667 13929
rect 10965 13883 11023 13889
rect 11609 13889 11621 13923
rect 11655 13920 11667 13923
rect 11698 13920 11704 13932
rect 11655 13892 11704 13920
rect 11655 13889 11667 13892
rect 11609 13883 11667 13889
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 7561 13855 7619 13861
rect 7561 13821 7573 13855
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13821 9827 13855
rect 10980 13852 11008 13883
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 12728 13929 12756 13960
rect 14090 13948 14096 14000
rect 14148 13988 14154 14000
rect 14458 13988 14464 14000
rect 14148 13960 14464 13988
rect 14148 13948 14154 13960
rect 14458 13948 14464 13960
rect 14516 13988 14522 14000
rect 15289 13991 15347 13997
rect 15289 13988 15301 13991
rect 14516 13960 15301 13988
rect 14516 13948 14522 13960
rect 15289 13957 15301 13960
rect 15335 13957 15347 13991
rect 15289 13951 15347 13957
rect 15473 13991 15531 13997
rect 15473 13957 15485 13991
rect 15519 13988 15531 13991
rect 15930 13988 15936 14000
rect 15519 13960 15936 13988
rect 15519 13957 15531 13960
rect 15473 13951 15531 13957
rect 15930 13948 15936 13960
rect 15988 13948 15994 14000
rect 16025 13991 16083 13997
rect 16025 13957 16037 13991
rect 16071 13988 16083 13991
rect 16206 13988 16212 14000
rect 16071 13960 16212 13988
rect 16071 13957 16083 13960
rect 16025 13951 16083 13957
rect 16206 13948 16212 13960
rect 16264 13948 16270 14000
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13988 17095 13991
rect 17494 13988 17500 14000
rect 17083 13960 17500 13988
rect 17083 13957 17095 13960
rect 17037 13951 17095 13957
rect 17494 13948 17500 13960
rect 17552 13948 17558 14000
rect 18322 13948 18328 14000
rect 18380 13988 18386 14000
rect 18960 13991 19018 13997
rect 18380 13960 18736 13988
rect 18380 13948 18386 13960
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13889 12771 13923
rect 12986 13920 12992 13932
rect 12947 13892 12992 13920
rect 12713 13883 12771 13889
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 13078 13880 13084 13932
rect 13136 13920 13142 13932
rect 13265 13923 13323 13929
rect 13136 13892 13181 13920
rect 13136 13880 13142 13892
rect 13265 13889 13277 13923
rect 13311 13889 13323 13923
rect 13265 13883 13323 13889
rect 12342 13852 12348 13864
rect 10980 13824 12348 13852
rect 9769 13815 9827 13821
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 6840 13784 6868 13815
rect 6788 13756 6868 13784
rect 6788 13744 6794 13756
rect 6638 13676 6644 13728
rect 6696 13716 6702 13728
rect 6932 13716 6960 13815
rect 6696 13688 6960 13716
rect 6696 13676 6702 13688
rect 7190 13676 7196 13728
rect 7248 13716 7254 13728
rect 7576 13716 7604 13815
rect 12342 13812 12348 13824
rect 12400 13852 12406 13864
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12400 13824 12449 13852
rect 12400 13812 12406 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 13280 13852 13308 13883
rect 13354 13880 13360 13932
rect 13412 13920 13418 13932
rect 13495 13923 13553 13929
rect 13412 13892 13457 13920
rect 13412 13880 13418 13892
rect 13495 13889 13507 13923
rect 13541 13920 13553 13923
rect 13722 13920 13728 13932
rect 13541 13892 13728 13920
rect 13541 13889 13553 13892
rect 13495 13883 13553 13889
rect 13722 13880 13728 13892
rect 13780 13920 13786 13932
rect 13780 13892 14504 13920
rect 13780 13880 13786 13892
rect 13630 13852 13636 13864
rect 13280 13824 13636 13852
rect 12437 13815 12495 13821
rect 13630 13812 13636 13824
rect 13688 13852 13694 13864
rect 14366 13852 14372 13864
rect 13688 13824 14372 13852
rect 13688 13812 13694 13824
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 14476 13861 14504 13892
rect 16758 13880 16764 13932
rect 16816 13920 16822 13932
rect 17405 13923 17463 13929
rect 17405 13920 17417 13923
rect 16816 13892 17417 13920
rect 16816 13880 16822 13892
rect 17405 13889 17417 13892
rect 17451 13889 17463 13923
rect 17405 13883 17463 13889
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 18414 13920 18420 13932
rect 17911 13892 18420 13920
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 18414 13880 18420 13892
rect 18472 13880 18478 13932
rect 18708 13929 18736 13960
rect 18960 13957 18972 13991
rect 19006 13988 19018 13991
rect 19242 13988 19248 14000
rect 19006 13960 19248 13988
rect 19006 13957 19018 13960
rect 18960 13951 19018 13957
rect 19242 13948 19248 13960
rect 19300 13948 19306 14000
rect 21082 13988 21088 14000
rect 20732 13960 21088 13988
rect 18693 13923 18751 13929
rect 18693 13889 18705 13923
rect 18739 13889 18751 13923
rect 20438 13920 20444 13932
rect 20399 13892 20444 13920
rect 18693 13883 18751 13889
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 20530 13880 20536 13932
rect 20588 13920 20594 13932
rect 20732 13929 20760 13960
rect 21082 13948 21088 13960
rect 21140 13948 21146 14000
rect 20717 13923 20775 13929
rect 20588 13892 20633 13920
rect 20588 13880 20594 13892
rect 20717 13889 20729 13923
rect 20763 13889 20775 13923
rect 20717 13883 20775 13889
rect 20806 13880 20812 13932
rect 20864 13920 20870 13932
rect 20864 13892 20909 13920
rect 20864 13880 20870 13892
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13821 14519 13855
rect 14461 13815 14519 13821
rect 14737 13855 14795 13861
rect 14737 13821 14749 13855
rect 14783 13821 14795 13855
rect 14737 13815 14795 13821
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13852 15623 13855
rect 17034 13852 17040 13864
rect 15611 13824 17040 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 11146 13784 11152 13796
rect 8496 13756 9812 13784
rect 11107 13756 11152 13784
rect 7834 13716 7840 13728
rect 7248 13688 7840 13716
rect 7248 13676 7254 13688
rect 7834 13676 7840 13688
rect 7892 13716 7898 13728
rect 8496 13716 8524 13756
rect 9784 13728 9812 13756
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 14090 13744 14096 13796
rect 14148 13784 14154 13796
rect 14752 13784 14780 13815
rect 14148 13756 14780 13784
rect 16025 13787 16083 13793
rect 14148 13744 14154 13756
rect 16025 13753 16037 13787
rect 16071 13784 16083 13787
rect 16574 13784 16580 13796
rect 16071 13756 16580 13784
rect 16071 13753 16083 13756
rect 16025 13747 16083 13753
rect 16574 13744 16580 13756
rect 16632 13744 16638 13796
rect 16868 13793 16896 13824
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 20456 13852 20484 13880
rect 21082 13852 21088 13864
rect 20456 13824 21088 13852
rect 21082 13812 21088 13824
rect 21140 13812 21146 13864
rect 21201 13852 21229 14028
rect 21284 14028 21640 14056
rect 21284 13929 21312 14028
rect 21634 14016 21640 14028
rect 21692 14016 21698 14068
rect 22554 14016 22560 14068
rect 22612 14056 22618 14068
rect 23290 14056 23296 14068
rect 22612 14028 22657 14056
rect 23251 14028 23296 14056
rect 22612 14016 22618 14028
rect 23290 14016 23296 14028
rect 23348 14016 23354 14068
rect 23658 14016 23664 14068
rect 23716 14056 23722 14068
rect 23716 14028 23980 14056
rect 23716 14016 23722 14028
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 21453 13923 21511 13929
rect 21453 13889 21465 13923
rect 21499 13920 21511 13923
rect 21542 13920 21548 13932
rect 21499 13892 21548 13920
rect 21499 13889 21511 13892
rect 21453 13883 21511 13889
rect 21542 13880 21548 13892
rect 21600 13880 21606 13932
rect 21634 13880 21640 13932
rect 21692 13920 21698 13932
rect 21810 13923 21868 13929
rect 21810 13920 21822 13923
rect 21692 13892 21822 13920
rect 21692 13880 21698 13892
rect 21810 13889 21822 13892
rect 21856 13889 21868 13923
rect 21810 13883 21868 13889
rect 22137 13923 22195 13929
rect 22137 13889 22149 13923
rect 22183 13920 22195 13923
rect 22278 13920 22284 13932
rect 22183 13892 22284 13920
rect 22183 13889 22195 13892
rect 22137 13883 22195 13889
rect 22278 13880 22284 13892
rect 22336 13880 22342 13932
rect 22925 13923 22983 13929
rect 22925 13889 22937 13923
rect 22971 13920 22983 13923
rect 23198 13920 23204 13932
rect 22971 13892 23204 13920
rect 22971 13889 22983 13892
rect 22925 13883 22983 13889
rect 23198 13880 23204 13892
rect 23256 13880 23262 13932
rect 23952 13929 23980 14028
rect 24118 14016 24124 14068
rect 24176 14056 24182 14068
rect 25225 14059 25283 14065
rect 24176 14028 24900 14056
rect 24176 14016 24182 14028
rect 24026 13948 24032 14000
rect 24084 13988 24090 14000
rect 24397 13991 24455 13997
rect 24397 13988 24409 13991
rect 24084 13960 24409 13988
rect 24084 13948 24090 13960
rect 24397 13957 24409 13960
rect 24443 13957 24455 13991
rect 24397 13951 24455 13957
rect 24578 13948 24584 14000
rect 24636 13988 24642 14000
rect 24765 13991 24823 13997
rect 24765 13988 24777 13991
rect 24636 13960 24777 13988
rect 24636 13948 24642 13960
rect 24765 13957 24777 13960
rect 24811 13957 24823 13991
rect 24765 13951 24823 13957
rect 23753 13923 23811 13929
rect 23753 13889 23765 13923
rect 23799 13889 23811 13923
rect 23753 13883 23811 13889
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 24210 13920 24216 13932
rect 24171 13892 24216 13920
rect 23937 13883 23995 13889
rect 22005 13855 22063 13861
rect 22005 13852 22017 13855
rect 21201 13824 22017 13852
rect 22005 13821 22017 13824
rect 22051 13852 22063 13855
rect 22833 13855 22891 13861
rect 22833 13852 22845 13855
rect 22051 13824 22845 13852
rect 22051 13821 22063 13824
rect 22005 13815 22063 13821
rect 22833 13821 22845 13824
rect 22879 13821 22891 13855
rect 22833 13815 22891 13821
rect 23014 13812 23020 13864
rect 23072 13852 23078 13864
rect 23566 13852 23572 13864
rect 23072 13824 23572 13852
rect 23072 13812 23078 13824
rect 23566 13812 23572 13824
rect 23624 13812 23630 13864
rect 23768 13852 23796 13883
rect 23952 13852 23980 13883
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 24489 13923 24547 13929
rect 24489 13889 24501 13923
rect 24535 13920 24547 13923
rect 24670 13920 24676 13932
rect 24535 13892 24676 13920
rect 24535 13889 24547 13892
rect 24489 13883 24547 13889
rect 24670 13880 24676 13892
rect 24728 13880 24734 13932
rect 24872 13920 24900 14028
rect 25225 14025 25237 14059
rect 25271 14056 25283 14059
rect 25866 14056 25872 14068
rect 25271 14028 25872 14056
rect 25271 14025 25283 14028
rect 25225 14019 25283 14025
rect 25866 14016 25872 14028
rect 25924 14016 25930 14068
rect 26786 14016 26792 14068
rect 26844 14056 26850 14068
rect 27433 14059 27491 14065
rect 27433 14056 27445 14059
rect 26844 14028 27445 14056
rect 26844 14016 26850 14028
rect 27433 14025 27445 14028
rect 27479 14025 27491 14059
rect 27433 14019 27491 14025
rect 26326 13988 26332 14000
rect 26287 13960 26332 13988
rect 26326 13948 26332 13960
rect 26384 13948 26390 14000
rect 27890 13988 27896 14000
rect 26528 13960 27896 13988
rect 25041 13923 25099 13929
rect 25041 13920 25053 13923
rect 24872 13892 25053 13920
rect 25041 13889 25053 13892
rect 25087 13889 25099 13923
rect 25041 13883 25099 13889
rect 26145 13923 26203 13929
rect 26145 13889 26157 13923
rect 26191 13889 26203 13923
rect 26145 13883 26203 13889
rect 24578 13852 24584 13864
rect 23768 13824 23888 13852
rect 23952 13824 24584 13852
rect 16853 13787 16911 13793
rect 16853 13753 16865 13787
rect 16899 13753 16911 13787
rect 23290 13784 23296 13796
rect 16853 13747 16911 13753
rect 16960 13756 17264 13784
rect 7892 13688 8524 13716
rect 7892 13676 7898 13688
rect 9766 13676 9772 13728
rect 9824 13676 9830 13728
rect 13633 13719 13691 13725
rect 13633 13685 13645 13719
rect 13679 13716 13691 13719
rect 13906 13716 13912 13728
rect 13679 13688 13912 13716
rect 13679 13685 13691 13688
rect 13633 13679 13691 13685
rect 13906 13676 13912 13688
rect 13964 13676 13970 13728
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 16960 13716 16988 13756
rect 15344 13688 16988 13716
rect 17037 13719 17095 13725
rect 15344 13676 15350 13688
rect 17037 13685 17049 13719
rect 17083 13716 17095 13719
rect 17126 13716 17132 13728
rect 17083 13688 17132 13716
rect 17083 13685 17095 13688
rect 17037 13679 17095 13685
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 17236 13716 17264 13756
rect 20548 13756 23296 13784
rect 20548 13716 20576 13756
rect 23290 13744 23296 13756
rect 23348 13744 23354 13796
rect 23860 13784 23888 13824
rect 24578 13812 24584 13824
rect 24636 13812 24642 13864
rect 24854 13852 24860 13864
rect 24815 13824 24860 13852
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 26160 13852 26188 13883
rect 26234 13880 26240 13932
rect 26292 13920 26298 13932
rect 26528 13929 26556 13960
rect 27890 13948 27896 13960
rect 27948 13948 27954 14000
rect 26513 13923 26571 13929
rect 26292 13892 26337 13920
rect 26292 13880 26298 13892
rect 26513 13889 26525 13923
rect 26559 13889 26571 13923
rect 26970 13920 26976 13932
rect 26931 13892 26976 13920
rect 26513 13883 26571 13889
rect 26970 13880 26976 13892
rect 27028 13880 27034 13932
rect 28258 13920 28264 13932
rect 28219 13892 28264 13920
rect 28258 13880 28264 13892
rect 28316 13880 28322 13932
rect 27062 13852 27068 13864
rect 26160 13824 27068 13852
rect 27062 13812 27068 13824
rect 27120 13812 27126 13864
rect 23860 13756 25084 13784
rect 25056 13728 25084 13756
rect 25682 13744 25688 13796
rect 25740 13784 25746 13796
rect 28077 13787 28135 13793
rect 28077 13784 28089 13787
rect 25740 13756 28089 13784
rect 25740 13744 25746 13756
rect 28077 13753 28089 13756
rect 28123 13753 28135 13787
rect 28077 13747 28135 13753
rect 17236 13688 20576 13716
rect 20622 13676 20628 13728
rect 20680 13716 20686 13728
rect 20993 13719 21051 13725
rect 20993 13716 21005 13719
rect 20680 13688 21005 13716
rect 20680 13676 20686 13688
rect 20993 13685 21005 13688
rect 21039 13685 21051 13719
rect 21450 13716 21456 13728
rect 21411 13688 21456 13716
rect 20993 13679 21051 13685
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 21726 13676 21732 13728
rect 21784 13716 21790 13728
rect 21821 13719 21879 13725
rect 21821 13716 21833 13719
rect 21784 13688 21833 13716
rect 21784 13676 21790 13688
rect 21821 13685 21833 13688
rect 21867 13685 21879 13719
rect 22278 13716 22284 13728
rect 22239 13688 22284 13716
rect 21821 13679 21879 13685
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 22370 13676 22376 13728
rect 22428 13716 22434 13728
rect 22741 13719 22799 13725
rect 22741 13716 22753 13719
rect 22428 13688 22753 13716
rect 22428 13676 22434 13688
rect 22741 13685 22753 13688
rect 22787 13685 22799 13719
rect 22741 13679 22799 13685
rect 24213 13719 24271 13725
rect 24213 13685 24225 13719
rect 24259 13716 24271 13719
rect 24486 13716 24492 13728
rect 24259 13688 24492 13716
rect 24259 13685 24271 13688
rect 24213 13679 24271 13685
rect 24486 13676 24492 13688
rect 24544 13676 24550 13728
rect 25038 13716 25044 13728
rect 24999 13688 25044 13716
rect 25038 13676 25044 13688
rect 25096 13676 25102 13728
rect 25958 13716 25964 13728
rect 25919 13688 25964 13716
rect 25958 13676 25964 13688
rect 26016 13676 26022 13728
rect 27154 13716 27160 13728
rect 27115 13688 27160 13716
rect 27154 13676 27160 13688
rect 27212 13676 27218 13728
rect 1104 13626 28888 13648
rect 1104 13574 5582 13626
rect 5634 13574 5646 13626
rect 5698 13574 5710 13626
rect 5762 13574 5774 13626
rect 5826 13574 5838 13626
rect 5890 13574 14846 13626
rect 14898 13574 14910 13626
rect 14962 13574 14974 13626
rect 15026 13574 15038 13626
rect 15090 13574 15102 13626
rect 15154 13574 24110 13626
rect 24162 13574 24174 13626
rect 24226 13574 24238 13626
rect 24290 13574 24302 13626
rect 24354 13574 24366 13626
rect 24418 13574 28888 13626
rect 1104 13552 28888 13574
rect 7190 13512 7196 13524
rect 5276 13484 7196 13512
rect 5166 13336 5172 13388
rect 5224 13376 5230 13388
rect 5276 13385 5304 13484
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7558 13472 7564 13524
rect 7616 13512 7622 13524
rect 7653 13515 7711 13521
rect 7653 13512 7665 13515
rect 7616 13484 7665 13512
rect 7616 13472 7622 13484
rect 7653 13481 7665 13484
rect 7699 13481 7711 13515
rect 7653 13475 7711 13481
rect 13725 13515 13783 13521
rect 13725 13481 13737 13515
rect 13771 13512 13783 13515
rect 15838 13512 15844 13524
rect 13771 13484 15844 13512
rect 13771 13481 13783 13484
rect 13725 13475 13783 13481
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 17126 13472 17132 13524
rect 17184 13512 17190 13524
rect 18325 13515 18383 13521
rect 18325 13512 18337 13515
rect 17184 13484 18337 13512
rect 17184 13472 17190 13484
rect 18325 13481 18337 13484
rect 18371 13512 18383 13515
rect 18598 13512 18604 13524
rect 18371 13484 18604 13512
rect 18371 13481 18383 13484
rect 18325 13475 18383 13481
rect 18598 13472 18604 13484
rect 18656 13472 18662 13524
rect 20254 13512 20260 13524
rect 18708 13484 20260 13512
rect 6641 13447 6699 13453
rect 6641 13413 6653 13447
rect 6687 13413 6699 13447
rect 9674 13444 9680 13456
rect 6641 13407 6699 13413
rect 9048 13416 9680 13444
rect 5261 13379 5319 13385
rect 5261 13376 5273 13379
rect 5224 13348 5273 13376
rect 5224 13336 5230 13348
rect 5261 13345 5273 13348
rect 5307 13345 5319 13379
rect 6656 13376 6684 13407
rect 6730 13376 6736 13388
rect 6643 13348 6736 13376
rect 5261 13339 5319 13345
rect 6730 13336 6736 13348
rect 6788 13376 6794 13388
rect 8113 13379 8171 13385
rect 8113 13376 8125 13379
rect 6788 13348 8125 13376
rect 6788 13336 6794 13348
rect 8113 13345 8125 13348
rect 8159 13345 8171 13379
rect 8113 13339 8171 13345
rect 8202 13336 8208 13388
rect 8260 13376 8266 13388
rect 9048 13385 9076 13416
rect 9674 13404 9680 13416
rect 9732 13404 9738 13456
rect 14458 13444 14464 13456
rect 13096 13416 14464 13444
rect 9033 13379 9091 13385
rect 8260 13348 8305 13376
rect 8260 13336 8266 13348
rect 9033 13345 9045 13379
rect 9079 13345 9091 13379
rect 9033 13339 9091 13345
rect 5528 13311 5586 13317
rect 5528 13277 5540 13311
rect 5574 13308 5586 13311
rect 5902 13308 5908 13320
rect 5574 13280 5908 13308
rect 5574 13277 5586 13280
rect 5528 13271 5586 13277
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13308 8079 13311
rect 8938 13308 8944 13320
rect 8067 13280 8944 13308
rect 8067 13277 8079 13280
rect 8021 13271 8079 13277
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 9214 13308 9220 13320
rect 9175 13280 9220 13308
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 9766 13308 9772 13320
rect 9723 13280 9772 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 13096 13317 13124 13416
rect 14458 13404 14464 13416
rect 14516 13404 14522 13456
rect 16209 13447 16267 13453
rect 16209 13413 16221 13447
rect 16255 13444 16267 13447
rect 16574 13444 16580 13456
rect 16255 13416 16580 13444
rect 16255 13413 16267 13416
rect 16209 13407 16267 13413
rect 16574 13404 16580 13416
rect 16632 13404 16638 13456
rect 18708 13453 18736 13484
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 21634 13512 21640 13524
rect 21140 13484 21640 13512
rect 21140 13472 21146 13484
rect 21634 13472 21640 13484
rect 21692 13512 21698 13524
rect 21729 13515 21787 13521
rect 21729 13512 21741 13515
rect 21692 13484 21741 13512
rect 21692 13472 21698 13484
rect 21729 13481 21741 13484
rect 21775 13512 21787 13515
rect 21818 13512 21824 13524
rect 21775 13484 21824 13512
rect 21775 13481 21787 13484
rect 21729 13475 21787 13481
rect 21818 13472 21824 13484
rect 21876 13472 21882 13524
rect 21910 13472 21916 13524
rect 21968 13512 21974 13524
rect 21968 13484 22094 13512
rect 21968 13472 21974 13484
rect 18693 13447 18751 13453
rect 18693 13444 18705 13447
rect 17052 13416 18705 13444
rect 14366 13376 14372 13388
rect 13372 13348 14136 13376
rect 14327 13348 14372 13376
rect 13372 13317 13400 13348
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11204 13280 11345 13308
rect 11204 13268 11210 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 13174 13311 13232 13317
rect 13174 13277 13186 13311
rect 13220 13277 13232 13311
rect 13174 13271 13232 13277
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 13587 13311 13645 13317
rect 13587 13277 13599 13311
rect 13633 13308 13645 13311
rect 13998 13308 14004 13320
rect 13633 13280 14004 13308
rect 13633 13277 13645 13280
rect 13587 13271 13645 13277
rect 7285 13243 7343 13249
rect 7285 13209 7297 13243
rect 7331 13240 7343 13243
rect 9122 13240 9128 13252
rect 7331 13212 9128 13240
rect 7331 13209 7343 13212
rect 7285 13203 7343 13209
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 9944 13243 10002 13249
rect 9944 13209 9956 13243
rect 9990 13240 10002 13243
rect 10870 13240 10876 13252
rect 9990 13212 10876 13240
rect 9990 13209 10002 13212
rect 9944 13203 10002 13209
rect 10870 13200 10876 13212
rect 10928 13200 10934 13252
rect 11606 13249 11612 13252
rect 11600 13203 11612 13249
rect 11664 13240 11670 13252
rect 13188 13240 13216 13271
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 14108 13317 14136 13348
rect 14366 13336 14372 13348
rect 14424 13336 14430 13388
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13376 15715 13379
rect 15930 13376 15936 13388
rect 15703 13348 15936 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 15930 13336 15936 13348
rect 15988 13336 15994 13388
rect 16758 13336 16764 13388
rect 16816 13376 16822 13388
rect 17052 13385 17080 13416
rect 17037 13379 17095 13385
rect 17037 13376 17049 13379
rect 16816 13348 17049 13376
rect 16816 13336 16822 13348
rect 17037 13345 17049 13348
rect 17083 13345 17095 13379
rect 17037 13339 17095 13345
rect 17221 13379 17279 13385
rect 17221 13345 17233 13379
rect 17267 13376 17279 13379
rect 17267 13348 17816 13376
rect 17267 13345 17279 13348
rect 17221 13339 17279 13345
rect 14093 13311 14151 13317
rect 14093 13277 14105 13311
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 11664 13212 11700 13240
rect 12406 13212 13216 13240
rect 11606 13200 11612 13203
rect 11664 13200 11670 13212
rect 9401 13175 9459 13181
rect 9401 13141 9413 13175
rect 9447 13172 9459 13175
rect 10962 13172 10968 13184
rect 9447 13144 10968 13172
rect 9447 13141 9459 13144
rect 9401 13135 9459 13141
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 12406 13172 12434 13212
rect 13446 13200 13452 13252
rect 13504 13240 13510 13252
rect 14108 13240 14136 13271
rect 14182 13268 14188 13320
rect 14240 13308 14246 13320
rect 17126 13308 17132 13320
rect 14240 13280 17132 13308
rect 14240 13268 14246 13280
rect 17126 13268 17132 13280
rect 17184 13308 17190 13320
rect 17788 13317 17816 13348
rect 17880 13317 17908 13416
rect 18693 13413 18705 13416
rect 18739 13413 18751 13447
rect 18693 13407 18751 13413
rect 19886 13404 19892 13456
rect 19944 13444 19950 13456
rect 20070 13444 20076 13456
rect 19944 13416 20076 13444
rect 19944 13404 19950 13416
rect 20070 13404 20076 13416
rect 20128 13404 20134 13456
rect 18414 13336 18420 13388
rect 18472 13376 18478 13388
rect 19245 13379 19303 13385
rect 19245 13376 19257 13379
rect 18472 13348 19257 13376
rect 18472 13336 18478 13348
rect 19245 13345 19257 13348
rect 19291 13376 19303 13379
rect 19794 13376 19800 13388
rect 19291 13348 19800 13376
rect 19291 13345 19303 13348
rect 19245 13339 19303 13345
rect 19794 13336 19800 13348
rect 19852 13336 19858 13388
rect 19978 13336 19984 13388
rect 20036 13376 20042 13388
rect 20349 13379 20407 13385
rect 20349 13376 20361 13379
rect 20036 13348 20361 13376
rect 20036 13336 20042 13348
rect 20349 13345 20361 13348
rect 20395 13345 20407 13379
rect 22066 13376 22094 13484
rect 22278 13472 22284 13524
rect 22336 13512 22342 13524
rect 23658 13512 23664 13524
rect 22336 13484 23664 13512
rect 22336 13472 22342 13484
rect 23658 13472 23664 13484
rect 23716 13512 23722 13524
rect 23845 13515 23903 13521
rect 23845 13512 23857 13515
rect 23716 13484 23857 13512
rect 23716 13472 23722 13484
rect 23845 13481 23857 13484
rect 23891 13481 23903 13515
rect 23845 13475 23903 13481
rect 23937 13515 23995 13521
rect 23937 13481 23949 13515
rect 23983 13512 23995 13515
rect 24026 13512 24032 13524
rect 23983 13484 24032 13512
rect 23983 13481 23995 13484
rect 23937 13475 23995 13481
rect 24026 13472 24032 13484
rect 24084 13472 24090 13524
rect 24397 13515 24455 13521
rect 24397 13481 24409 13515
rect 24443 13481 24455 13515
rect 24397 13475 24455 13481
rect 23566 13404 23572 13456
rect 23624 13444 23630 13456
rect 24412 13444 24440 13475
rect 24670 13472 24676 13524
rect 24728 13512 24734 13524
rect 24765 13515 24823 13521
rect 24765 13512 24777 13515
rect 24728 13484 24777 13512
rect 24728 13472 24734 13484
rect 24765 13481 24777 13484
rect 24811 13481 24823 13515
rect 24765 13475 24823 13481
rect 26421 13515 26479 13521
rect 26421 13481 26433 13515
rect 26467 13512 26479 13515
rect 26970 13512 26976 13524
rect 26467 13484 26976 13512
rect 26467 13481 26479 13484
rect 26421 13475 26479 13481
rect 26970 13472 26976 13484
rect 27028 13472 27034 13524
rect 28353 13515 28411 13521
rect 28353 13481 28365 13515
rect 28399 13512 28411 13515
rect 28442 13512 28448 13524
rect 28399 13484 28448 13512
rect 28399 13481 28411 13484
rect 28353 13475 28411 13481
rect 28442 13472 28448 13484
rect 28500 13472 28506 13524
rect 23624 13416 24440 13444
rect 23624 13404 23630 13416
rect 22373 13379 22431 13385
rect 22373 13376 22385 13379
rect 22066 13348 22385 13376
rect 20349 13339 20407 13345
rect 22373 13345 22385 13348
rect 22419 13376 22431 13379
rect 24029 13379 24087 13385
rect 22419 13348 23796 13376
rect 22419 13345 22431 13348
rect 22373 13339 22431 13345
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 17184 13280 17693 13308
rect 17184 13268 17190 13280
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 17865 13311 17923 13317
rect 17865 13277 17877 13311
rect 17911 13277 17923 13311
rect 17865 13271 17923 13277
rect 16206 13240 16212 13252
rect 13504 13212 13549 13240
rect 14108 13212 14872 13240
rect 16167 13212 16212 13240
rect 13504 13200 13510 13212
rect 14844 13184 14872 13212
rect 16206 13200 16212 13212
rect 16264 13200 16270 13252
rect 17788 13240 17816 13271
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 19521 13311 19579 13317
rect 19521 13308 19533 13311
rect 19392 13280 19533 13308
rect 19392 13268 19398 13280
rect 19521 13277 19533 13280
rect 19567 13308 19579 13311
rect 19886 13308 19892 13320
rect 19567 13280 19892 13308
rect 19567 13277 19579 13280
rect 19521 13271 19579 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 22189 13311 22247 13317
rect 22189 13277 22201 13311
rect 22235 13308 22247 13311
rect 22649 13311 22707 13317
rect 22235 13280 22600 13308
rect 22235 13277 22247 13280
rect 22189 13271 22247 13277
rect 18506 13240 18512 13252
rect 17788 13212 18512 13240
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 20438 13200 20444 13252
rect 20496 13240 20502 13252
rect 20594 13243 20652 13249
rect 20594 13240 20606 13243
rect 20496 13212 20606 13240
rect 20496 13200 20502 13212
rect 20594 13209 20606 13212
rect 20640 13209 20652 13243
rect 22572 13240 22600 13280
rect 22649 13277 22661 13311
rect 22695 13308 22707 13311
rect 22738 13308 22744 13320
rect 22695 13280 22744 13308
rect 22695 13277 22707 13280
rect 22649 13271 22707 13277
rect 22738 13268 22744 13280
rect 22796 13268 22802 13320
rect 22925 13311 22983 13317
rect 22925 13277 22937 13311
rect 22971 13308 22983 13311
rect 23198 13308 23204 13320
rect 22971 13280 23204 13308
rect 22971 13277 22983 13280
rect 22925 13271 22983 13277
rect 22940 13240 22968 13271
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 23768 13317 23796 13348
rect 24029 13345 24041 13379
rect 24075 13376 24087 13379
rect 25038 13376 25044 13388
rect 24075 13348 25044 13376
rect 24075 13345 24087 13348
rect 24029 13339 24087 13345
rect 25038 13336 25044 13348
rect 25096 13336 25102 13388
rect 26142 13336 26148 13388
rect 26200 13376 26206 13388
rect 26973 13379 27031 13385
rect 26973 13376 26985 13379
rect 26200 13348 26985 13376
rect 26200 13336 26206 13348
rect 26973 13345 26985 13348
rect 27019 13345 27031 13379
rect 26973 13339 27031 13345
rect 23753 13311 23811 13317
rect 23753 13277 23765 13311
rect 23799 13277 23811 13311
rect 24394 13308 24400 13320
rect 24355 13280 24400 13308
rect 23753 13271 23811 13277
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 24489 13311 24547 13317
rect 24489 13277 24501 13311
rect 24535 13277 24547 13311
rect 25866 13308 25872 13320
rect 24489 13271 24547 13277
rect 24596 13280 25872 13308
rect 24504 13240 24532 13271
rect 22572 13212 22968 13240
rect 23216 13212 24532 13240
rect 20594 13203 20652 13209
rect 12710 13172 12716 13184
rect 11112 13144 12434 13172
rect 12671 13144 12716 13172
rect 11112 13132 11118 13144
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 15473 13175 15531 13181
rect 15473 13172 15485 13175
rect 14884 13144 15485 13172
rect 14884 13132 14890 13144
rect 15473 13141 15485 13144
rect 15519 13141 15531 13175
rect 15473 13135 15531 13141
rect 15749 13175 15807 13181
rect 15749 13141 15761 13175
rect 15795 13172 15807 13175
rect 16022 13172 16028 13184
rect 15795 13144 16028 13172
rect 15795 13141 15807 13144
rect 15749 13135 15807 13141
rect 16022 13132 16028 13144
rect 16080 13172 16086 13184
rect 16853 13175 16911 13181
rect 16853 13172 16865 13175
rect 16080 13144 16865 13172
rect 16080 13132 16086 13144
rect 16853 13141 16865 13144
rect 16899 13141 16911 13175
rect 18046 13172 18052 13184
rect 18007 13144 18052 13172
rect 16853 13135 16911 13141
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 20346 13132 20352 13184
rect 20404 13172 20410 13184
rect 21082 13172 21088 13184
rect 20404 13144 21088 13172
rect 20404 13132 20410 13144
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 21818 13132 21824 13184
rect 21876 13172 21882 13184
rect 22370 13172 22376 13184
rect 21876 13144 22376 13172
rect 21876 13132 21882 13144
rect 22370 13132 22376 13144
rect 22428 13132 22434 13184
rect 22462 13132 22468 13184
rect 22520 13172 22526 13184
rect 23216 13172 23244 13212
rect 22520 13144 23244 13172
rect 22520 13132 22526 13144
rect 23290 13132 23296 13184
rect 23348 13172 23354 13184
rect 24596 13172 24624 13280
rect 25866 13268 25872 13280
rect 25924 13308 25930 13320
rect 26053 13311 26111 13317
rect 26053 13308 26065 13311
rect 25924 13280 26065 13308
rect 25924 13268 25930 13280
rect 26053 13277 26065 13280
rect 26099 13277 26111 13311
rect 26053 13271 26111 13277
rect 26237 13311 26295 13317
rect 26237 13277 26249 13311
rect 26283 13277 26295 13311
rect 26237 13271 26295 13277
rect 25314 13200 25320 13252
rect 25372 13240 25378 13252
rect 25501 13243 25559 13249
rect 25501 13240 25513 13243
rect 25372 13212 25513 13240
rect 25372 13200 25378 13212
rect 25501 13209 25513 13212
rect 25547 13209 25559 13243
rect 25682 13240 25688 13252
rect 25643 13212 25688 13240
rect 25501 13203 25559 13209
rect 25682 13200 25688 13212
rect 25740 13200 25746 13252
rect 25958 13200 25964 13252
rect 26016 13240 26022 13252
rect 26252 13240 26280 13271
rect 27246 13249 27252 13252
rect 26016 13212 26280 13240
rect 26016 13200 26022 13212
rect 27240 13203 27252 13249
rect 27304 13240 27310 13252
rect 27304 13212 27340 13240
rect 27246 13200 27252 13203
rect 27304 13200 27310 13212
rect 23348 13144 24624 13172
rect 23348 13132 23354 13144
rect 1104 13082 28888 13104
rect 1104 13030 10214 13082
rect 10266 13030 10278 13082
rect 10330 13030 10342 13082
rect 10394 13030 10406 13082
rect 10458 13030 10470 13082
rect 10522 13030 19478 13082
rect 19530 13030 19542 13082
rect 19594 13030 19606 13082
rect 19658 13030 19670 13082
rect 19722 13030 19734 13082
rect 19786 13030 28888 13082
rect 1104 13008 28888 13030
rect 6730 12968 6736 12980
rect 6691 12940 6736 12968
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 9272 12940 9965 12968
rect 9272 12928 9278 12940
rect 9953 12937 9965 12940
rect 9999 12937 10011 12971
rect 9953 12931 10011 12937
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10928 12940 10977 12968
rect 10928 12928 10934 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 11517 12971 11575 12977
rect 11517 12937 11529 12971
rect 11563 12968 11575 12971
rect 11606 12968 11612 12980
rect 11563 12940 11612 12968
rect 11563 12937 11575 12940
rect 11517 12931 11575 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 12492 12940 12633 12968
rect 12492 12928 12498 12940
rect 12621 12937 12633 12940
rect 12667 12937 12679 12971
rect 12621 12931 12679 12937
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 14277 12971 14335 12977
rect 12768 12940 13860 12968
rect 12768 12928 12774 12940
rect 5810 12860 5816 12912
rect 5868 12900 5874 12912
rect 5994 12900 6000 12912
rect 5868 12872 6000 12900
rect 5868 12860 5874 12872
rect 5994 12860 6000 12872
rect 6052 12900 6058 12912
rect 6546 12900 6552 12912
rect 6052 12872 6552 12900
rect 6052 12860 6058 12872
rect 6546 12860 6552 12872
rect 6604 12900 6610 12912
rect 7377 12903 7435 12909
rect 7377 12900 7389 12903
rect 6604 12872 7389 12900
rect 6604 12860 6610 12872
rect 7377 12869 7389 12872
rect 7423 12869 7435 12903
rect 7377 12863 7435 12869
rect 10321 12903 10379 12909
rect 10321 12869 10333 12903
rect 10367 12900 10379 12903
rect 11054 12900 11060 12912
rect 10367 12872 11060 12900
rect 10367 12869 10379 12872
rect 10321 12863 10379 12869
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 12406 12872 13768 12900
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12832 5043 12835
rect 5445 12835 5503 12841
rect 5445 12832 5457 12835
rect 5031 12804 5457 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5445 12801 5457 12804
rect 5491 12801 5503 12835
rect 5445 12795 5503 12801
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12832 5687 12835
rect 5675 12804 6408 12832
rect 5675 12801 5687 12804
rect 5629 12795 5687 12801
rect 5810 12764 5816 12776
rect 5771 12736 5816 12764
rect 5810 12724 5816 12736
rect 5868 12724 5874 12776
rect 6380 12705 6408 12804
rect 6638 12792 6644 12844
rect 6696 12832 6702 12844
rect 7834 12832 7840 12844
rect 6696 12804 6960 12832
rect 7795 12804 7840 12832
rect 6696 12792 6702 12804
rect 6546 12724 6552 12776
rect 6604 12764 6610 12776
rect 6932 12773 6960 12804
rect 7834 12792 7840 12804
rect 7892 12792 7898 12844
rect 7926 12792 7932 12844
rect 7984 12832 7990 12844
rect 8093 12835 8151 12841
rect 8093 12832 8105 12835
rect 7984 12804 8105 12832
rect 7984 12792 7990 12804
rect 8093 12801 8105 12804
rect 8139 12801 8151 12835
rect 8093 12795 8151 12801
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12832 9735 12835
rect 9950 12832 9956 12844
rect 9723 12804 9956 12832
rect 9723 12801 9735 12804
rect 9677 12795 9735 12801
rect 9950 12792 9956 12804
rect 10008 12792 10014 12844
rect 10962 12792 10968 12844
rect 11020 12832 11026 12844
rect 11149 12835 11207 12841
rect 11149 12832 11161 12835
rect 11020 12804 11161 12832
rect 11020 12792 11026 12804
rect 11149 12801 11161 12804
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12832 11759 12835
rect 11790 12832 11796 12844
rect 11747 12804 11796 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6604 12736 6837 12764
rect 6604 12724 6610 12736
rect 6825 12733 6837 12736
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 9858 12724 9864 12776
rect 9916 12764 9922 12776
rect 10413 12767 10471 12773
rect 10413 12764 10425 12767
rect 9916 12736 10425 12764
rect 9916 12724 9922 12736
rect 10413 12733 10425 12736
rect 10459 12733 10471 12767
rect 10594 12764 10600 12776
rect 10555 12736 10600 12764
rect 10413 12727 10471 12733
rect 10594 12724 10600 12736
rect 10652 12764 10658 12776
rect 11054 12764 11060 12776
rect 10652 12736 11060 12764
rect 10652 12724 10658 12736
rect 11054 12724 11060 12736
rect 11112 12724 11118 12776
rect 11974 12764 11980 12776
rect 11935 12736 11980 12764
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 6365 12699 6423 12705
rect 6365 12665 6377 12699
rect 6411 12665 6423 12699
rect 6365 12659 6423 12665
rect 9217 12699 9275 12705
rect 9217 12665 9229 12699
rect 9263 12696 9275 12699
rect 9306 12696 9312 12708
rect 9263 12668 9312 12696
rect 9263 12665 9275 12668
rect 9217 12659 9275 12665
rect 9306 12656 9312 12668
rect 9364 12656 9370 12708
rect 9493 12699 9551 12705
rect 9493 12665 9505 12699
rect 9539 12696 9551 12699
rect 9582 12696 9588 12708
rect 9539 12668 9588 12696
rect 9539 12665 9551 12668
rect 9493 12659 9551 12665
rect 9582 12656 9588 12668
rect 9640 12656 9646 12708
rect 12406 12696 12434 12872
rect 13740 12841 13768 12872
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 13726 12835 13784 12841
rect 13726 12801 13738 12835
rect 13772 12801 13784 12835
rect 13832 12832 13860 12940
rect 14277 12937 14289 12971
rect 14323 12968 14335 12971
rect 14550 12968 14556 12980
rect 14323 12940 14556 12968
rect 14323 12937 14335 12940
rect 14277 12931 14335 12937
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 15197 12971 15255 12977
rect 15197 12937 15209 12971
rect 15243 12968 15255 12971
rect 15470 12968 15476 12980
rect 15243 12940 15476 12968
rect 15243 12937 15255 12940
rect 15197 12931 15255 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 16574 12968 16580 12980
rect 15764 12940 16580 12968
rect 13909 12903 13967 12909
rect 13909 12869 13921 12903
rect 13955 12900 13967 12903
rect 14826 12900 14832 12912
rect 13955 12872 14832 12900
rect 13955 12869 13967 12872
rect 13909 12863 13967 12869
rect 14826 12860 14832 12872
rect 14884 12860 14890 12912
rect 13998 12832 14004 12844
rect 13832 12804 14004 12832
rect 13726 12795 13784 12801
rect 12894 12764 12900 12776
rect 12855 12736 12900 12764
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13648 12764 13676 12795
rect 13998 12792 14004 12804
rect 14056 12792 14062 12844
rect 14090 12792 14096 12844
rect 14148 12841 14154 12844
rect 14148 12832 14156 12841
rect 14148 12804 14193 12832
rect 14148 12795 14156 12804
rect 14148 12792 14154 12795
rect 14458 12792 14464 12844
rect 14516 12832 14522 12844
rect 14553 12835 14611 12841
rect 14553 12832 14565 12835
rect 14516 12804 14565 12832
rect 14516 12792 14522 12804
rect 14553 12801 14565 12804
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 14642 12792 14648 12844
rect 14700 12832 14706 12844
rect 14921 12835 14979 12841
rect 14700 12804 14745 12832
rect 14700 12792 14706 12804
rect 14921 12801 14933 12835
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 15059 12835 15117 12841
rect 15059 12801 15071 12835
rect 15105 12832 15117 12835
rect 15657 12835 15715 12841
rect 15105 12804 15240 12832
rect 15105 12801 15117 12804
rect 15059 12795 15117 12801
rect 14476 12764 14504 12792
rect 13648 12736 14504 12764
rect 14182 12696 14188 12708
rect 9784 12668 12434 12696
rect 13280 12668 14188 12696
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12628 5227 12631
rect 5258 12628 5264 12640
rect 5215 12600 5264 12628
rect 5215 12597 5227 12600
rect 5169 12591 5227 12597
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 9784 12628 9812 12668
rect 9456 12600 9812 12628
rect 11885 12631 11943 12637
rect 9456 12588 9462 12600
rect 11885 12597 11897 12631
rect 11931 12628 11943 12631
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 11931 12600 12265 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 12253 12597 12265 12600
rect 12299 12597 12311 12631
rect 12253 12591 12311 12597
rect 12802 12588 12808 12640
rect 12860 12628 12866 12640
rect 13280 12637 13308 12668
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 14936 12696 14964 12795
rect 15102 12696 15108 12708
rect 14936 12668 15108 12696
rect 15102 12656 15108 12668
rect 15160 12656 15166 12708
rect 15212 12696 15240 12804
rect 15657 12801 15669 12835
rect 15703 12832 15715 12835
rect 15764 12832 15792 12940
rect 16574 12928 16580 12940
rect 16632 12968 16638 12980
rect 17862 12968 17868 12980
rect 16632 12940 17868 12968
rect 16632 12928 16638 12940
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 19705 12971 19763 12977
rect 19705 12937 19717 12971
rect 19751 12968 19763 12971
rect 19978 12968 19984 12980
rect 19751 12940 19984 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 20438 12928 20444 12980
rect 20496 12977 20502 12980
rect 20496 12968 20505 12977
rect 21358 12968 21364 12980
rect 20496 12940 20541 12968
rect 21319 12940 21364 12968
rect 20496 12931 20505 12940
rect 20496 12928 20502 12931
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 22554 12968 22560 12980
rect 22515 12940 22560 12968
rect 22554 12928 22560 12940
rect 22612 12928 22618 12980
rect 25038 12928 25044 12980
rect 25096 12968 25102 12980
rect 25593 12971 25651 12977
rect 25593 12968 25605 12971
rect 25096 12940 25605 12968
rect 25096 12928 25102 12940
rect 25593 12937 25605 12940
rect 25639 12937 25651 12971
rect 25866 12968 25872 12980
rect 25827 12940 25872 12968
rect 25593 12931 25651 12937
rect 25866 12928 25872 12940
rect 25924 12928 25930 12980
rect 27890 12928 27896 12980
rect 27948 12968 27954 12980
rect 28353 12971 28411 12977
rect 28353 12968 28365 12971
rect 27948 12940 28365 12968
rect 27948 12928 27954 12940
rect 28353 12937 28365 12940
rect 28399 12937 28411 12971
rect 28353 12931 28411 12937
rect 16942 12860 16948 12912
rect 17000 12900 17006 12912
rect 17405 12903 17463 12909
rect 17405 12900 17417 12903
rect 17000 12872 17417 12900
rect 17000 12860 17006 12872
rect 17405 12869 17417 12872
rect 17451 12869 17463 12903
rect 20070 12900 20076 12912
rect 17405 12863 17463 12869
rect 19168 12872 20076 12900
rect 15703 12804 15792 12832
rect 15841 12835 15899 12841
rect 15703 12801 15715 12804
rect 15657 12795 15715 12801
rect 15841 12801 15853 12835
rect 15887 12832 15899 12835
rect 16206 12832 16212 12844
rect 15887 12804 16212 12832
rect 15887 12801 15899 12804
rect 15841 12795 15899 12801
rect 16206 12792 16212 12804
rect 16264 12792 16270 12844
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12832 16359 12835
rect 16666 12832 16672 12844
rect 16347 12804 16672 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 16666 12792 16672 12804
rect 16724 12832 16730 12844
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16724 12804 16865 12832
rect 16724 12792 16730 12804
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 17770 12792 17776 12844
rect 17828 12832 17834 12844
rect 17865 12835 17923 12841
rect 17865 12832 17877 12835
rect 17828 12804 17877 12832
rect 17828 12792 17834 12804
rect 17865 12801 17877 12804
rect 17911 12801 17923 12835
rect 17865 12795 17923 12801
rect 18693 12835 18751 12841
rect 18693 12801 18705 12835
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 15746 12764 15752 12776
rect 15707 12736 15752 12764
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 16022 12724 16028 12776
rect 16080 12764 16086 12776
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 16080 12736 16957 12764
rect 16080 12724 16086 12736
rect 16945 12733 16957 12736
rect 16991 12733 17003 12767
rect 17954 12764 17960 12776
rect 17915 12736 17960 12764
rect 16945 12727 17003 12733
rect 17954 12724 17960 12736
rect 18012 12764 18018 12776
rect 18708 12764 18736 12795
rect 19058 12792 19064 12844
rect 19116 12832 19122 12844
rect 19168 12841 19196 12872
rect 20070 12860 20076 12872
rect 20128 12860 20134 12912
rect 20346 12900 20352 12912
rect 20307 12872 20352 12900
rect 20346 12860 20352 12872
rect 20404 12860 20410 12912
rect 20533 12903 20591 12909
rect 20533 12869 20545 12903
rect 20579 12900 20591 12903
rect 21913 12903 21971 12909
rect 21913 12900 21925 12903
rect 20579 12872 21925 12900
rect 20579 12869 20591 12872
rect 20533 12863 20591 12869
rect 21913 12869 21925 12872
rect 21959 12869 21971 12903
rect 21913 12863 21971 12869
rect 22465 12903 22523 12909
rect 22465 12869 22477 12903
rect 22511 12900 22523 12903
rect 23198 12900 23204 12912
rect 22511 12872 23204 12900
rect 22511 12869 22523 12872
rect 22465 12863 22523 12869
rect 23198 12860 23204 12872
rect 23256 12860 23262 12912
rect 23750 12900 23756 12912
rect 23400 12872 23756 12900
rect 19153 12835 19211 12841
rect 19153 12832 19165 12835
rect 19116 12804 19165 12832
rect 19116 12792 19122 12804
rect 19153 12801 19165 12804
rect 19199 12801 19211 12835
rect 19153 12795 19211 12801
rect 19334 12792 19340 12844
rect 19392 12832 19398 12844
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 19392 12804 19809 12832
rect 19392 12792 19398 12804
rect 19797 12801 19809 12804
rect 19843 12801 19855 12835
rect 19797 12795 19855 12801
rect 20622 12792 20628 12844
rect 20680 12832 20686 12844
rect 20901 12835 20959 12841
rect 20680 12804 20725 12832
rect 20680 12792 20686 12804
rect 20901 12801 20913 12835
rect 20947 12801 20959 12835
rect 21082 12832 21088 12844
rect 21043 12804 21088 12832
rect 20901 12795 20959 12801
rect 18966 12764 18972 12776
rect 18012 12736 18736 12764
rect 18927 12736 18972 12764
rect 18012 12724 18018 12736
rect 18966 12724 18972 12736
rect 19024 12724 19030 12776
rect 19426 12724 19432 12776
rect 19484 12764 19490 12776
rect 20916 12764 20944 12795
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 21818 12832 21824 12844
rect 21779 12804 21824 12832
rect 21818 12792 21824 12804
rect 21876 12792 21882 12844
rect 22002 12832 22008 12844
rect 21963 12804 22008 12832
rect 22002 12792 22008 12804
rect 22060 12832 22066 12844
rect 23400 12832 23428 12872
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 24486 12909 24492 12912
rect 24480 12900 24492 12909
rect 24447 12872 24492 12900
rect 24480 12863 24492 12872
rect 24486 12860 24492 12863
rect 24544 12860 24550 12912
rect 27154 12860 27160 12912
rect 27212 12909 27218 12912
rect 27212 12903 27276 12909
rect 27212 12869 27230 12903
rect 27264 12869 27276 12903
rect 27212 12863 27276 12869
rect 27212 12860 27218 12863
rect 22060 12804 22416 12832
rect 22060 12792 22066 12804
rect 19484 12736 20944 12764
rect 19484 12724 19490 12736
rect 16669 12699 16727 12705
rect 16669 12696 16681 12699
rect 15212 12668 16681 12696
rect 13265 12631 13323 12637
rect 13265 12628 13277 12631
rect 12860 12600 13277 12628
rect 12860 12588 12866 12600
rect 13265 12597 13277 12600
rect 13311 12597 13323 12631
rect 13265 12591 13323 12597
rect 14090 12588 14096 12640
rect 14148 12628 14154 12640
rect 15212 12628 15240 12668
rect 16669 12665 16681 12668
rect 16715 12665 16727 12699
rect 16669 12659 16727 12665
rect 17405 12699 17463 12705
rect 17405 12665 17417 12699
rect 17451 12696 17463 12699
rect 18138 12696 18144 12708
rect 17451 12668 18144 12696
rect 17451 12665 17463 12668
rect 17405 12659 17463 12665
rect 14148 12600 15240 12628
rect 14148 12588 14154 12600
rect 15930 12588 15936 12640
rect 15988 12628 15994 12640
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15988 12600 16129 12628
rect 15988 12588 15994 12600
rect 16117 12597 16129 12600
rect 16163 12597 16175 12631
rect 16117 12591 16175 12597
rect 16206 12588 16212 12640
rect 16264 12628 16270 12640
rect 17420 12628 17448 12659
rect 18138 12656 18144 12668
rect 18196 12696 18202 12708
rect 18509 12699 18567 12705
rect 18509 12696 18521 12699
rect 18196 12668 18521 12696
rect 18196 12656 18202 12668
rect 18509 12665 18521 12668
rect 18555 12665 18567 12699
rect 18509 12659 18567 12665
rect 19337 12699 19395 12705
rect 19337 12665 19349 12699
rect 19383 12696 19395 12699
rect 20622 12696 20628 12708
rect 19383 12668 20628 12696
rect 19383 12665 19395 12668
rect 19337 12659 19395 12665
rect 20622 12656 20628 12668
rect 20680 12656 20686 12708
rect 21100 12696 21128 12792
rect 22388 12764 22416 12804
rect 23124 12804 23428 12832
rect 22646 12764 22652 12776
rect 22388 12736 22652 12764
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 22925 12767 22983 12773
rect 22925 12733 22937 12767
rect 22971 12764 22983 12767
rect 23124 12764 23152 12804
rect 23474 12792 23480 12844
rect 23532 12832 23538 12844
rect 24213 12835 24271 12841
rect 24213 12832 24225 12835
rect 23532 12804 24225 12832
rect 23532 12792 23538 12804
rect 24213 12801 24225 12804
rect 24259 12801 24271 12835
rect 24213 12795 24271 12801
rect 22971 12736 23152 12764
rect 23201 12767 23259 12773
rect 22971 12733 22983 12736
rect 22925 12727 22983 12733
rect 23201 12733 23213 12767
rect 23247 12764 23259 12767
rect 23566 12764 23572 12776
rect 23247 12736 23572 12764
rect 23247 12733 23259 12736
rect 23201 12727 23259 12733
rect 23566 12724 23572 12736
rect 23624 12724 23630 12776
rect 25222 12724 25228 12776
rect 25280 12764 25286 12776
rect 26142 12764 26148 12776
rect 25280 12736 26148 12764
rect 25280 12724 25286 12736
rect 26142 12724 26148 12736
rect 26200 12764 26206 12776
rect 26973 12767 27031 12773
rect 26973 12764 26985 12767
rect 26200 12736 26985 12764
rect 26200 12724 26206 12736
rect 26973 12733 26985 12736
rect 27019 12733 27031 12767
rect 26973 12727 27031 12733
rect 23658 12696 23664 12708
rect 21100 12668 21496 12696
rect 18046 12628 18052 12640
rect 16264 12600 17448 12628
rect 18007 12600 18052 12628
rect 16264 12588 16270 12600
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 18230 12628 18236 12640
rect 18191 12600 18236 12628
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 20070 12588 20076 12640
rect 20128 12628 20134 12640
rect 20254 12628 20260 12640
rect 20128 12600 20260 12628
rect 20128 12588 20134 12600
rect 20254 12588 20260 12600
rect 20312 12588 20318 12640
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 20901 12631 20959 12637
rect 20901 12628 20913 12631
rect 20772 12600 20913 12628
rect 20772 12588 20778 12600
rect 20901 12597 20913 12600
rect 20947 12597 20959 12631
rect 21468 12628 21496 12668
rect 22066 12668 23664 12696
rect 22066 12628 22094 12668
rect 23658 12656 23664 12668
rect 23716 12656 23722 12708
rect 21468 12600 22094 12628
rect 20901 12591 20959 12597
rect 22738 12588 22744 12640
rect 22796 12628 22802 12640
rect 23106 12628 23112 12640
rect 22796 12600 23112 12628
rect 22796 12588 22802 12600
rect 23106 12588 23112 12600
rect 23164 12628 23170 12640
rect 24854 12628 24860 12640
rect 23164 12600 24860 12628
rect 23164 12588 23170 12600
rect 24854 12588 24860 12600
rect 24912 12588 24918 12640
rect 1104 12538 28888 12560
rect 1104 12486 5582 12538
rect 5634 12486 5646 12538
rect 5698 12486 5710 12538
rect 5762 12486 5774 12538
rect 5826 12486 5838 12538
rect 5890 12486 14846 12538
rect 14898 12486 14910 12538
rect 14962 12486 14974 12538
rect 15026 12486 15038 12538
rect 15090 12486 15102 12538
rect 15154 12486 24110 12538
rect 24162 12486 24174 12538
rect 24226 12486 24238 12538
rect 24290 12486 24302 12538
rect 24354 12486 24366 12538
rect 24418 12486 28888 12538
rect 1104 12464 28888 12486
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9398 12424 9404 12436
rect 8904 12396 9404 12424
rect 8904 12384 8910 12396
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 11204 12396 13645 12424
rect 11204 12384 11210 12396
rect 13633 12393 13645 12396
rect 13679 12424 13691 12427
rect 14182 12424 14188 12436
rect 13679 12396 14188 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 16390 12424 16396 12436
rect 16351 12396 16396 12424
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 18138 12424 18144 12436
rect 18099 12396 18144 12424
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 18506 12384 18512 12436
rect 18564 12424 18570 12436
rect 18785 12427 18843 12433
rect 18785 12424 18797 12427
rect 18564 12396 18797 12424
rect 18564 12384 18570 12396
rect 18785 12393 18797 12396
rect 18831 12393 18843 12427
rect 19426 12424 19432 12436
rect 18785 12387 18843 12393
rect 18984 12396 19432 12424
rect 6546 12356 6552 12368
rect 6459 12328 6552 12356
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 8941 12359 8999 12365
rect 8941 12325 8953 12359
rect 8987 12325 8999 12359
rect 10229 12359 10287 12365
rect 10229 12356 10241 12359
rect 8941 12319 8999 12325
rect 9048 12328 10241 12356
rect 5166 12288 5172 12300
rect 5127 12260 5172 12288
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5258 12180 5264 12232
rect 5316 12220 5322 12232
rect 5425 12223 5483 12229
rect 5425 12220 5437 12223
rect 5316 12192 5437 12220
rect 5316 12180 5322 12192
rect 5425 12189 5437 12192
rect 5471 12189 5483 12223
rect 6564 12220 6592 12316
rect 6638 12248 6644 12300
rect 6696 12288 6702 12300
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 6696 12260 7389 12288
rect 6696 12248 6702 12260
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 8956 12288 8984 12319
rect 7377 12251 7435 12257
rect 8128 12260 8984 12288
rect 8128 12229 8156 12260
rect 8113 12223 8171 12229
rect 6564 12192 7236 12220
rect 5425 12183 5483 12189
rect 7208 12161 7236 12192
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 8202 12180 8208 12232
rect 8260 12220 8266 12232
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 8260 12192 8309 12220
rect 8260 12180 8266 12192
rect 8297 12189 8309 12192
rect 8343 12220 8355 12223
rect 9048 12220 9076 12328
rect 10229 12325 10241 12328
rect 10275 12356 10287 12359
rect 10275 12328 12848 12356
rect 10275 12325 10287 12328
rect 10229 12319 10287 12325
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 9180 12260 9505 12288
rect 9180 12248 9186 12260
rect 9493 12257 9505 12260
rect 9539 12288 9551 12291
rect 10873 12291 10931 12297
rect 10873 12288 10885 12291
rect 9539 12260 10885 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 10873 12257 10885 12260
rect 10919 12288 10931 12291
rect 12066 12288 12072 12300
rect 10919 12260 12072 12288
rect 10919 12257 10931 12260
rect 10873 12251 10931 12257
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 9306 12220 9312 12232
rect 8343 12192 9076 12220
rect 9267 12192 9312 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 11054 12220 11060 12232
rect 11015 12192 11060 12220
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11882 12220 11888 12232
rect 11843 12192 11888 12220
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12220 12035 12223
rect 12023 12192 12480 12220
rect 12023 12189 12035 12192
rect 11977 12183 12035 12189
rect 7193 12155 7251 12161
rect 7193 12121 7205 12155
rect 7239 12152 7251 12155
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 7239 12124 9413 12152
rect 7239 12121 7251 12124
rect 7193 12115 7251 12121
rect 9401 12121 9413 12124
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 9950 12112 9956 12164
rect 10008 12152 10014 12164
rect 10045 12155 10103 12161
rect 10045 12152 10057 12155
rect 10008 12124 10057 12152
rect 10008 12112 10014 12124
rect 10045 12121 10057 12124
rect 10091 12152 10103 12155
rect 12342 12152 12348 12164
rect 10091 12124 12348 12152
rect 10091 12121 10103 12124
rect 10045 12115 10103 12121
rect 12342 12112 12348 12124
rect 12400 12112 12406 12164
rect 1578 12044 1584 12096
rect 1636 12084 1642 12096
rect 1762 12084 1768 12096
rect 1636 12056 1768 12084
rect 1636 12044 1642 12056
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 6638 12044 6644 12096
rect 6696 12084 6702 12096
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 6696 12056 6837 12084
rect 6696 12044 6702 12056
rect 6825 12053 6837 12056
rect 6871 12053 6883 12087
rect 7282 12084 7288 12096
rect 7243 12056 7288 12084
rect 6825 12047 6883 12053
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 7929 12087 7987 12093
rect 7929 12084 7941 12087
rect 7800 12056 7941 12084
rect 7800 12044 7806 12056
rect 7929 12053 7941 12056
rect 7975 12053 7987 12087
rect 7929 12047 7987 12053
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10505 12087 10563 12093
rect 10505 12084 10517 12087
rect 9732 12056 10517 12084
rect 9732 12044 9738 12056
rect 10505 12053 10517 12056
rect 10551 12053 10563 12087
rect 11514 12084 11520 12096
rect 11475 12056 11520 12084
rect 10505 12047 10563 12053
rect 11514 12044 11520 12056
rect 11572 12044 11578 12096
rect 12158 12084 12164 12096
rect 12119 12056 12164 12084
rect 12158 12044 12164 12056
rect 12216 12044 12222 12096
rect 12452 12093 12480 12192
rect 12820 12152 12848 12328
rect 12986 12248 12992 12300
rect 13044 12288 13050 12300
rect 13081 12291 13139 12297
rect 13081 12288 13093 12291
rect 13044 12260 13093 12288
rect 13044 12248 13050 12260
rect 13081 12257 13093 12260
rect 13127 12288 13139 12291
rect 14093 12291 14151 12297
rect 14093 12288 14105 12291
rect 13127 12260 14105 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 14093 12257 14105 12260
rect 14139 12257 14151 12291
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 14093 12251 14151 12257
rect 14476 12260 15301 12288
rect 12894 12180 12900 12232
rect 12952 12220 12958 12232
rect 14274 12220 14280 12232
rect 12952 12192 14141 12220
rect 14235 12192 14280 12220
rect 12952 12180 12958 12192
rect 12820 12124 13492 12152
rect 12437 12087 12495 12093
rect 12437 12053 12449 12087
rect 12483 12053 12495 12087
rect 12437 12047 12495 12053
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 12805 12087 12863 12093
rect 12805 12084 12817 12087
rect 12768 12056 12817 12084
rect 12768 12044 12774 12056
rect 12805 12053 12817 12056
rect 12851 12053 12863 12087
rect 12805 12047 12863 12053
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 13464 12084 13492 12124
rect 13538 12112 13544 12164
rect 13596 12152 13602 12164
rect 14113 12152 14141 12192
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14476 12161 14504 12260
rect 15289 12257 15301 12260
rect 15335 12288 15347 12291
rect 16183 12291 16241 12297
rect 16183 12288 16195 12291
rect 15335 12260 16195 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 16183 12257 16195 12260
rect 16229 12257 16241 12291
rect 16408 12288 16436 12384
rect 16945 12291 17003 12297
rect 16945 12288 16957 12291
rect 16408 12260 16957 12288
rect 16183 12251 16241 12257
rect 16945 12257 16957 12260
rect 16991 12257 17003 12291
rect 16945 12251 17003 12257
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 18141 12291 18199 12297
rect 18141 12288 18153 12291
rect 18104 12260 18153 12288
rect 18104 12248 18110 12260
rect 18141 12257 18153 12260
rect 18187 12257 18199 12291
rect 18141 12251 18199 12257
rect 15838 12220 15844 12232
rect 14568 12192 15844 12220
rect 14461 12155 14519 12161
rect 14461 12152 14473 12155
rect 13596 12124 13641 12152
rect 14113 12124 14473 12152
rect 13596 12112 13602 12124
rect 14461 12121 14473 12124
rect 14507 12121 14519 12155
rect 14461 12115 14519 12121
rect 14568 12084 14596 12192
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 16022 12220 16028 12232
rect 15983 12192 16028 12220
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 16574 12220 16580 12232
rect 16535 12192 16580 12220
rect 16393 12183 16451 12189
rect 14642 12112 14648 12164
rect 14700 12152 14706 12164
rect 15105 12155 15163 12161
rect 15105 12152 15117 12155
rect 14700 12124 15117 12152
rect 14700 12112 14706 12124
rect 15105 12121 15117 12124
rect 15151 12121 15163 12155
rect 16408 12152 16436 12183
rect 16574 12180 16580 12192
rect 16632 12220 16638 12232
rect 16850 12220 16856 12232
rect 16632 12192 16856 12220
rect 16632 12180 16638 12192
rect 16850 12180 16856 12192
rect 16908 12180 16914 12232
rect 17221 12223 17279 12229
rect 17221 12189 17233 12223
rect 17267 12220 17279 12223
rect 17770 12220 17776 12232
rect 17267 12192 17776 12220
rect 17267 12189 17279 12192
rect 17221 12183 17279 12189
rect 17770 12180 17776 12192
rect 17828 12220 17834 12232
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 17828 12192 18092 12220
rect 17828 12180 17834 12192
rect 17954 12152 17960 12164
rect 16408 12124 17960 12152
rect 15105 12115 15163 12121
rect 17954 12112 17960 12124
rect 18012 12112 18018 12164
rect 18064 12161 18092 12192
rect 18156 12192 18337 12220
rect 18049 12155 18107 12161
rect 18049 12121 18061 12155
rect 18095 12121 18107 12155
rect 18049 12115 18107 12121
rect 14734 12084 14740 12096
rect 12952 12056 12997 12084
rect 13464 12056 14596 12084
rect 14695 12056 14740 12084
rect 12952 12044 12958 12056
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15197 12087 15255 12093
rect 15197 12053 15209 12087
rect 15243 12084 15255 12087
rect 17770 12084 17776 12096
rect 15243 12056 17776 12084
rect 15243 12053 15255 12056
rect 15197 12047 15255 12053
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18156 12084 18184 12192
rect 18325 12189 18337 12192
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 17920 12056 18184 12084
rect 18509 12087 18567 12093
rect 17920 12044 17926 12056
rect 18509 12053 18521 12087
rect 18555 12084 18567 12087
rect 18984 12084 19012 12396
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 19886 12384 19892 12436
rect 19944 12424 19950 12436
rect 20254 12424 20260 12436
rect 19944 12396 20260 12424
rect 19944 12384 19950 12396
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 21085 12427 21143 12433
rect 21085 12393 21097 12427
rect 21131 12393 21143 12427
rect 21085 12387 21143 12393
rect 22097 12427 22155 12433
rect 22097 12393 22109 12427
rect 22143 12424 22155 12427
rect 23198 12424 23204 12436
rect 22143 12396 23204 12424
rect 22143 12393 22155 12396
rect 22097 12387 22155 12393
rect 20625 12359 20683 12365
rect 20625 12325 20637 12359
rect 20671 12325 20683 12359
rect 21100 12356 21128 12387
rect 23198 12384 23204 12396
rect 23256 12384 23262 12436
rect 23290 12384 23296 12436
rect 23348 12424 23354 12436
rect 25222 12424 25228 12436
rect 23348 12396 25228 12424
rect 23348 12384 23354 12396
rect 25222 12384 25228 12396
rect 25280 12384 25286 12436
rect 27246 12424 27252 12436
rect 27207 12396 27252 12424
rect 27246 12384 27252 12396
rect 27304 12384 27310 12436
rect 22465 12359 22523 12365
rect 22465 12356 22477 12359
rect 21100 12328 22477 12356
rect 20625 12319 20683 12325
rect 22465 12325 22477 12328
rect 22511 12325 22523 12359
rect 22465 12319 22523 12325
rect 24397 12359 24455 12365
rect 24397 12325 24409 12359
rect 24443 12356 24455 12359
rect 24578 12356 24584 12368
rect 24443 12328 24584 12356
rect 24443 12325 24455 12328
rect 24397 12319 24455 12325
rect 20640 12288 20668 12319
rect 24578 12316 24584 12328
rect 24636 12316 24642 12368
rect 25777 12359 25835 12365
rect 25777 12356 25789 12359
rect 24688 12328 25789 12356
rect 20640 12260 21864 12288
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 19886 12220 19892 12232
rect 19291 12192 19892 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 20622 12180 20628 12232
rect 20680 12220 20686 12232
rect 21726 12220 21732 12232
rect 20680 12192 20944 12220
rect 21687 12192 21732 12220
rect 20680 12180 20686 12192
rect 19512 12155 19570 12161
rect 19512 12121 19524 12155
rect 19558 12152 19570 12155
rect 20714 12152 20720 12164
rect 19558 12124 20720 12152
rect 19558 12121 19570 12124
rect 19512 12115 19570 12121
rect 20714 12112 20720 12124
rect 20772 12112 20778 12164
rect 20916 12161 20944 12192
rect 21726 12180 21732 12192
rect 21784 12180 21790 12232
rect 20901 12155 20959 12161
rect 20901 12121 20913 12155
rect 20947 12121 20959 12155
rect 20901 12115 20959 12121
rect 21117 12155 21175 12161
rect 21117 12121 21129 12155
rect 21163 12152 21175 12155
rect 21163 12124 21588 12152
rect 21163 12121 21175 12124
rect 21117 12115 21175 12121
rect 18555 12056 19012 12084
rect 18555 12053 18567 12056
rect 18509 12047 18567 12053
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 20162 12084 20168 12096
rect 19300 12056 20168 12084
rect 19300 12044 19306 12056
rect 20162 12044 20168 12056
rect 20220 12044 20226 12096
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 21560 12093 21588 12124
rect 21269 12087 21327 12093
rect 21269 12084 21281 12087
rect 21048 12056 21281 12084
rect 21048 12044 21054 12056
rect 21269 12053 21281 12056
rect 21315 12053 21327 12087
rect 21269 12047 21327 12053
rect 21545 12087 21603 12093
rect 21545 12053 21557 12087
rect 21591 12053 21603 12087
rect 21836 12084 21864 12260
rect 22204 12260 23152 12288
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12220 21971 12223
rect 22094 12220 22100 12232
rect 21959 12192 22100 12220
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 22094 12180 22100 12192
rect 22152 12180 22158 12232
rect 22204 12229 22232 12260
rect 22189 12223 22247 12229
rect 22189 12189 22201 12223
rect 22235 12189 22247 12223
rect 22189 12183 22247 12189
rect 22002 12112 22008 12164
rect 22060 12152 22066 12164
rect 22204 12152 22232 12183
rect 22462 12180 22468 12232
rect 22520 12220 22526 12232
rect 22603 12223 22661 12229
rect 22603 12220 22615 12223
rect 22520 12192 22615 12220
rect 22520 12180 22526 12192
rect 22603 12189 22615 12192
rect 22649 12189 22661 12223
rect 22603 12183 22661 12189
rect 22922 12180 22928 12232
rect 22980 12230 22986 12232
rect 22980 12229 23060 12230
rect 23124 12229 23152 12260
rect 23198 12248 23204 12300
rect 23256 12288 23262 12300
rect 24688 12288 24716 12328
rect 25777 12325 25789 12328
rect 25823 12325 25835 12359
rect 25777 12319 25835 12325
rect 23256 12260 23428 12288
rect 23256 12248 23262 12260
rect 23400 12229 23428 12260
rect 23492 12260 24716 12288
rect 22980 12223 23074 12229
rect 22980 12202 23028 12223
rect 22980 12180 22986 12202
rect 23016 12189 23028 12202
rect 23062 12189 23074 12223
rect 23016 12183 23074 12189
rect 23109 12223 23167 12229
rect 23109 12189 23121 12223
rect 23155 12189 23167 12223
rect 23109 12183 23167 12189
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12189 23443 12223
rect 23385 12183 23443 12189
rect 22738 12152 22744 12164
rect 22060 12124 22232 12152
rect 22296 12124 22744 12152
rect 22060 12112 22066 12124
rect 22296 12084 22324 12124
rect 22738 12112 22744 12124
rect 22796 12112 22802 12164
rect 22833 12155 22891 12161
rect 22833 12121 22845 12155
rect 22879 12152 22891 12155
rect 22879 12124 23152 12152
rect 22879 12121 22891 12124
rect 22833 12115 22891 12121
rect 21836 12056 22324 12084
rect 21545 12047 21603 12053
rect 22554 12044 22560 12096
rect 22612 12084 22618 12096
rect 22922 12084 22928 12096
rect 22612 12056 22928 12084
rect 22612 12044 22618 12056
rect 22922 12044 22928 12056
rect 22980 12044 22986 12096
rect 23124 12084 23152 12124
rect 23198 12112 23204 12164
rect 23256 12152 23262 12164
rect 23492 12152 23520 12260
rect 25038 12248 25044 12300
rect 25096 12288 25102 12300
rect 25961 12291 26019 12297
rect 25961 12288 25973 12291
rect 25096 12260 25973 12288
rect 25096 12248 25102 12260
rect 25961 12257 25973 12260
rect 26007 12288 26019 12291
rect 26237 12291 26295 12297
rect 26237 12288 26249 12291
rect 26007 12260 26249 12288
rect 26007 12257 26019 12260
rect 25961 12251 26019 12257
rect 26237 12257 26249 12260
rect 26283 12257 26295 12291
rect 28350 12288 28356 12300
rect 28311 12260 28356 12288
rect 26237 12251 26295 12257
rect 28350 12248 28356 12260
rect 28408 12248 28414 12300
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12220 23627 12223
rect 23750 12220 23756 12232
rect 23615 12192 23756 12220
rect 23615 12189 23627 12192
rect 23569 12183 23627 12189
rect 23750 12180 23756 12192
rect 23808 12180 23814 12232
rect 24670 12220 24676 12232
rect 24631 12192 24676 12220
rect 24670 12180 24676 12192
rect 24728 12180 24734 12232
rect 25682 12220 25688 12232
rect 25643 12192 25688 12220
rect 25682 12180 25688 12192
rect 25740 12180 25746 12232
rect 27062 12220 27068 12232
rect 27023 12192 27068 12220
rect 27062 12180 27068 12192
rect 27120 12180 27126 12232
rect 23256 12124 23520 12152
rect 23256 12112 23262 12124
rect 23658 12112 23664 12164
rect 23716 12152 23722 12164
rect 24397 12155 24455 12161
rect 24397 12152 24409 12155
rect 23716 12124 24409 12152
rect 23716 12112 23722 12124
rect 24397 12121 24409 12124
rect 24443 12152 24455 12155
rect 24486 12152 24492 12164
rect 24443 12124 24492 12152
rect 24443 12121 24455 12124
rect 24397 12115 24455 12121
rect 24486 12112 24492 12124
rect 24544 12112 24550 12164
rect 24762 12112 24768 12164
rect 24820 12152 24826 12164
rect 25041 12155 25099 12161
rect 25041 12152 25053 12155
rect 24820 12124 25053 12152
rect 24820 12112 24826 12124
rect 25041 12121 25053 12124
rect 25087 12121 25099 12155
rect 25222 12152 25228 12164
rect 25183 12124 25228 12152
rect 25041 12115 25099 12121
rect 25222 12112 25228 12124
rect 25280 12112 25286 12164
rect 23477 12087 23535 12093
rect 23477 12084 23489 12087
rect 23124 12056 23489 12084
rect 23477 12053 23489 12056
rect 23523 12084 23535 12087
rect 23566 12084 23572 12096
rect 23523 12056 23572 12084
rect 23523 12053 23535 12056
rect 23477 12047 23535 12053
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 23842 12084 23848 12096
rect 23803 12056 23848 12084
rect 23842 12044 23848 12056
rect 23900 12044 23906 12096
rect 24581 12087 24639 12093
rect 24581 12053 24593 12087
rect 24627 12084 24639 12087
rect 24946 12084 24952 12096
rect 24627 12056 24952 12084
rect 24627 12053 24639 12056
rect 24581 12047 24639 12053
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 25685 12087 25743 12093
rect 25685 12053 25697 12087
rect 25731 12084 25743 12087
rect 26142 12084 26148 12096
rect 25731 12056 26148 12084
rect 25731 12053 25743 12056
rect 25685 12047 25743 12053
rect 26142 12044 26148 12056
rect 26200 12044 26206 12096
rect 1104 11994 28888 12016
rect 1104 11942 10214 11994
rect 10266 11942 10278 11994
rect 10330 11942 10342 11994
rect 10394 11942 10406 11994
rect 10458 11942 10470 11994
rect 10522 11942 19478 11994
rect 19530 11942 19542 11994
rect 19594 11942 19606 11994
rect 19658 11942 19670 11994
rect 19722 11942 19734 11994
rect 19786 11942 28888 11994
rect 1104 11920 28888 11942
rect 5994 11880 6000 11892
rect 5955 11852 6000 11880
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 7926 11880 7932 11892
rect 7887 11852 7932 11880
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 8570 11840 8576 11892
rect 8628 11840 8634 11892
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 11238 11880 11244 11892
rect 10928 11852 11244 11880
rect 10928 11840 10934 11852
rect 11238 11840 11244 11852
rect 11296 11880 11302 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 11296 11852 11529 11880
rect 11296 11840 11302 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 11517 11843 11575 11849
rect 12066 11840 12072 11892
rect 12124 11880 12130 11892
rect 15654 11880 15660 11892
rect 12124 11852 13584 11880
rect 12124 11840 12130 11852
rect 6012 11744 6040 11840
rect 8588 11812 8616 11840
rect 9401 11815 9459 11821
rect 9401 11812 9413 11815
rect 8588 11784 9413 11812
rect 9401 11781 9413 11784
rect 9447 11781 9459 11815
rect 9401 11775 9459 11781
rect 6457 11747 6515 11753
rect 6457 11744 6469 11747
rect 6012 11716 6469 11744
rect 6457 11713 6469 11716
rect 6503 11713 6515 11747
rect 6638 11744 6644 11756
rect 6599 11716 6644 11744
rect 6457 11707 6515 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11744 6883 11747
rect 7101 11747 7159 11753
rect 7101 11744 7113 11747
rect 6871 11716 7113 11744
rect 6871 11713 6883 11716
rect 6825 11707 6883 11713
rect 7101 11713 7113 11716
rect 7147 11713 7159 11747
rect 7742 11744 7748 11756
rect 7703 11716 7748 11744
rect 7101 11707 7159 11713
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 8573 11747 8631 11753
rect 8573 11713 8585 11747
rect 8619 11744 8631 11747
rect 8846 11744 8852 11756
rect 8619 11716 8852 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 10025 11747 10083 11753
rect 10025 11744 10037 11747
rect 9548 11716 10037 11744
rect 9548 11704 9554 11716
rect 10025 11713 10037 11716
rect 10071 11713 10083 11747
rect 10025 11707 10083 11713
rect 12152 11747 12210 11753
rect 12152 11713 12164 11747
rect 12198 11744 12210 11747
rect 12526 11744 12532 11756
rect 12198 11716 12532 11744
rect 12198 11713 12210 11716
rect 12152 11707 12210 11713
rect 12526 11704 12532 11716
rect 12584 11704 12590 11756
rect 13556 11753 13584 11852
rect 14384 11852 15660 11880
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 7340 11648 8677 11676
rect 7340 11636 7346 11648
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 9122 11676 9128 11688
rect 8803 11648 9128 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9306 11636 9312 11688
rect 9364 11676 9370 11688
rect 9769 11679 9827 11685
rect 9769 11676 9781 11679
rect 9364 11648 9781 11676
rect 9364 11636 9370 11648
rect 9769 11645 9781 11648
rect 9815 11645 9827 11679
rect 9769 11639 9827 11645
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 11885 11679 11943 11685
rect 11885 11676 11897 11679
rect 11204 11648 11897 11676
rect 11204 11636 11210 11648
rect 11885 11645 11897 11648
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 12894 11636 12900 11688
rect 12952 11676 12958 11688
rect 13556 11676 13584 11707
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 14277 11747 14335 11753
rect 14277 11744 14289 11747
rect 14240 11716 14289 11744
rect 14240 11704 14246 11716
rect 14277 11713 14289 11716
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 13722 11676 13728 11688
rect 12952 11648 13032 11676
rect 13556 11648 13728 11676
rect 12952 11636 12958 11648
rect 9214 11608 9220 11620
rect 9175 11580 9220 11608
rect 9214 11568 9220 11580
rect 9272 11568 9278 11620
rect 13004 11608 13032 11648
rect 13722 11636 13728 11648
rect 13780 11636 13786 11688
rect 14384 11676 14412 11852
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 16301 11883 16359 11889
rect 16301 11849 16313 11883
rect 16347 11880 16359 11883
rect 16390 11880 16396 11892
rect 16347 11852 16396 11880
rect 16347 11849 16359 11852
rect 16301 11843 16359 11849
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 16666 11880 16672 11892
rect 16627 11852 16672 11880
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 19242 11880 19248 11892
rect 19203 11852 19248 11880
rect 19242 11840 19248 11852
rect 19300 11840 19306 11892
rect 20622 11880 20628 11892
rect 19444 11852 20628 11880
rect 16574 11772 16580 11824
rect 16632 11812 16638 11824
rect 16632 11784 18000 11812
rect 16632 11772 16638 11784
rect 14550 11753 14556 11756
rect 14544 11707 14556 11753
rect 14608 11744 14614 11756
rect 16114 11744 16120 11756
rect 14608 11716 14644 11744
rect 16027 11716 16120 11744
rect 14550 11704 14556 11707
rect 14608 11704 14614 11716
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 16206 11704 16212 11756
rect 16264 11744 16270 11756
rect 16301 11747 16359 11753
rect 16301 11744 16313 11747
rect 16264 11716 16313 11744
rect 16264 11704 16270 11716
rect 16301 11713 16313 11716
rect 16347 11713 16359 11747
rect 16301 11707 16359 11713
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11744 17739 11747
rect 17862 11744 17868 11756
rect 17727 11716 17868 11744
rect 17727 11713 17739 11716
rect 17681 11707 17739 11713
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 17972 11744 18000 11784
rect 18230 11772 18236 11824
rect 18288 11812 18294 11824
rect 18693 11815 18751 11821
rect 18693 11812 18705 11815
rect 18288 11784 18705 11812
rect 18288 11772 18294 11784
rect 18693 11781 18705 11784
rect 18739 11781 18751 11815
rect 18693 11775 18751 11781
rect 18509 11747 18567 11753
rect 18509 11744 18521 11747
rect 17972 11716 18521 11744
rect 18509 11713 18521 11716
rect 18555 11713 18567 11747
rect 18509 11707 18567 11713
rect 19058 11704 19064 11756
rect 19116 11744 19122 11756
rect 19444 11753 19472 11852
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 23842 11880 23848 11892
rect 21928 11852 23848 11880
rect 21928 11821 21956 11852
rect 23842 11840 23848 11852
rect 23900 11840 23906 11892
rect 24489 11883 24547 11889
rect 24489 11849 24501 11883
rect 24535 11880 24547 11883
rect 24854 11880 24860 11892
rect 24535 11852 24860 11880
rect 24535 11849 24547 11852
rect 24489 11843 24547 11849
rect 24854 11840 24860 11852
rect 24912 11840 24918 11892
rect 21913 11815 21971 11821
rect 21913 11812 21925 11815
rect 19904 11784 21925 11812
rect 19429 11747 19487 11753
rect 19429 11744 19441 11747
rect 19116 11716 19441 11744
rect 19116 11704 19122 11716
rect 19429 11713 19441 11716
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 19794 11704 19800 11756
rect 19852 11744 19858 11756
rect 19904 11753 19932 11784
rect 21913 11781 21925 11784
rect 21959 11781 21971 11815
rect 21913 11775 21971 11781
rect 22097 11815 22155 11821
rect 22097 11781 22109 11815
rect 22143 11812 22155 11815
rect 24762 11812 24768 11824
rect 22143 11784 24768 11812
rect 22143 11781 22155 11784
rect 22097 11775 22155 11781
rect 24762 11772 24768 11784
rect 24820 11772 24826 11824
rect 19889 11747 19947 11753
rect 19889 11744 19901 11747
rect 19852 11716 19901 11744
rect 19852 11704 19858 11716
rect 19889 11713 19901 11716
rect 19935 11713 19947 11747
rect 20990 11744 20996 11756
rect 20951 11716 20996 11744
rect 19889 11707 19947 11713
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 21453 11747 21511 11753
rect 21453 11713 21465 11747
rect 21499 11744 21511 11747
rect 21726 11744 21732 11756
rect 21499 11716 21732 11744
rect 21499 11713 21511 11716
rect 21453 11707 21511 11713
rect 21726 11704 21732 11716
rect 21784 11744 21790 11756
rect 22370 11744 22376 11756
rect 21784 11716 22376 11744
rect 21784 11704 21790 11716
rect 22370 11704 22376 11716
rect 22428 11704 22434 11756
rect 22554 11704 22560 11756
rect 22612 11744 22618 11756
rect 22830 11744 22836 11756
rect 22612 11716 22705 11744
rect 22791 11716 22836 11744
rect 22612 11704 22618 11716
rect 22830 11704 22836 11716
rect 22888 11704 22894 11756
rect 23014 11744 23020 11756
rect 22975 11716 23020 11744
rect 23014 11704 23020 11716
rect 23072 11704 23078 11756
rect 23569 11747 23627 11753
rect 23569 11713 23581 11747
rect 23615 11744 23627 11747
rect 23750 11744 23756 11756
rect 23615 11716 23756 11744
rect 23615 11713 23627 11716
rect 23569 11707 23627 11713
rect 23750 11704 23756 11716
rect 23808 11704 23814 11756
rect 24026 11704 24032 11756
rect 24084 11744 24090 11756
rect 24581 11747 24639 11753
rect 24084 11716 24532 11744
rect 24084 11704 24090 11716
rect 14292 11648 14412 11676
rect 16132 11676 16160 11704
rect 17126 11676 17132 11688
rect 16132 11648 17132 11676
rect 13446 11608 13452 11620
rect 13004 11580 13452 11608
rect 7285 11543 7343 11549
rect 7285 11509 7297 11543
rect 7331 11540 7343 11543
rect 7374 11540 7380 11552
rect 7331 11512 7380 11540
rect 7331 11509 7343 11512
rect 7285 11503 7343 11509
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 8202 11540 8208 11552
rect 8163 11512 8208 11540
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11540 11207 11543
rect 11238 11540 11244 11552
rect 11195 11512 11244 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 13280 11549 13308 11580
rect 13446 11568 13452 11580
rect 13504 11568 13510 11620
rect 14292 11608 14320 11648
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 17402 11676 17408 11688
rect 17363 11648 17408 11676
rect 17402 11636 17408 11648
rect 17460 11636 17466 11688
rect 17770 11636 17776 11688
rect 17828 11676 17834 11688
rect 20530 11676 20536 11688
rect 17828 11648 20536 11676
rect 17828 11636 17834 11648
rect 20530 11636 20536 11648
rect 20588 11636 20594 11688
rect 21361 11679 21419 11685
rect 21361 11645 21373 11679
rect 21407 11676 21419 11679
rect 22572 11676 22600 11704
rect 21407 11648 22600 11676
rect 22741 11679 22799 11685
rect 21407 11645 21419 11648
rect 21361 11639 21419 11645
rect 22741 11645 22753 11679
rect 22787 11676 22799 11679
rect 23382 11676 23388 11688
rect 22787 11648 23388 11676
rect 22787 11645 22799 11648
rect 22741 11639 22799 11645
rect 23382 11636 23388 11648
rect 23440 11636 23446 11688
rect 23474 11636 23480 11688
rect 23532 11676 23538 11688
rect 23661 11679 23719 11685
rect 23661 11676 23673 11679
rect 23532 11648 23673 11676
rect 23532 11636 23538 11648
rect 23661 11645 23673 11648
rect 23707 11676 23719 11679
rect 24213 11679 24271 11685
rect 24213 11676 24225 11679
rect 23707 11648 24225 11676
rect 23707 11645 23719 11648
rect 23661 11639 23719 11645
rect 24213 11645 24225 11648
rect 24259 11645 24271 11679
rect 24504 11676 24532 11716
rect 24581 11713 24593 11747
rect 24627 11744 24639 11747
rect 25498 11744 25504 11756
rect 24627 11716 25504 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 25498 11704 25504 11716
rect 25556 11704 25562 11756
rect 25409 11679 25467 11685
rect 25409 11676 25421 11679
rect 24504 11648 25421 11676
rect 24213 11639 24271 11645
rect 25409 11645 25421 11648
rect 25455 11645 25467 11679
rect 25409 11639 25467 11645
rect 25682 11636 25688 11688
rect 25740 11676 25746 11688
rect 25869 11679 25927 11685
rect 25869 11676 25881 11679
rect 25740 11648 25881 11676
rect 25740 11636 25746 11648
rect 25869 11645 25881 11648
rect 25915 11645 25927 11679
rect 25869 11639 25927 11645
rect 13648 11580 14320 11608
rect 13265 11543 13323 11549
rect 13265 11509 13277 11543
rect 13311 11509 13323 11543
rect 13265 11503 13323 11509
rect 13354 11500 13360 11552
rect 13412 11540 13418 11552
rect 13648 11549 13676 11580
rect 16206 11568 16212 11620
rect 16264 11608 16270 11620
rect 16761 11611 16819 11617
rect 16761 11608 16773 11611
rect 16264 11580 16773 11608
rect 16264 11568 16270 11580
rect 16761 11577 16773 11580
rect 16807 11608 16819 11611
rect 18966 11608 18972 11620
rect 16807 11580 18972 11608
rect 16807 11577 16819 11580
rect 16761 11571 16819 11577
rect 18966 11568 18972 11580
rect 19024 11608 19030 11620
rect 19024 11580 19380 11608
rect 19024 11568 19030 11580
rect 13633 11543 13691 11549
rect 13633 11540 13645 11543
rect 13412 11512 13645 11540
rect 13412 11500 13418 11512
rect 13633 11509 13645 11512
rect 13679 11509 13691 11543
rect 13633 11503 13691 11509
rect 14001 11543 14059 11549
rect 14001 11509 14013 11543
rect 14047 11540 14059 11543
rect 14274 11540 14280 11552
rect 14047 11512 14280 11540
rect 14047 11509 14059 11512
rect 14001 11503 14059 11509
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 18782 11540 18788 11552
rect 18743 11512 18788 11540
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 19352 11540 19380 11580
rect 19518 11568 19524 11620
rect 19576 11608 19582 11620
rect 19705 11611 19763 11617
rect 19705 11608 19717 11611
rect 19576 11580 19717 11608
rect 19576 11568 19582 11580
rect 19705 11577 19717 11580
rect 19751 11577 19763 11611
rect 19705 11571 19763 11577
rect 22002 11568 22008 11620
rect 22060 11608 22066 11620
rect 22060 11580 22600 11608
rect 22060 11568 22066 11580
rect 20257 11543 20315 11549
rect 20257 11540 20269 11543
rect 19352 11512 20269 11540
rect 20257 11509 20269 11512
rect 20303 11509 20315 11543
rect 20806 11540 20812 11552
rect 20767 11512 20812 11540
rect 20257 11503 20315 11509
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 22370 11540 22376 11552
rect 22331 11512 22376 11540
rect 22370 11500 22376 11512
rect 22428 11500 22434 11552
rect 22572 11540 22600 11580
rect 22646 11568 22652 11620
rect 22704 11608 22710 11620
rect 23198 11608 23204 11620
rect 22704 11580 23204 11608
rect 22704 11568 22710 11580
rect 23198 11568 23204 11580
rect 23256 11568 23262 11620
rect 24305 11611 24363 11617
rect 24305 11608 24317 11611
rect 23584 11580 24317 11608
rect 23584 11549 23612 11580
rect 24305 11577 24317 11580
rect 24351 11577 24363 11611
rect 24305 11571 24363 11577
rect 23569 11543 23627 11549
rect 23569 11540 23581 11543
rect 22572 11512 23581 11540
rect 23569 11509 23581 11512
rect 23615 11509 23627 11543
rect 23569 11503 23627 11509
rect 23937 11543 23995 11549
rect 23937 11509 23949 11543
rect 23983 11540 23995 11543
rect 24026 11540 24032 11552
rect 23983 11512 24032 11540
rect 23983 11509 23995 11512
rect 23937 11503 23995 11509
rect 24026 11500 24032 11512
rect 24084 11500 24090 11552
rect 24397 11543 24455 11549
rect 24397 11509 24409 11543
rect 24443 11540 24455 11543
rect 24946 11540 24952 11552
rect 24443 11512 24952 11540
rect 24443 11509 24455 11512
rect 24397 11503 24455 11509
rect 24946 11500 24952 11512
rect 25004 11500 25010 11552
rect 1104 11450 28888 11472
rect 1104 11398 5582 11450
rect 5634 11398 5646 11450
rect 5698 11398 5710 11450
rect 5762 11398 5774 11450
rect 5826 11398 5838 11450
rect 5890 11398 14846 11450
rect 14898 11398 14910 11450
rect 14962 11398 14974 11450
rect 15026 11398 15038 11450
rect 15090 11398 15102 11450
rect 15154 11398 24110 11450
rect 24162 11398 24174 11450
rect 24226 11398 24238 11450
rect 24290 11398 24302 11450
rect 24354 11398 24366 11450
rect 24418 11398 28888 11450
rect 1104 11376 28888 11398
rect 6273 11339 6331 11345
rect 6273 11305 6285 11339
rect 6319 11336 6331 11339
rect 7282 11336 7288 11348
rect 6319 11308 7288 11336
rect 6319 11305 6331 11308
rect 6273 11299 6331 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8628 11308 8953 11336
rect 8628 11296 8634 11308
rect 8941 11305 8953 11308
rect 8987 11336 8999 11339
rect 10134 11336 10140 11348
rect 8987 11308 10140 11336
rect 8987 11305 8999 11308
rect 8941 11299 8999 11305
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 12158 11296 12164 11348
rect 12216 11336 12222 11348
rect 12710 11336 12716 11348
rect 12216 11308 12716 11336
rect 12216 11296 12222 11308
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 14458 11336 14464 11348
rect 13504 11308 14464 11336
rect 13504 11296 13510 11308
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 14550 11296 14556 11348
rect 14608 11336 14614 11348
rect 14829 11339 14887 11345
rect 14829 11336 14841 11339
rect 14608 11308 14841 11336
rect 14608 11296 14614 11308
rect 14829 11305 14841 11308
rect 14875 11305 14887 11339
rect 17218 11336 17224 11348
rect 17179 11308 17224 11336
rect 14829 11299 14887 11305
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 17957 11339 18015 11345
rect 17957 11305 17969 11339
rect 18003 11336 18015 11339
rect 18598 11336 18604 11348
rect 18003 11308 18604 11336
rect 18003 11305 18015 11308
rect 17957 11299 18015 11305
rect 18598 11296 18604 11308
rect 18656 11296 18662 11348
rect 22002 11336 22008 11348
rect 20640 11308 21588 11336
rect 21963 11308 22008 11336
rect 9490 11268 9496 11280
rect 9451 11240 9496 11268
rect 9490 11228 9496 11240
rect 9548 11228 9554 11280
rect 10505 11271 10563 11277
rect 10505 11237 10517 11271
rect 10551 11237 10563 11271
rect 10505 11231 10563 11237
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 8294 11200 8300 11212
rect 7699 11172 8300 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 10520 11200 10548 11231
rect 13170 11228 13176 11280
rect 13228 11268 13234 11280
rect 13357 11271 13415 11277
rect 13357 11268 13369 11271
rect 13228 11240 13369 11268
rect 13228 11228 13234 11240
rect 13357 11237 13369 11240
rect 13403 11237 13415 11271
rect 16206 11268 16212 11280
rect 13357 11231 13415 11237
rect 14200 11240 14872 11268
rect 16167 11240 16212 11268
rect 9968 11172 10548 11200
rect 11149 11203 11207 11209
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 7374 11092 7380 11144
rect 7432 11141 7438 11144
rect 7432 11132 7444 11141
rect 8018 11132 8024 11144
rect 7432 11104 7477 11132
rect 7979 11104 8024 11132
rect 7432 11095 7444 11104
rect 7432 11092 7438 11095
rect 8018 11092 8024 11104
rect 8076 11092 8082 11144
rect 8202 11132 8208 11144
rect 8163 11104 8208 11132
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 9968 11141 9996 11172
rect 11149 11169 11161 11203
rect 11195 11200 11207 11203
rect 12434 11200 12440 11212
rect 11195 11172 12440 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 12434 11160 12440 11172
rect 12492 11200 12498 11212
rect 12805 11203 12863 11209
rect 12805 11200 12817 11203
rect 12492 11172 12817 11200
rect 12492 11160 12498 11172
rect 12805 11169 12817 11172
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 14200 11144 14228 11240
rect 14734 11200 14740 11212
rect 14476 11172 14740 11200
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9355 11104 9781 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11101 10103 11135
rect 10870 11132 10876 11144
rect 10831 11104 10876 11132
rect 10045 11095 10103 11101
rect 8389 11067 8447 11073
rect 8389 11033 8401 11067
rect 8435 11064 8447 11067
rect 8754 11064 8760 11076
rect 8435 11036 8760 11064
rect 8435 11033 8447 11036
rect 8389 11027 8447 11033
rect 8754 11024 8760 11036
rect 8812 11024 8818 11076
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 10060 11064 10088 11095
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 11882 11092 11888 11144
rect 11940 11132 11946 11144
rect 12069 11135 12127 11141
rect 12069 11132 12081 11135
rect 11940 11104 12081 11132
rect 11940 11092 11946 11104
rect 12069 11101 12081 11104
rect 12115 11101 12127 11135
rect 12342 11132 12348 11144
rect 12303 11104 12348 11132
rect 12069 11095 12127 11101
rect 9916 11036 10088 11064
rect 12084 11064 12112 11095
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12986 11132 12992 11144
rect 12947 11104 12992 11132
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 13412 11104 13553 11132
rect 13412 11092 13418 11104
rect 13541 11101 13553 11104
rect 13587 11101 13599 11135
rect 14182 11132 14188 11144
rect 14095 11104 14188 11132
rect 13541 11095 13599 11101
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 14274 11092 14280 11144
rect 14332 11132 14338 11144
rect 14476 11141 14504 11172
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 14844 11200 14872 11240
rect 16206 11228 16212 11240
rect 16264 11228 16270 11280
rect 16669 11271 16727 11277
rect 16669 11237 16681 11271
rect 16715 11268 16727 11271
rect 17126 11268 17132 11280
rect 16715 11240 17132 11268
rect 16715 11237 16727 11240
rect 16669 11231 16727 11237
rect 17126 11228 17132 11240
rect 17184 11228 17190 11280
rect 19242 11268 19248 11280
rect 17236 11240 19248 11268
rect 17236 11200 17264 11240
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 19337 11271 19395 11277
rect 19337 11237 19349 11271
rect 19383 11268 19395 11271
rect 20070 11268 20076 11280
rect 19383 11240 20076 11268
rect 19383 11237 19395 11240
rect 19337 11231 19395 11237
rect 20070 11228 20076 11240
rect 20128 11228 20134 11280
rect 14844 11172 17264 11200
rect 17862 11160 17868 11212
rect 17920 11200 17926 11212
rect 18601 11203 18659 11209
rect 17920 11172 18460 11200
rect 17920 11160 17926 11172
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 14332 11104 14381 11132
rect 14332 11092 14338 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11101 14611 11135
rect 15286 11132 15292 11144
rect 15247 11104 15292 11132
rect 14553 11095 14611 11101
rect 13262 11064 13268 11076
rect 12084 11036 13268 11064
rect 9916 11024 9922 11036
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 13722 11024 13728 11076
rect 13780 11064 13786 11076
rect 14568 11064 14596 11095
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 15382 11135 15440 11141
rect 15382 11101 15394 11135
rect 15428 11101 15440 11135
rect 15654 11132 15660 11144
rect 15615 11104 15660 11132
rect 15382 11095 15440 11101
rect 13780 11036 14596 11064
rect 13780 11024 13786 11036
rect 15194 11024 15200 11076
rect 15252 11064 15258 11076
rect 15396 11064 15424 11095
rect 15654 11092 15660 11104
rect 15712 11092 15718 11144
rect 15746 11092 15752 11144
rect 15804 11141 15810 11144
rect 15804 11132 15812 11141
rect 18230 11132 18236 11144
rect 15804 11104 15849 11132
rect 18191 11104 18236 11132
rect 15804 11095 15812 11104
rect 15804 11092 15810 11095
rect 18230 11092 18236 11104
rect 18288 11092 18294 11144
rect 18432 11141 18460 11172
rect 18601 11169 18613 11203
rect 18647 11200 18659 11203
rect 20162 11200 20168 11212
rect 18647 11172 20168 11200
rect 18647 11169 18659 11172
rect 18601 11163 18659 11169
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 18417 11135 18475 11141
rect 18417 11101 18429 11135
rect 18463 11101 18475 11135
rect 18417 11095 18475 11101
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11132 19763 11135
rect 19978 11132 19984 11144
rect 19751 11104 19984 11132
rect 19751 11101 19763 11104
rect 19705 11095 19763 11101
rect 19978 11092 19984 11104
rect 20036 11092 20042 11144
rect 20640 11141 20668 11308
rect 21560 11268 21588 11308
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 22278 11336 22284 11348
rect 22239 11308 22284 11336
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22830 11296 22836 11348
rect 22888 11336 22894 11348
rect 23109 11339 23167 11345
rect 23109 11336 23121 11339
rect 22888 11308 23121 11336
rect 22888 11296 22894 11308
rect 23109 11305 23121 11308
rect 23155 11305 23167 11339
rect 23109 11299 23167 11305
rect 23385 11339 23443 11345
rect 23385 11305 23397 11339
rect 23431 11305 23443 11339
rect 23385 11299 23443 11305
rect 23198 11268 23204 11280
rect 21560 11240 23204 11268
rect 23198 11228 23204 11240
rect 23256 11228 23262 11280
rect 23400 11268 23428 11299
rect 23842 11296 23848 11348
rect 23900 11336 23906 11348
rect 23937 11339 23995 11345
rect 23937 11336 23949 11339
rect 23900 11308 23949 11336
rect 23900 11296 23906 11308
rect 23937 11305 23949 11308
rect 23983 11305 23995 11339
rect 24670 11336 24676 11348
rect 24631 11308 24676 11336
rect 23937 11299 23995 11305
rect 24670 11296 24676 11308
rect 24728 11296 24734 11348
rect 25498 11296 25504 11348
rect 25556 11336 25562 11348
rect 25961 11339 26019 11345
rect 25961 11336 25973 11339
rect 25556 11308 25973 11336
rect 25556 11296 25562 11308
rect 25961 11305 25973 11308
rect 26007 11305 26019 11339
rect 25961 11299 26019 11305
rect 23400 11240 23520 11268
rect 22462 11160 22468 11212
rect 22520 11200 22526 11212
rect 23382 11200 23388 11212
rect 22520 11172 23388 11200
rect 22520 11160 22526 11172
rect 23382 11160 23388 11172
rect 23440 11160 23446 11212
rect 20625 11135 20683 11141
rect 20625 11101 20637 11135
rect 20671 11101 20683 11135
rect 20625 11095 20683 11101
rect 20892 11135 20950 11141
rect 20892 11101 20904 11135
rect 20938 11101 20950 11135
rect 22646 11132 22652 11144
rect 22607 11104 22652 11132
rect 20892 11095 20950 11101
rect 15565 11067 15623 11073
rect 15565 11064 15577 11067
rect 15252 11036 15424 11064
rect 15488 11036 15577 11064
rect 15252 11024 15258 11036
rect 10965 10999 11023 11005
rect 10965 10965 10977 10999
rect 11011 10996 11023 10999
rect 11238 10996 11244 11008
rect 11011 10968 11244 10996
rect 11011 10965 11023 10968
rect 10965 10959 11023 10965
rect 11238 10956 11244 10968
rect 11296 10996 11302 11008
rect 13906 10996 13912 11008
rect 11296 10968 13912 10996
rect 11296 10956 11302 10968
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 14642 10956 14648 11008
rect 14700 10996 14706 11008
rect 15102 10996 15108 11008
rect 14700 10968 15108 10996
rect 14700 10956 14706 10968
rect 15102 10956 15108 10968
rect 15160 10996 15166 11008
rect 15488 10996 15516 11036
rect 15565 11033 15577 11036
rect 15611 11033 15623 11067
rect 17402 11064 17408 11076
rect 17363 11036 17408 11064
rect 15565 11027 15623 11033
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 17589 11067 17647 11073
rect 17589 11033 17601 11067
rect 17635 11064 17647 11067
rect 17954 11064 17960 11076
rect 17635 11036 17960 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 17954 11024 17960 11036
rect 18012 11064 18018 11076
rect 18506 11064 18512 11076
rect 18012 11036 18512 11064
rect 18012 11024 18018 11036
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 18598 11024 18604 11076
rect 18656 11064 18662 11076
rect 19889 11067 19947 11073
rect 18656 11036 19334 11064
rect 18656 11024 18662 11036
rect 15930 10996 15936 11008
rect 15160 10968 15516 10996
rect 15891 10968 15936 10996
rect 15160 10956 15166 10968
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 19306 10996 19334 11036
rect 19889 11033 19901 11067
rect 19935 11064 19947 11067
rect 20073 11067 20131 11073
rect 19935 11036 19969 11064
rect 19935 11033 19947 11036
rect 19889 11027 19947 11033
rect 20073 11033 20085 11067
rect 20119 11064 20131 11067
rect 20714 11064 20720 11076
rect 20119 11036 20720 11064
rect 20119 11033 20131 11036
rect 20073 11027 20131 11033
rect 19904 10996 19932 11027
rect 20714 11024 20720 11036
rect 20772 11024 20778 11076
rect 20806 11024 20812 11076
rect 20864 11064 20870 11076
rect 20916 11064 20944 11095
rect 22646 11092 22652 11104
rect 22704 11092 22710 11144
rect 22833 11135 22891 11141
rect 22833 11101 22845 11135
rect 22879 11132 22891 11135
rect 23106 11132 23112 11144
rect 22879 11104 23112 11132
rect 22879 11101 22891 11104
rect 22833 11095 22891 11101
rect 23106 11092 23112 11104
rect 23164 11092 23170 11144
rect 23290 11092 23296 11144
rect 23348 11132 23354 11144
rect 23492 11132 23520 11240
rect 24026 11228 24032 11280
rect 24084 11268 24090 11280
rect 24765 11271 24823 11277
rect 24765 11268 24777 11271
rect 24084 11240 24777 11268
rect 24084 11228 24090 11240
rect 24765 11237 24777 11240
rect 24811 11237 24823 11271
rect 25516 11268 25544 11296
rect 24765 11231 24823 11237
rect 24872 11240 25544 11268
rect 24581 11203 24639 11209
rect 24581 11169 24593 11203
rect 24627 11200 24639 11203
rect 24670 11200 24676 11212
rect 24627 11172 24676 11200
rect 24627 11169 24639 11172
rect 24581 11163 24639 11169
rect 24670 11160 24676 11172
rect 24728 11160 24734 11212
rect 24872 11141 24900 11240
rect 23348 11104 23520 11132
rect 23661 11135 23719 11141
rect 23348 11092 23354 11104
rect 23661 11101 23673 11135
rect 23707 11132 23719 11135
rect 24857 11135 24915 11141
rect 23707 11104 24440 11132
rect 23707 11101 23719 11104
rect 23661 11095 23719 11101
rect 20864 11036 20944 11064
rect 20864 11024 20870 11036
rect 22278 11024 22284 11076
rect 22336 11064 22342 11076
rect 22741 11067 22799 11073
rect 22741 11064 22753 11067
rect 22336 11036 22753 11064
rect 22336 11024 22342 11036
rect 22741 11033 22753 11036
rect 22787 11064 22799 11067
rect 24026 11064 24032 11076
rect 22787 11036 24032 11064
rect 22787 11033 22799 11036
rect 22741 11027 22799 11033
rect 24026 11024 24032 11036
rect 24084 11024 24090 11076
rect 20254 10996 20260 11008
rect 19306 10968 20260 10996
rect 20254 10956 20260 10968
rect 20312 10956 20318 11008
rect 24412 10996 24440 11104
rect 24857 11101 24869 11135
rect 24903 11101 24915 11135
rect 24857 11095 24915 11101
rect 25222 11092 25228 11144
rect 25280 11132 25286 11144
rect 27341 11135 27399 11141
rect 27341 11132 27353 11135
rect 25280 11104 27353 11132
rect 25280 11092 25286 11104
rect 27341 11101 27353 11104
rect 27387 11101 27399 11135
rect 28350 11132 28356 11144
rect 28311 11104 28356 11132
rect 27341 11095 27399 11101
rect 28350 11092 28356 11104
rect 28408 11092 28414 11144
rect 24486 11024 24492 11076
rect 24544 11064 24550 11076
rect 25133 11067 25191 11073
rect 25133 11064 25145 11067
rect 24544 11036 25145 11064
rect 24544 11024 24550 11036
rect 25133 11033 25145 11036
rect 25179 11033 25191 11067
rect 25314 11064 25320 11076
rect 25275 11036 25320 11064
rect 25133 11027 25191 11033
rect 25314 11024 25320 11036
rect 25372 11024 25378 11076
rect 26142 11024 26148 11076
rect 26200 11064 26206 11076
rect 27074 11067 27132 11073
rect 27074 11064 27086 11067
rect 26200 11036 27086 11064
rect 26200 11024 26206 11036
rect 27074 11033 27086 11036
rect 27120 11033 27132 11067
rect 27074 11027 27132 11033
rect 24854 10996 24860 11008
rect 24412 10968 24860 10996
rect 24854 10956 24860 10968
rect 24912 10956 24918 11008
rect 1104 10906 28888 10928
rect 1104 10854 10214 10906
rect 10266 10854 10278 10906
rect 10330 10854 10342 10906
rect 10394 10854 10406 10906
rect 10458 10854 10470 10906
rect 10522 10854 19478 10906
rect 19530 10854 19542 10906
rect 19594 10854 19606 10906
rect 19658 10854 19670 10906
rect 19722 10854 19734 10906
rect 19786 10854 28888 10906
rect 1104 10832 28888 10854
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 8904 10764 9229 10792
rect 8904 10752 8910 10764
rect 9217 10761 9229 10764
rect 9263 10761 9275 10795
rect 9217 10755 9275 10761
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 10192 10764 10333 10792
rect 10192 10752 10198 10764
rect 10321 10761 10333 10764
rect 10367 10792 10379 10795
rect 16298 10792 16304 10804
rect 10367 10764 16304 10792
rect 10367 10761 10379 10764
rect 10321 10755 10379 10761
rect 8294 10724 8300 10736
rect 7852 10696 8300 10724
rect 7852 10665 7880 10696
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 10870 10684 10876 10736
rect 10928 10724 10934 10736
rect 12084 10733 12112 10764
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 16850 10792 16856 10804
rect 16811 10764 16856 10792
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 23293 10795 23351 10801
rect 23293 10761 23305 10795
rect 23339 10792 23351 10795
rect 23382 10792 23388 10804
rect 23339 10764 23388 10792
rect 23339 10761 23351 10764
rect 23293 10755 23351 10761
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 24486 10792 24492 10804
rect 23952 10764 24492 10792
rect 11057 10727 11115 10733
rect 11057 10724 11069 10727
rect 10928 10696 11069 10724
rect 10928 10684 10934 10696
rect 11057 10693 11069 10696
rect 11103 10693 11115 10727
rect 11057 10687 11115 10693
rect 12069 10727 12127 10733
rect 12069 10693 12081 10727
rect 12115 10693 12127 10727
rect 12069 10687 12127 10693
rect 12253 10727 12311 10733
rect 12253 10693 12265 10727
rect 12299 10724 12311 10727
rect 12986 10724 12992 10736
rect 12299 10696 12992 10724
rect 12299 10693 12311 10696
rect 12253 10687 12311 10693
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 8104 10659 8162 10665
rect 8104 10625 8116 10659
rect 8150 10656 8162 10659
rect 8570 10656 8576 10668
rect 8150 10628 8576 10656
rect 8150 10625 8162 10628
rect 8104 10619 8162 10625
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10656 9827 10659
rect 10042 10656 10048 10668
rect 9815 10628 10048 10656
rect 9815 10625 9827 10628
rect 9769 10619 9827 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 9953 10591 10011 10597
rect 9953 10588 9965 10591
rect 9916 10560 9965 10588
rect 9916 10548 9922 10560
rect 9953 10557 9965 10560
rect 9999 10557 10011 10591
rect 11072 10588 11100 10687
rect 12986 10684 12992 10696
rect 13044 10724 13050 10736
rect 13538 10724 13544 10736
rect 13044 10696 13544 10724
rect 13044 10684 13050 10696
rect 13538 10684 13544 10696
rect 13596 10684 13602 10736
rect 15470 10724 15476 10736
rect 14660 10696 15476 10724
rect 11698 10656 11704 10668
rect 11659 10628 11704 10656
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 12710 10656 12716 10668
rect 12671 10628 12716 10656
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13219 10628 13676 10656
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 12989 10591 13047 10597
rect 11072 10560 12945 10588
rect 9953 10551 10011 10557
rect 10781 10523 10839 10529
rect 10781 10489 10793 10523
rect 10827 10520 10839 10523
rect 12526 10520 12532 10532
rect 10827 10492 12434 10520
rect 12487 10492 12532 10520
rect 10827 10489 10839 10492
rect 10781 10483 10839 10489
rect 9585 10455 9643 10461
rect 9585 10421 9597 10455
rect 9631 10452 9643 10455
rect 9766 10452 9772 10464
rect 9631 10424 9772 10452
rect 9631 10421 9643 10424
rect 9585 10415 9643 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 11422 10412 11428 10464
rect 11480 10452 11486 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 11480 10424 11529 10452
rect 11480 10412 11486 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 12406 10452 12434 10492
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 12710 10452 12716 10464
rect 12406 10424 12716 10452
rect 11517 10415 11575 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 12917 10452 12945 10560
rect 12989 10557 13001 10591
rect 13035 10557 13047 10591
rect 13354 10588 13360 10600
rect 13315 10560 13360 10588
rect 12989 10551 13047 10557
rect 13004 10520 13032 10551
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 13262 10520 13268 10532
rect 13004 10492 13268 10520
rect 13262 10480 13268 10492
rect 13320 10480 13326 10532
rect 13648 10529 13676 10628
rect 13740 10628 14013 10656
rect 13633 10523 13691 10529
rect 13633 10489 13645 10523
rect 13679 10489 13691 10523
rect 13633 10483 13691 10489
rect 13740 10452 13768 10628
rect 14001 10625 14013 10628
rect 14047 10625 14059 10659
rect 14001 10619 14059 10625
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10656 14151 10659
rect 14274 10656 14280 10668
rect 14139 10628 14280 10656
rect 14139 10625 14151 10628
rect 14093 10619 14151 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10588 14243 10591
rect 14660 10588 14688 10696
rect 15470 10684 15476 10696
rect 15528 10724 15534 10736
rect 17497 10727 17555 10733
rect 15528 10696 15976 10724
rect 15528 10684 15534 10696
rect 14734 10616 14740 10668
rect 14792 10656 14798 10668
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14792 10628 15025 10656
rect 14792 10616 14798 10628
rect 15013 10625 15025 10628
rect 15059 10656 15071 10659
rect 15657 10659 15715 10665
rect 15657 10656 15669 10659
rect 15059 10628 15669 10656
rect 15059 10625 15071 10628
rect 15013 10619 15071 10625
rect 14231 10560 14688 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 12917 10424 13768 10452
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 15378 10452 15384 10464
rect 15335 10424 15384 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 15488 10452 15516 10628
rect 15657 10625 15669 10628
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 15746 10588 15752 10600
rect 15707 10560 15752 10588
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 15948 10597 15976 10696
rect 17497 10693 17509 10727
rect 17543 10724 17555 10727
rect 18598 10724 18604 10736
rect 17543 10696 18604 10724
rect 17543 10693 17555 10696
rect 17497 10687 17555 10693
rect 18598 10684 18604 10696
rect 18656 10684 18662 10736
rect 22180 10727 22238 10733
rect 22180 10693 22192 10727
rect 22226 10724 22238 10727
rect 22370 10724 22376 10736
rect 22226 10696 22376 10724
rect 22226 10693 22238 10696
rect 22180 10687 22238 10693
rect 22370 10684 22376 10696
rect 22428 10684 22434 10736
rect 16669 10659 16727 10665
rect 16669 10625 16681 10659
rect 16715 10625 16727 10659
rect 17678 10656 17684 10668
rect 17639 10628 17684 10656
rect 16669 10619 16727 10625
rect 15933 10591 15991 10597
rect 15933 10557 15945 10591
rect 15979 10557 15991 10591
rect 15933 10551 15991 10557
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 16684 10520 16712 10619
rect 17678 10616 17684 10628
rect 17736 10616 17742 10668
rect 19058 10656 19064 10668
rect 19116 10665 19122 10668
rect 19028 10628 19064 10656
rect 19058 10616 19064 10628
rect 19116 10619 19128 10665
rect 20248 10659 20306 10665
rect 20248 10625 20260 10659
rect 20294 10656 20306 10659
rect 20622 10656 20628 10668
rect 20294 10628 20628 10656
rect 20294 10625 20306 10628
rect 20248 10619 20306 10625
rect 19116 10616 19122 10619
rect 20622 10616 20628 10628
rect 20680 10616 20686 10668
rect 23952 10656 23980 10764
rect 24486 10752 24492 10764
rect 24544 10752 24550 10804
rect 24670 10752 24676 10804
rect 24728 10792 24734 10804
rect 24946 10792 24952 10804
rect 24728 10764 24952 10792
rect 24728 10752 24734 10764
rect 24946 10752 24952 10764
rect 25004 10792 25010 10804
rect 25409 10795 25467 10801
rect 25409 10792 25421 10795
rect 25004 10764 25421 10792
rect 25004 10752 25010 10764
rect 25409 10761 25421 10764
rect 25455 10761 25467 10795
rect 25409 10755 25467 10761
rect 26234 10752 26240 10804
rect 26292 10792 26298 10804
rect 27249 10795 27307 10801
rect 27249 10792 27261 10795
rect 26292 10764 27261 10792
rect 26292 10752 26298 10764
rect 27249 10761 27261 10764
rect 27295 10761 27307 10795
rect 27249 10755 27307 10761
rect 25222 10724 25228 10736
rect 24044 10696 25228 10724
rect 24044 10665 24072 10696
rect 25222 10684 25228 10696
rect 25280 10684 25286 10736
rect 25314 10684 25320 10736
rect 25372 10724 25378 10736
rect 26145 10727 26203 10733
rect 26145 10724 26157 10727
rect 25372 10696 26157 10724
rect 25372 10684 25378 10696
rect 26145 10693 26157 10696
rect 26191 10693 26203 10727
rect 26145 10687 26203 10693
rect 26329 10727 26387 10733
rect 26329 10693 26341 10727
rect 26375 10724 26387 10727
rect 26375 10696 27936 10724
rect 26375 10693 26387 10696
rect 26329 10687 26387 10693
rect 21008 10628 23980 10656
rect 24029 10659 24087 10665
rect 19337 10591 19395 10597
rect 19337 10557 19349 10591
rect 19383 10588 19395 10591
rect 19426 10588 19432 10600
rect 19383 10560 19432 10588
rect 19383 10557 19395 10560
rect 19337 10551 19395 10557
rect 19426 10548 19432 10560
rect 19484 10588 19490 10600
rect 19886 10588 19892 10600
rect 19484 10560 19892 10588
rect 19484 10548 19490 10560
rect 19886 10548 19892 10560
rect 19944 10588 19950 10600
rect 19981 10591 20039 10597
rect 19981 10588 19993 10591
rect 19944 10560 19993 10588
rect 19944 10548 19950 10560
rect 19981 10557 19993 10560
rect 20027 10557 20039 10591
rect 19981 10551 20039 10557
rect 18322 10520 18328 10532
rect 15620 10492 16712 10520
rect 16776 10492 18328 10520
rect 15620 10480 15626 10492
rect 16776 10452 16804 10492
rect 18322 10480 18328 10492
rect 18380 10480 18386 10532
rect 17310 10452 17316 10464
rect 15488 10424 16804 10452
rect 17271 10424 17316 10452
rect 17310 10412 17316 10424
rect 17368 10412 17374 10464
rect 17954 10452 17960 10464
rect 17915 10424 17960 10452
rect 17954 10412 17960 10424
rect 18012 10412 18018 10464
rect 18046 10412 18052 10464
rect 18104 10452 18110 10464
rect 18966 10452 18972 10464
rect 18104 10424 18972 10452
rect 18104 10412 18110 10424
rect 18966 10412 18972 10424
rect 19024 10452 19030 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 19024 10424 19625 10452
rect 19024 10412 19030 10424
rect 19613 10421 19625 10424
rect 19659 10452 19671 10455
rect 21008 10452 21036 10628
rect 24029 10625 24041 10659
rect 24075 10625 24087 10659
rect 24029 10619 24087 10625
rect 24296 10659 24354 10665
rect 24296 10625 24308 10659
rect 24342 10656 24354 10659
rect 24578 10656 24584 10668
rect 24342 10628 24584 10656
rect 24342 10625 24354 10628
rect 24296 10619 24354 10625
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 25774 10616 25780 10668
rect 25832 10656 25838 10668
rect 25961 10659 26019 10665
rect 25961 10656 25973 10659
rect 25832 10628 25973 10656
rect 25832 10616 25838 10628
rect 25961 10625 25973 10628
rect 26007 10625 26019 10659
rect 25961 10619 26019 10625
rect 26786 10616 26792 10668
rect 26844 10656 26850 10668
rect 27908 10665 27936 10696
rect 27341 10659 27399 10665
rect 27341 10656 27353 10659
rect 26844 10628 27353 10656
rect 26844 10616 26850 10628
rect 27341 10625 27353 10628
rect 27387 10625 27399 10659
rect 27341 10619 27399 10625
rect 27893 10659 27951 10665
rect 27893 10625 27905 10659
rect 27939 10625 27951 10659
rect 27893 10619 27951 10625
rect 21913 10591 21971 10597
rect 21913 10557 21925 10591
rect 21959 10557 21971 10591
rect 21913 10551 21971 10557
rect 19659 10424 21036 10452
rect 19659 10421 19671 10424
rect 19613 10415 19671 10421
rect 21266 10412 21272 10464
rect 21324 10452 21330 10464
rect 21361 10455 21419 10461
rect 21361 10452 21373 10455
rect 21324 10424 21373 10452
rect 21324 10412 21330 10424
rect 21361 10421 21373 10424
rect 21407 10421 21419 10455
rect 21928 10452 21956 10551
rect 22094 10452 22100 10464
rect 21928 10424 22100 10452
rect 21361 10415 21419 10421
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 23290 10412 23296 10464
rect 23348 10452 23354 10464
rect 26234 10452 26240 10464
rect 23348 10424 26240 10452
rect 23348 10412 23354 10424
rect 26234 10412 26240 10424
rect 26292 10412 26298 10464
rect 27338 10412 27344 10464
rect 27396 10452 27402 10464
rect 27709 10455 27767 10461
rect 27709 10452 27721 10455
rect 27396 10424 27721 10452
rect 27396 10412 27402 10424
rect 27709 10421 27721 10424
rect 27755 10421 27767 10455
rect 27709 10415 27767 10421
rect 1104 10362 28888 10384
rect 1104 10310 5582 10362
rect 5634 10310 5646 10362
rect 5698 10310 5710 10362
rect 5762 10310 5774 10362
rect 5826 10310 5838 10362
rect 5890 10310 14846 10362
rect 14898 10310 14910 10362
rect 14962 10310 14974 10362
rect 15026 10310 15038 10362
rect 15090 10310 15102 10362
rect 15154 10310 24110 10362
rect 24162 10310 24174 10362
rect 24226 10310 24238 10362
rect 24290 10310 24302 10362
rect 24354 10310 24366 10362
rect 24418 10310 28888 10362
rect 1104 10288 28888 10310
rect 9674 10248 9680 10260
rect 2746 10220 9680 10248
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 2746 10044 2774 10220
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 13078 10248 13084 10260
rect 12575 10220 13084 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 14182 10248 14188 10260
rect 13188 10220 14188 10248
rect 12710 10140 12716 10192
rect 12768 10180 12774 10192
rect 13188 10180 13216 10220
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 14829 10251 14887 10257
rect 14829 10217 14841 10251
rect 14875 10248 14887 10251
rect 15286 10248 15292 10260
rect 14875 10220 15292 10248
rect 14875 10217 14887 10220
rect 14829 10211 14887 10217
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 15562 10248 15568 10260
rect 15523 10220 15568 10248
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 16025 10251 16083 10257
rect 16025 10248 16037 10251
rect 15804 10220 16037 10248
rect 15804 10208 15810 10220
rect 16025 10217 16037 10220
rect 16071 10217 16083 10251
rect 17678 10248 17684 10260
rect 17639 10220 17684 10248
rect 16025 10211 16083 10217
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 18877 10251 18935 10257
rect 18877 10217 18889 10251
rect 18923 10248 18935 10251
rect 19058 10248 19064 10260
rect 18923 10220 19064 10248
rect 18923 10217 18935 10220
rect 18877 10211 18935 10217
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 19613 10251 19671 10257
rect 19613 10217 19625 10251
rect 19659 10248 19671 10251
rect 19978 10248 19984 10260
rect 19659 10220 19984 10248
rect 19659 10217 19671 10220
rect 19613 10211 19671 10217
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 20622 10248 20628 10260
rect 20583 10220 20628 10248
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 25774 10248 25780 10260
rect 25735 10220 25780 10248
rect 25774 10208 25780 10220
rect 25832 10208 25838 10260
rect 12768 10152 13216 10180
rect 12768 10140 12774 10152
rect 13262 10140 13268 10192
rect 13320 10180 13326 10192
rect 19426 10180 19432 10192
rect 13320 10152 15240 10180
rect 13320 10140 13326 10152
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10112 8263 10115
rect 8294 10112 8300 10124
rect 8251 10084 8300 10112
rect 8251 10081 8263 10084
rect 8205 10075 8263 10081
rect 8294 10072 8300 10084
rect 8352 10112 8358 10124
rect 8938 10112 8944 10124
rect 8352 10084 8944 10112
rect 8352 10072 8358 10084
rect 8938 10072 8944 10084
rect 8996 10112 9002 10124
rect 9306 10112 9312 10124
rect 8996 10084 9312 10112
rect 8996 10072 9002 10084
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 11146 10112 11152 10124
rect 11107 10084 11152 10112
rect 11146 10072 11152 10084
rect 11204 10072 11210 10124
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 13357 10115 13415 10121
rect 13357 10112 13369 10115
rect 12492 10084 13369 10112
rect 12492 10072 12498 10084
rect 13357 10081 13369 10084
rect 13403 10081 13415 10115
rect 13357 10075 13415 10081
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 15212 10121 15240 10152
rect 17420 10152 19432 10180
rect 15197 10115 15255 10121
rect 14056 10084 14596 10112
rect 14056 10072 14062 10084
rect 1903 10016 2774 10044
rect 8389 10047 8447 10053
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 9214 10044 9220 10056
rect 8435 10016 9220 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 11422 10053 11428 10056
rect 11416 10044 11428 10053
rect 11383 10016 11428 10044
rect 11416 10007 11428 10016
rect 11422 10004 11428 10007
rect 11480 10004 11486 10056
rect 11532 10016 13032 10044
rect 1578 9936 1584 9988
rect 1636 9976 1642 9988
rect 9582 9985 9588 9988
rect 1673 9979 1731 9985
rect 1673 9976 1685 9979
rect 1636 9948 1685 9976
rect 1636 9936 1642 9948
rect 1673 9945 1685 9948
rect 1719 9976 1731 9979
rect 2133 9979 2191 9985
rect 2133 9976 2145 9979
rect 1719 9948 2145 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 2133 9945 2145 9948
rect 2179 9945 2191 9979
rect 2133 9939 2191 9945
rect 9576 9939 9588 9985
rect 9640 9976 9646 9988
rect 9640 9948 9676 9976
rect 9582 9936 9588 9939
rect 9640 9936 9646 9948
rect 10686 9908 10692 9920
rect 10599 9880 10692 9908
rect 10686 9868 10692 9880
rect 10744 9908 10750 9920
rect 11532 9908 11560 10016
rect 11790 9936 11796 9988
rect 11848 9976 11854 9988
rect 13004 9976 13032 10016
rect 13078 10004 13084 10056
rect 13136 10044 13142 10056
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 13136 10016 13277 10044
rect 13136 10004 13142 10016
rect 13265 10013 13277 10016
rect 13311 10044 13323 10047
rect 13814 10044 13820 10056
rect 13311 10016 13820 10044
rect 13311 10013 13323 10016
rect 13265 10007 13323 10013
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 14182 10044 14188 10056
rect 14143 10016 14188 10044
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14274 10004 14280 10056
rect 14332 10044 14338 10056
rect 14568 10053 14596 10084
rect 15197 10081 15209 10115
rect 15243 10112 15255 10115
rect 16206 10112 16212 10124
rect 15243 10084 16212 10112
rect 15243 10081 15255 10084
rect 15197 10075 15255 10081
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 17420 10121 17448 10152
rect 19426 10140 19432 10152
rect 19484 10140 19490 10192
rect 21266 10180 21272 10192
rect 20088 10152 21272 10180
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 18230 10072 18236 10124
rect 18288 10112 18294 10124
rect 18325 10115 18383 10121
rect 18325 10112 18337 10115
rect 18288 10084 18337 10112
rect 18288 10072 18294 10084
rect 18325 10081 18337 10084
rect 18371 10112 18383 10115
rect 18782 10112 18788 10124
rect 18371 10084 18788 10112
rect 18371 10081 18383 10084
rect 18325 10075 18383 10081
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 20088 10121 20116 10152
rect 21266 10140 21272 10152
rect 21324 10140 21330 10192
rect 23566 10140 23572 10192
rect 23624 10180 23630 10192
rect 26786 10180 26792 10192
rect 23624 10152 26792 10180
rect 23624 10140 23630 10152
rect 20073 10115 20131 10121
rect 20073 10081 20085 10115
rect 20119 10081 20131 10115
rect 20073 10075 20131 10081
rect 20162 10072 20168 10124
rect 20220 10112 20226 10124
rect 21545 10115 21603 10121
rect 21545 10112 21557 10115
rect 20220 10084 20265 10112
rect 20548 10084 21557 10112
rect 20220 10072 20226 10084
rect 14553 10047 14611 10053
rect 14332 10016 14377 10044
rect 14332 10004 14338 10016
rect 14553 10013 14565 10047
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 14691 10047 14749 10053
rect 14691 10013 14703 10047
rect 14737 10044 14749 10047
rect 15378 10044 15384 10056
rect 14737 10016 15148 10044
rect 15339 10016 15384 10044
rect 14737 10013 14749 10016
rect 14691 10007 14749 10013
rect 11848 9948 12848 9976
rect 13004 9948 13769 9976
rect 11848 9936 11854 9948
rect 12820 9917 12848 9948
rect 10744 9880 11560 9908
rect 12805 9911 12863 9917
rect 10744 9868 10750 9880
rect 12805 9877 12817 9911
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 13173 9911 13231 9917
rect 13173 9877 13185 9911
rect 13219 9908 13231 9911
rect 13446 9908 13452 9920
rect 13219 9880 13452 9908
rect 13219 9877 13231 9880
rect 13173 9871 13231 9877
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 13741 9908 13769 9948
rect 13906 9936 13912 9988
rect 13964 9976 13970 9988
rect 14461 9979 14519 9985
rect 14461 9976 14473 9979
rect 13964 9948 14473 9976
rect 13964 9936 13970 9948
rect 14461 9945 14473 9948
rect 14507 9945 14519 9979
rect 15120 9976 15148 10016
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17138 10047 17196 10053
rect 17138 10044 17150 10047
rect 16908 10016 17150 10044
rect 16908 10004 16914 10016
rect 17138 10013 17150 10016
rect 17184 10013 17196 10047
rect 17138 10007 17196 10013
rect 17310 10004 17316 10056
rect 17368 10044 17374 10056
rect 18693 10047 18751 10053
rect 18693 10044 18705 10047
rect 17368 10016 18705 10044
rect 17368 10004 17374 10016
rect 18693 10013 18705 10016
rect 18739 10013 18751 10047
rect 19978 10044 19984 10056
rect 19939 10016 19984 10044
rect 18693 10007 18751 10013
rect 19978 10004 19984 10016
rect 20036 10044 20042 10056
rect 20548 10044 20576 10084
rect 21545 10081 21557 10084
rect 21591 10081 21603 10115
rect 21545 10075 21603 10081
rect 22741 10115 22799 10121
rect 22741 10081 22753 10115
rect 22787 10112 22799 10115
rect 23290 10112 23296 10124
rect 22787 10084 23296 10112
rect 22787 10081 22799 10084
rect 22741 10075 22799 10081
rect 23290 10072 23296 10084
rect 23348 10072 23354 10124
rect 24670 10072 24676 10124
rect 24728 10112 24734 10124
rect 26344 10121 26372 10152
rect 26786 10140 26792 10152
rect 26844 10140 26850 10192
rect 26329 10115 26387 10121
rect 24728 10084 25452 10112
rect 24728 10072 24734 10084
rect 20036 10016 20576 10044
rect 20036 10004 20042 10016
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 20809 10047 20867 10053
rect 20809 10044 20821 10047
rect 20772 10016 20821 10044
rect 20772 10004 20778 10016
rect 20809 10013 20821 10016
rect 20855 10013 20867 10047
rect 20809 10007 20867 10013
rect 21085 10047 21143 10053
rect 21085 10013 21097 10047
rect 21131 10013 21143 10047
rect 21085 10007 21143 10013
rect 23753 10047 23811 10053
rect 23753 10013 23765 10047
rect 23799 10044 23811 10047
rect 23934 10044 23940 10056
rect 23799 10016 23940 10044
rect 23799 10013 23811 10016
rect 23753 10007 23811 10013
rect 17954 9976 17960 9988
rect 15120 9948 17960 9976
rect 14461 9939 14519 9945
rect 17954 9936 17960 9948
rect 18012 9976 18018 9988
rect 18141 9979 18199 9985
rect 18141 9976 18153 9979
rect 18012 9948 18153 9976
rect 18012 9936 18018 9948
rect 18141 9945 18153 9948
rect 18187 9945 18199 9979
rect 18141 9939 18199 9945
rect 18414 9936 18420 9988
rect 18472 9976 18478 9988
rect 21100 9976 21128 10007
rect 23934 10004 23940 10016
rect 23992 10044 23998 10056
rect 25130 10044 25136 10056
rect 23992 10016 25136 10044
rect 23992 10004 23998 10016
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 25314 10044 25320 10056
rect 25275 10016 25320 10044
rect 25314 10004 25320 10016
rect 25372 10004 25378 10056
rect 25424 10044 25452 10084
rect 26329 10081 26341 10115
rect 26375 10081 26387 10115
rect 26329 10075 26387 10081
rect 26789 10047 26847 10053
rect 26789 10044 26801 10047
rect 25424 10016 26801 10044
rect 26789 10013 26801 10016
rect 26835 10013 26847 10047
rect 26789 10007 26847 10013
rect 27056 10047 27114 10053
rect 27056 10013 27068 10047
rect 27102 10044 27114 10047
rect 27338 10044 27344 10056
rect 27102 10016 27344 10044
rect 27102 10013 27114 10016
rect 27056 10007 27114 10013
rect 27338 10004 27344 10016
rect 27396 10004 27402 10056
rect 23566 9976 23572 9988
rect 18472 9948 21128 9976
rect 23527 9948 23572 9976
rect 18472 9936 18478 9948
rect 23566 9936 23572 9948
rect 23624 9936 23630 9988
rect 24026 9936 24032 9988
rect 24084 9976 24090 9988
rect 24673 9979 24731 9985
rect 24673 9976 24685 9979
rect 24084 9948 24685 9976
rect 24084 9936 24090 9948
rect 24673 9945 24685 9948
rect 24719 9945 24731 9979
rect 24854 9976 24860 9988
rect 24815 9948 24860 9976
rect 24673 9939 24731 9945
rect 24854 9936 24860 9948
rect 24912 9936 24918 9988
rect 26145 9979 26203 9985
rect 26145 9945 26157 9979
rect 26191 9976 26203 9979
rect 26191 9948 28120 9976
rect 26191 9945 26203 9948
rect 26145 9939 26203 9945
rect 28092 9920 28120 9948
rect 14642 9908 14648 9920
rect 13741 9880 14648 9908
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 18046 9908 18052 9920
rect 18007 9880 18052 9908
rect 18046 9868 18052 9880
rect 18104 9868 18110 9920
rect 19337 9911 19395 9917
rect 19337 9877 19349 9911
rect 19383 9908 19395 9911
rect 19886 9908 19892 9920
rect 19383 9880 19892 9908
rect 19383 9877 19395 9880
rect 19337 9871 19395 9877
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 21174 9868 21180 9920
rect 21232 9908 21238 9920
rect 21269 9911 21327 9917
rect 21269 9908 21281 9911
rect 21232 9880 21281 9908
rect 21232 9868 21238 9880
rect 21269 9877 21281 9880
rect 21315 9877 21327 9911
rect 21269 9871 21327 9877
rect 22097 9911 22155 9917
rect 22097 9877 22109 9911
rect 22143 9908 22155 9911
rect 22186 9908 22192 9920
rect 22143 9880 22192 9908
rect 22143 9877 22155 9880
rect 22097 9871 22155 9877
rect 22186 9868 22192 9880
rect 22244 9868 22250 9920
rect 22462 9908 22468 9920
rect 22423 9880 22468 9908
rect 22462 9868 22468 9880
rect 22520 9868 22526 9920
rect 22557 9911 22615 9917
rect 22557 9877 22569 9911
rect 22603 9908 22615 9911
rect 23474 9908 23480 9920
rect 22603 9880 23480 9908
rect 22603 9877 22615 9880
rect 22557 9871 22615 9877
rect 23474 9868 23480 9880
rect 23532 9868 23538 9920
rect 23842 9868 23848 9920
rect 23900 9908 23906 9920
rect 23937 9911 23995 9917
rect 23937 9908 23949 9911
rect 23900 9880 23949 9908
rect 23900 9868 23906 9880
rect 23937 9877 23949 9880
rect 23983 9877 23995 9911
rect 25498 9908 25504 9920
rect 25459 9880 25504 9908
rect 23937 9871 23995 9877
rect 25498 9868 25504 9880
rect 25556 9868 25562 9920
rect 26237 9911 26295 9917
rect 26237 9877 26249 9911
rect 26283 9908 26295 9911
rect 26510 9908 26516 9920
rect 26283 9880 26516 9908
rect 26283 9877 26295 9880
rect 26237 9871 26295 9877
rect 26510 9868 26516 9880
rect 26568 9868 26574 9920
rect 28074 9868 28080 9920
rect 28132 9908 28138 9920
rect 28169 9911 28227 9917
rect 28169 9908 28181 9911
rect 28132 9880 28181 9908
rect 28132 9868 28138 9880
rect 28169 9877 28181 9880
rect 28215 9877 28227 9911
rect 28169 9871 28227 9877
rect 1104 9818 28888 9840
rect 1104 9766 10214 9818
rect 10266 9766 10278 9818
rect 10330 9766 10342 9818
rect 10394 9766 10406 9818
rect 10458 9766 10470 9818
rect 10522 9766 19478 9818
rect 19530 9766 19542 9818
rect 19594 9766 19606 9818
rect 19658 9766 19670 9818
rect 19722 9766 19734 9818
rect 19786 9766 28888 9818
rect 1104 9744 28888 9766
rect 8570 9704 8576 9716
rect 8531 9676 8576 9704
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 9582 9704 9588 9716
rect 9543 9676 9588 9704
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 10042 9704 10048 9716
rect 10003 9676 10048 9704
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 10505 9707 10563 9713
rect 10505 9673 10517 9707
rect 10551 9704 10563 9707
rect 10686 9704 10692 9716
rect 10551 9676 10692 9704
rect 10551 9673 10563 9676
rect 10505 9667 10563 9673
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 11517 9707 11575 9713
rect 11517 9673 11529 9707
rect 11563 9704 11575 9707
rect 11698 9704 11704 9716
rect 11563 9676 11704 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 11974 9664 11980 9716
rect 12032 9704 12038 9716
rect 12161 9707 12219 9713
rect 12161 9704 12173 9707
rect 12032 9676 12173 9704
rect 12032 9664 12038 9676
rect 12161 9673 12173 9676
rect 12207 9673 12219 9707
rect 14274 9704 14280 9716
rect 14235 9676 14280 9704
rect 12161 9667 12219 9673
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 15657 9707 15715 9713
rect 15657 9673 15669 9707
rect 15703 9673 15715 9707
rect 19061 9707 19119 9713
rect 19061 9704 19073 9707
rect 15657 9667 15715 9673
rect 18800 9676 19073 9704
rect 11238 9636 11244 9648
rect 10704 9608 11244 9636
rect 8754 9568 8760 9580
rect 8715 9540 8760 9568
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 9766 9568 9772 9580
rect 9727 9540 9772 9568
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10428 9432 10456 9531
rect 10704 9509 10732 9608
rect 11238 9596 11244 9608
rect 11296 9636 11302 9648
rect 12434 9636 12440 9648
rect 11296 9608 12440 9636
rect 11296 9596 11302 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 12621 9639 12679 9645
rect 12621 9605 12633 9639
rect 12667 9636 12679 9639
rect 12710 9636 12716 9648
rect 12667 9608 12716 9636
rect 12667 9605 12679 9608
rect 12621 9599 12679 9605
rect 12710 9596 12716 9608
rect 12768 9596 12774 9648
rect 13170 9645 13176 9648
rect 13164 9636 13176 9645
rect 13131 9608 13176 9636
rect 13164 9599 13176 9608
rect 13170 9596 13176 9599
rect 13228 9596 13234 9648
rect 13262 9596 13268 9648
rect 13320 9596 13326 9648
rect 13446 9596 13452 9648
rect 13504 9636 13510 9648
rect 14553 9639 14611 9645
rect 14553 9636 14565 9639
rect 13504 9608 14565 9636
rect 13504 9596 13510 9608
rect 14553 9605 14565 9608
rect 14599 9605 14611 9639
rect 14553 9599 14611 9605
rect 15289 9639 15347 9645
rect 15289 9605 15301 9639
rect 15335 9636 15347 9639
rect 15562 9636 15568 9648
rect 15335 9608 15568 9636
rect 15335 9605 15347 9608
rect 15289 9599 15347 9605
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9568 11759 9571
rect 11790 9568 11796 9580
rect 11747 9540 11796 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9568 11943 9571
rect 13280 9568 13308 9596
rect 11931 9540 13308 9568
rect 14568 9568 14596 9599
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 15672 9568 15700 9667
rect 15746 9596 15752 9648
rect 15804 9636 15810 9648
rect 17954 9636 17960 9648
rect 15804 9608 17960 9636
rect 15804 9596 15810 9608
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 18800 9645 18828 9676
rect 19061 9673 19073 9676
rect 19107 9673 19119 9707
rect 19061 9667 19119 9673
rect 22462 9664 22468 9716
rect 22520 9704 22526 9716
rect 22833 9707 22891 9713
rect 22833 9704 22845 9707
rect 22520 9676 22845 9704
rect 22520 9664 22526 9676
rect 22833 9673 22845 9676
rect 22879 9673 22891 9707
rect 22833 9667 22891 9673
rect 18049 9639 18107 9645
rect 18049 9605 18061 9639
rect 18095 9636 18107 9639
rect 18785 9639 18843 9645
rect 18095 9608 18736 9636
rect 18095 9605 18107 9608
rect 18049 9599 18107 9605
rect 16117 9571 16175 9577
rect 16117 9568 16129 9571
rect 14568 9540 15332 9568
rect 15672 9540 16129 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9469 10747 9503
rect 12894 9500 12900 9512
rect 12855 9472 12900 9500
rect 10689 9463 10747 9469
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9469 15071 9503
rect 15194 9500 15200 9512
rect 15155 9472 15200 9500
rect 15013 9463 15071 9469
rect 10778 9432 10784 9444
rect 10428 9404 10784 9432
rect 9214 9364 9220 9376
rect 9175 9336 9220 9364
rect 9214 9324 9220 9336
rect 9272 9364 9278 9376
rect 10428 9364 10456 9404
rect 10778 9392 10784 9404
rect 10836 9432 10842 9444
rect 12710 9432 12716 9444
rect 10836 9404 12716 9432
rect 10836 9392 10842 9404
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 15028 9432 15056 9463
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 15304 9500 15332 9540
rect 16117 9537 16129 9540
rect 16163 9537 16175 9571
rect 16117 9531 16175 9537
rect 16206 9528 16212 9580
rect 16264 9568 16270 9580
rect 16264 9540 16309 9568
rect 16264 9528 16270 9540
rect 17034 9528 17040 9580
rect 17092 9568 17098 9580
rect 17313 9571 17371 9577
rect 17313 9568 17325 9571
rect 17092 9540 17325 9568
rect 17092 9528 17098 9540
rect 17313 9537 17325 9540
rect 17359 9537 17371 9571
rect 18414 9568 18420 9580
rect 18375 9540 18420 9568
rect 17313 9531 17371 9537
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 18598 9568 18604 9580
rect 18559 9540 18604 9568
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 18708 9566 18736 9608
rect 18785 9605 18797 9639
rect 18831 9605 18843 9639
rect 18785 9599 18843 9605
rect 20070 9596 20076 9648
rect 20128 9636 20134 9648
rect 25400 9639 25458 9645
rect 20128 9608 25176 9636
rect 20128 9596 20134 9608
rect 19334 9568 19340 9580
rect 18892 9566 19340 9568
rect 18708 9540 19340 9566
rect 18708 9538 18920 9540
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9568 19487 9571
rect 19886 9568 19892 9580
rect 19475 9540 19892 9568
rect 19475 9537 19487 9540
rect 19429 9531 19487 9537
rect 15304 9472 18736 9500
rect 15470 9432 15476 9444
rect 15028 9404 15476 9432
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 17862 9432 17868 9444
rect 17823 9404 17868 9432
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 18708 9432 18736 9472
rect 19444 9432 19472 9531
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 21174 9528 21180 9580
rect 21232 9577 21238 9580
rect 21232 9568 21244 9577
rect 21453 9571 21511 9577
rect 21232 9540 21277 9568
rect 21232 9531 21244 9540
rect 21453 9537 21465 9571
rect 21499 9568 21511 9571
rect 22094 9568 22100 9580
rect 21499 9540 22100 9568
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 21232 9528 21238 9531
rect 22094 9528 22100 9540
rect 22152 9528 22158 9580
rect 22278 9568 22284 9580
rect 22204 9540 22284 9568
rect 19521 9503 19579 9509
rect 19521 9469 19533 9503
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 18708 9404 19472 9432
rect 19536 9432 19564 9463
rect 19702 9460 19708 9512
rect 19760 9500 19766 9512
rect 20162 9500 20168 9512
rect 19760 9472 20168 9500
rect 19760 9460 19766 9472
rect 20162 9460 20168 9472
rect 20220 9460 20226 9512
rect 22204 9509 22232 9540
rect 22278 9528 22284 9540
rect 22336 9528 22342 9580
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9537 22523 9571
rect 22465 9531 22523 9537
rect 22189 9503 22247 9509
rect 22189 9469 22201 9503
rect 22235 9469 22247 9503
rect 22370 9500 22376 9512
rect 22331 9472 22376 9500
rect 22189 9463 22247 9469
rect 22370 9460 22376 9472
rect 22428 9460 22434 9512
rect 19536 9404 20116 9432
rect 9272 9336 10456 9364
rect 9272 9324 9278 9336
rect 13538 9324 13544 9376
rect 13596 9364 13602 9376
rect 15933 9367 15991 9373
rect 15933 9364 15945 9367
rect 13596 9336 15945 9364
rect 13596 9324 13602 9336
rect 15933 9333 15945 9336
rect 15979 9333 15991 9367
rect 16666 9364 16672 9376
rect 16627 9336 16672 9364
rect 15933 9327 15991 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 20088 9373 20116 9404
rect 20073 9367 20131 9373
rect 20073 9333 20085 9367
rect 20119 9364 20131 9367
rect 22480 9364 22508 9531
rect 24026 9528 24032 9580
rect 24084 9568 24090 9580
rect 24590 9571 24648 9577
rect 24590 9568 24602 9571
rect 24084 9540 24602 9568
rect 24084 9528 24090 9540
rect 24590 9537 24602 9540
rect 24636 9537 24648 9571
rect 25148 9568 25176 9608
rect 25400 9605 25412 9639
rect 25446 9636 25458 9639
rect 25498 9636 25504 9648
rect 25446 9608 25504 9636
rect 25446 9605 25458 9608
rect 25400 9599 25458 9605
rect 25498 9596 25504 9608
rect 25556 9596 25562 9648
rect 28077 9639 28135 9645
rect 28077 9636 28089 9639
rect 25608 9608 28089 9636
rect 25608 9568 25636 9608
rect 28077 9605 28089 9608
rect 28123 9605 28135 9639
rect 28077 9599 28135 9605
rect 25148 9540 25636 9568
rect 27801 9571 27859 9577
rect 24590 9531 24648 9537
rect 27801 9537 27813 9571
rect 27847 9568 27859 9571
rect 28258 9568 28264 9580
rect 27847 9540 28264 9568
rect 27847 9537 27859 9540
rect 27801 9531 27859 9537
rect 28258 9528 28264 9540
rect 28316 9528 28322 9580
rect 24857 9503 24915 9509
rect 24857 9469 24869 9503
rect 24903 9500 24915 9503
rect 25133 9503 25191 9509
rect 25133 9500 25145 9503
rect 24903 9472 25145 9500
rect 24903 9469 24915 9472
rect 24857 9463 24915 9469
rect 25133 9469 25145 9472
rect 25179 9469 25191 9503
rect 25133 9463 25191 9469
rect 23474 9432 23480 9444
rect 23435 9404 23480 9432
rect 23474 9392 23480 9404
rect 23532 9392 23538 9444
rect 20119 9336 22508 9364
rect 20119 9333 20131 9336
rect 20073 9327 20131 9333
rect 24670 9324 24676 9376
rect 24728 9364 24734 9376
rect 24872 9364 24900 9463
rect 26510 9432 26516 9444
rect 26471 9404 26516 9432
rect 26510 9392 26516 9404
rect 26568 9392 26574 9444
rect 24728 9336 24900 9364
rect 24728 9324 24734 9336
rect 1104 9274 28888 9296
rect 1104 9222 5582 9274
rect 5634 9222 5646 9274
rect 5698 9222 5710 9274
rect 5762 9222 5774 9274
rect 5826 9222 5838 9274
rect 5890 9222 14846 9274
rect 14898 9222 14910 9274
rect 14962 9222 14974 9274
rect 15026 9222 15038 9274
rect 15090 9222 15102 9274
rect 15154 9222 24110 9274
rect 24162 9222 24174 9274
rect 24226 9222 24238 9274
rect 24290 9222 24302 9274
rect 24354 9222 24366 9274
rect 24418 9222 28888 9274
rect 1104 9200 28888 9222
rect 14550 9160 14556 9172
rect 12636 9132 14556 9160
rect 12636 9104 12664 9132
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 15194 9120 15200 9172
rect 15252 9160 15258 9172
rect 16393 9163 16451 9169
rect 16393 9160 16405 9163
rect 15252 9132 16405 9160
rect 15252 9120 15258 9132
rect 16393 9129 16405 9132
rect 16439 9129 16451 9163
rect 17034 9160 17040 9172
rect 16995 9132 17040 9160
rect 16393 9123 16451 9129
rect 17034 9120 17040 9132
rect 17092 9120 17098 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 18693 9163 18751 9169
rect 18693 9160 18705 9163
rect 17368 9132 18705 9160
rect 17368 9120 17374 9132
rect 18693 9129 18705 9132
rect 18739 9160 18751 9163
rect 23293 9163 23351 9169
rect 18739 9132 22876 9160
rect 18739 9129 18751 9132
rect 18693 9123 18751 9129
rect 10321 9095 10379 9101
rect 10321 9061 10333 9095
rect 10367 9092 10379 9095
rect 12618 9092 12624 9104
rect 10367 9064 12624 9092
rect 10367 9061 10379 9064
rect 10321 9055 10379 9061
rect 8938 9024 8944 9036
rect 8899 8996 8944 9024
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 11072 9033 11100 9064
rect 12618 9052 12624 9064
rect 12676 9052 12682 9104
rect 12894 9052 12900 9104
rect 12952 9092 12958 9104
rect 12952 9064 15056 9092
rect 12952 9052 12958 9064
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 8993 11115 9027
rect 11238 9024 11244 9036
rect 11199 8996 11244 9024
rect 11057 8987 11115 8993
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 13170 9024 13176 9036
rect 13131 8996 13176 9024
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 15028 9033 15056 9064
rect 18598 9052 18604 9104
rect 18656 9092 18662 9104
rect 20806 9092 20812 9104
rect 18656 9064 20812 9092
rect 18656 9052 18662 9064
rect 20806 9052 20812 9064
rect 20864 9052 20870 9104
rect 22370 9052 22376 9104
rect 22428 9092 22434 9104
rect 22649 9095 22707 9101
rect 22649 9092 22661 9095
rect 22428 9064 22661 9092
rect 22428 9052 22434 9064
rect 22649 9061 22661 9064
rect 22695 9061 22707 9095
rect 22649 9055 22707 9061
rect 15013 9027 15071 9033
rect 13872 8996 14320 9024
rect 13872 8984 13878 8996
rect 8386 8956 8392 8968
rect 8347 8928 8392 8956
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 11606 8956 11612 8968
rect 11011 8928 11612 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 11606 8916 11612 8928
rect 11664 8956 11670 8968
rect 11882 8956 11888 8968
rect 11664 8928 11888 8956
rect 11664 8916 11670 8928
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 11974 8916 11980 8968
rect 12032 8956 12038 8968
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 12032 8928 12081 8956
rect 12032 8916 12038 8928
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8956 12955 8959
rect 13446 8956 13452 8968
rect 12943 8928 13452 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 14292 8965 14320 8996
rect 15013 8993 15025 9027
rect 15059 8993 15071 9027
rect 15013 8987 15071 8993
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19702 9024 19708 9036
rect 19392 8996 19708 9024
rect 19392 8984 19398 8996
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 19889 9027 19947 9033
rect 19889 8993 19901 9027
rect 19935 9024 19947 9027
rect 19935 8996 21404 9024
rect 19935 8993 19947 8996
rect 19889 8987 19947 8993
rect 21376 8968 21404 8996
rect 14093 8959 14151 8965
rect 13596 8928 13641 8956
rect 14093 8952 14105 8959
rect 13596 8916 13602 8928
rect 14016 8925 14105 8952
rect 14139 8925 14151 8959
rect 14016 8924 14151 8925
rect 9186 8891 9244 8897
rect 9186 8888 9198 8891
rect 8588 8860 9198 8888
rect 8588 8829 8616 8860
rect 9186 8857 9198 8860
rect 9232 8857 9244 8891
rect 9186 8851 9244 8857
rect 12989 8891 13047 8897
rect 12989 8857 13001 8891
rect 13035 8888 13047 8891
rect 13078 8888 13084 8900
rect 13035 8860 13084 8888
rect 13035 8857 13047 8860
rect 12989 8851 13047 8857
rect 13078 8848 13084 8860
rect 13136 8888 13142 8900
rect 14016 8888 14044 8924
rect 14093 8919 14151 8924
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8925 14335 8959
rect 14458 8956 14464 8968
rect 14419 8928 14464 8956
rect 14277 8919 14335 8925
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 15896 8928 16681 8956
rect 15896 8916 15902 8928
rect 16669 8925 16681 8928
rect 16715 8925 16727 8959
rect 16850 8956 16856 8968
rect 16811 8928 16856 8956
rect 16669 8919 16727 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 17580 8959 17638 8965
rect 17580 8925 17592 8959
rect 17626 8925 17638 8959
rect 17580 8919 17638 8925
rect 13136 8860 14044 8888
rect 13136 8848 13142 8860
rect 14366 8848 14372 8900
rect 14424 8888 14430 8900
rect 15258 8891 15316 8897
rect 15258 8888 15270 8891
rect 14424 8860 14469 8888
rect 14568 8860 15270 8888
rect 14424 8848 14430 8860
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8789 8631 8823
rect 10594 8820 10600 8832
rect 10555 8792 10600 8820
rect 8573 8783 8631 8789
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 11882 8820 11888 8832
rect 11843 8792 11888 8820
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 12526 8820 12532 8832
rect 12487 8792 12532 8820
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 14568 8820 14596 8860
rect 15258 8857 15270 8860
rect 15304 8857 15316 8891
rect 15258 8851 15316 8857
rect 13771 8792 14596 8820
rect 14645 8823 14703 8829
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 14645 8789 14657 8823
rect 14691 8820 14703 8823
rect 14918 8820 14924 8832
rect 14691 8792 14924 8820
rect 14691 8789 14703 8792
rect 14645 8783 14703 8789
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 17328 8820 17356 8919
rect 17494 8848 17500 8900
rect 17552 8888 17558 8900
rect 17604 8888 17632 8919
rect 20346 8916 20352 8968
rect 20404 8956 20410 8968
rect 21269 8959 21327 8965
rect 21269 8956 21281 8959
rect 20404 8928 21281 8956
rect 20404 8916 20410 8928
rect 21269 8925 21281 8928
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 21358 8916 21364 8968
rect 21416 8916 21422 8968
rect 22848 8956 22876 9132
rect 23293 9129 23305 9163
rect 23339 9160 23351 9163
rect 23566 9160 23572 9172
rect 23339 9132 23572 9160
rect 23339 9129 23351 9132
rect 23293 9123 23351 9129
rect 23566 9120 23572 9132
rect 23624 9120 23630 9172
rect 25314 9160 25320 9172
rect 25275 9132 25320 9160
rect 25314 9120 25320 9132
rect 25372 9120 25378 9172
rect 26510 9052 26516 9104
rect 26568 9052 26574 9104
rect 23474 8984 23480 9036
rect 23532 9024 23538 9036
rect 23753 9027 23811 9033
rect 23753 9024 23765 9027
rect 23532 8996 23765 9024
rect 23532 8984 23538 8996
rect 23753 8993 23765 8996
rect 23799 8993 23811 9027
rect 23753 8987 23811 8993
rect 23937 9027 23995 9033
rect 23937 8993 23949 9027
rect 23983 9024 23995 9027
rect 24854 9024 24860 9036
rect 23983 8996 24860 9024
rect 23983 8993 23995 8996
rect 23937 8987 23995 8993
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 25130 8984 25136 9036
rect 25188 9024 25194 9036
rect 25869 9027 25927 9033
rect 25869 9024 25881 9027
rect 25188 8996 25881 9024
rect 25188 8984 25194 8996
rect 25869 8993 25881 8996
rect 25915 8993 25927 9027
rect 26528 9024 26556 9052
rect 26697 9027 26755 9033
rect 26697 9024 26709 9027
rect 26528 8996 26709 9024
rect 25869 8987 25927 8993
rect 26697 8993 26709 8996
rect 26743 8993 26755 9027
rect 26697 8987 26755 8993
rect 23661 8959 23719 8965
rect 23661 8956 23673 8959
rect 22848 8928 23673 8956
rect 23661 8925 23673 8928
rect 23707 8925 23719 8959
rect 23661 8919 23719 8925
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8956 24639 8959
rect 24762 8956 24768 8968
rect 24627 8928 24768 8956
rect 24627 8925 24639 8928
rect 24581 8919 24639 8925
rect 24762 8916 24768 8928
rect 24820 8916 24826 8968
rect 24872 8956 24900 8984
rect 25590 8956 25596 8968
rect 24872 8928 25596 8956
rect 25590 8916 25596 8928
rect 25648 8956 25654 8968
rect 26513 8959 26571 8965
rect 26513 8956 26525 8959
rect 25648 8928 26525 8956
rect 25648 8916 25654 8928
rect 26513 8925 26525 8928
rect 26559 8925 26571 8959
rect 26513 8919 26571 8925
rect 17552 8860 17632 8888
rect 17552 8848 17558 8860
rect 18322 8848 18328 8900
rect 18380 8888 18386 8900
rect 20625 8891 20683 8897
rect 18380 8860 20024 8888
rect 18380 8848 18386 8860
rect 19996 8832 20024 8860
rect 20625 8857 20637 8891
rect 20671 8857 20683 8891
rect 20806 8888 20812 8900
rect 20767 8860 20812 8888
rect 20625 8851 20683 8857
rect 17862 8820 17868 8832
rect 17328 8792 17868 8820
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18138 8780 18144 8832
rect 18196 8820 18202 8832
rect 19245 8823 19303 8829
rect 19245 8820 19257 8823
rect 18196 8792 19257 8820
rect 18196 8780 18202 8792
rect 19245 8789 19257 8792
rect 19291 8789 19303 8823
rect 19978 8820 19984 8832
rect 19939 8792 19984 8820
rect 19245 8783 19303 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 20349 8823 20407 8829
rect 20349 8789 20361 8823
rect 20395 8820 20407 8823
rect 20640 8820 20668 8851
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 21536 8891 21594 8897
rect 21536 8857 21548 8891
rect 21582 8888 21594 8891
rect 21818 8888 21824 8900
rect 21582 8860 21824 8888
rect 21582 8857 21594 8860
rect 21536 8851 21594 8857
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 22094 8848 22100 8900
rect 22152 8888 22158 8900
rect 24397 8891 24455 8897
rect 24397 8888 24409 8891
rect 22152 8860 24409 8888
rect 22152 8848 22158 8860
rect 24397 8857 24409 8860
rect 24443 8888 24455 8891
rect 24670 8888 24676 8900
rect 24443 8860 24676 8888
rect 24443 8857 24455 8860
rect 24397 8851 24455 8857
rect 24670 8848 24676 8860
rect 24728 8848 24734 8900
rect 25685 8891 25743 8897
rect 25685 8857 25697 8891
rect 25731 8888 25743 8891
rect 26329 8891 26387 8897
rect 26329 8888 26341 8891
rect 25731 8860 26341 8888
rect 25731 8857 25743 8860
rect 25685 8851 25743 8857
rect 26329 8857 26341 8860
rect 26375 8857 26387 8891
rect 26329 8851 26387 8857
rect 20990 8820 20996 8832
rect 20395 8792 20668 8820
rect 20951 8792 20996 8820
rect 20395 8789 20407 8792
rect 20349 8783 20407 8789
rect 20990 8780 20996 8792
rect 21048 8780 21054 8832
rect 21082 8780 21088 8832
rect 21140 8820 21146 8832
rect 22370 8820 22376 8832
rect 21140 8792 22376 8820
rect 21140 8780 21146 8792
rect 22370 8780 22376 8792
rect 22428 8780 22434 8832
rect 25774 8820 25780 8832
rect 25735 8792 25780 8820
rect 25774 8780 25780 8792
rect 25832 8780 25838 8832
rect 1104 8730 28888 8752
rect 1104 8678 10214 8730
rect 10266 8678 10278 8730
rect 10330 8678 10342 8730
rect 10394 8678 10406 8730
rect 10458 8678 10470 8730
rect 10522 8678 19478 8730
rect 19530 8678 19542 8730
rect 19594 8678 19606 8730
rect 19658 8678 19670 8730
rect 19722 8678 19734 8730
rect 19786 8678 28888 8730
rect 1104 8656 28888 8678
rect 8386 8576 8392 8628
rect 8444 8616 8450 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 8444 8588 9413 8616
rect 8444 8576 8450 8588
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 9401 8579 9459 8585
rect 12989 8619 13047 8625
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13078 8616 13084 8628
rect 13035 8588 13084 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 13630 8616 13636 8628
rect 13591 8588 13636 8616
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 14182 8576 14188 8628
rect 14240 8616 14246 8628
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 14240 8588 14289 8616
rect 14240 8576 14246 8588
rect 14277 8585 14289 8588
rect 14323 8585 14335 8619
rect 14277 8579 14335 8585
rect 14366 8576 14372 8628
rect 14424 8576 14430 8628
rect 14550 8576 14556 8628
rect 14608 8616 14614 8628
rect 16850 8616 16856 8628
rect 14608 8588 14688 8616
rect 16811 8588 16856 8616
rect 14608 8576 14614 8588
rect 12894 8548 12900 8560
rect 11624 8520 12900 8548
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8480 1455 8483
rect 1486 8480 1492 8492
rect 1443 8452 1492 8480
rect 1443 8449 1455 8452
rect 1397 8443 1455 8449
rect 1486 8440 1492 8452
rect 1544 8440 1550 8492
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 10594 8480 10600 8492
rect 9631 8452 10600 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 10778 8480 10784 8492
rect 10739 8452 10784 8480
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 11514 8480 11520 8492
rect 10919 8452 11520 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 11624 8489 11652 8520
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 14384 8548 14412 8576
rect 14660 8557 14688 8588
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 17310 8616 17316 8628
rect 17271 8588 17316 8616
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 18506 8616 18512 8628
rect 18467 8588 18512 8616
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 19889 8619 19947 8625
rect 19889 8585 19901 8619
rect 19935 8616 19947 8619
rect 21082 8616 21088 8628
rect 19935 8588 21088 8616
rect 19935 8585 19947 8588
rect 19889 8579 19947 8585
rect 21082 8576 21088 8588
rect 21140 8576 21146 8628
rect 21818 8616 21824 8628
rect 21779 8588 21824 8616
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 24026 8616 24032 8628
rect 23987 8588 24032 8616
rect 24026 8576 24032 8588
rect 24084 8576 24090 8628
rect 13740 8520 14412 8548
rect 14645 8551 14703 8557
rect 11882 8489 11888 8492
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8449 11667 8483
rect 11876 8480 11888 8489
rect 11843 8452 11888 8480
rect 11609 8443 11667 8449
rect 11876 8443 11888 8452
rect 11882 8440 11888 8443
rect 11940 8440 11946 8492
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 9858 8412 9864 8424
rect 9815 8384 9864 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 10137 8415 10195 8421
rect 10137 8381 10149 8415
rect 10183 8412 10195 8415
rect 10796 8412 10824 8440
rect 10183 8384 10824 8412
rect 10965 8415 11023 8421
rect 10183 8381 10195 8384
rect 10137 8375 10195 8381
rect 10965 8381 10977 8415
rect 11011 8412 11023 8415
rect 11238 8412 11244 8424
rect 11011 8384 11244 8412
rect 11011 8381 11023 8384
rect 10965 8375 11023 8381
rect 11238 8372 11244 8384
rect 11296 8372 11302 8424
rect 13354 8372 13360 8424
rect 13412 8412 13418 8424
rect 13740 8421 13768 8520
rect 14645 8517 14657 8551
rect 14691 8517 14703 8551
rect 15470 8548 15476 8560
rect 15431 8520 15476 8548
rect 14645 8511 14703 8517
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 18230 8548 18236 8560
rect 15856 8520 18236 8548
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 14415 8483 14473 8489
rect 14415 8480 14427 8483
rect 14332 8452 14427 8480
rect 14332 8440 14338 8452
rect 14415 8449 14427 8452
rect 14461 8449 14473 8483
rect 14550 8480 14556 8492
rect 14511 8452 14556 8480
rect 14415 8443 14473 8449
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 14773 8483 14831 8489
rect 14773 8480 14785 8483
rect 14752 8449 14785 8480
rect 14819 8449 14831 8483
rect 14752 8443 14831 8449
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 13412 8384 13737 8412
rect 13412 8372 13418 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 13909 8415 13967 8421
rect 13909 8381 13921 8415
rect 13955 8412 13967 8415
rect 14752 8412 14780 8443
rect 14918 8440 14924 8492
rect 14976 8480 14982 8492
rect 15289 8483 15347 8489
rect 14976 8452 15021 8480
rect 14976 8440 14982 8452
rect 15289 8449 15301 8483
rect 15335 8480 15347 8483
rect 15856 8480 15884 8520
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 19978 8508 19984 8560
rect 20036 8548 20042 8560
rect 20901 8551 20959 8557
rect 20901 8548 20913 8551
rect 20036 8520 20913 8548
rect 20036 8508 20042 8520
rect 20901 8517 20913 8520
rect 20947 8517 20959 8551
rect 20901 8511 20959 8517
rect 22278 8508 22284 8560
rect 22336 8548 22342 8560
rect 22925 8551 22983 8557
rect 22925 8548 22937 8551
rect 22336 8520 22937 8548
rect 22336 8508 22342 8520
rect 22925 8517 22937 8520
rect 22971 8517 22983 8551
rect 22925 8511 22983 8517
rect 23290 8508 23296 8560
rect 23348 8548 23354 8560
rect 23477 8551 23535 8557
rect 23477 8548 23489 8551
rect 23348 8520 23489 8548
rect 23348 8508 23354 8520
rect 23477 8517 23489 8520
rect 23523 8548 23535 8551
rect 25501 8551 25559 8557
rect 25501 8548 25513 8551
rect 23523 8520 25513 8548
rect 23523 8517 23535 8520
rect 23477 8511 23535 8517
rect 25501 8517 25513 8520
rect 25547 8517 25559 8551
rect 25501 8511 25559 8517
rect 15335 8452 15884 8480
rect 16117 8483 16175 8489
rect 15335 8449 15347 8452
rect 15289 8443 15347 8449
rect 16117 8449 16129 8483
rect 16163 8480 16175 8483
rect 17126 8480 17132 8492
rect 16163 8452 17132 8480
rect 16163 8449 16175 8452
rect 16117 8443 16175 8449
rect 13955 8384 14412 8412
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 1578 8344 1584 8356
rect 1539 8316 1584 8344
rect 1578 8304 1584 8316
rect 1636 8304 1642 8356
rect 13170 8304 13176 8356
rect 13228 8344 13234 8356
rect 13924 8344 13952 8375
rect 13228 8316 13952 8344
rect 13228 8304 13234 8316
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10413 8279 10471 8285
rect 10413 8276 10425 8279
rect 10192 8248 10425 8276
rect 10192 8236 10198 8248
rect 10413 8245 10425 8248
rect 10459 8245 10471 8279
rect 13262 8276 13268 8288
rect 13223 8248 13268 8276
rect 10413 8239 10471 8245
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 14384 8276 14412 8384
rect 14476 8384 14780 8412
rect 14476 8356 14504 8384
rect 14458 8304 14464 8356
rect 14516 8304 14522 8356
rect 15304 8344 15332 8443
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8449 17279 8483
rect 18046 8480 18052 8492
rect 18007 8452 18052 8480
rect 17221 8443 17279 8449
rect 15838 8372 15844 8424
rect 15896 8412 15902 8424
rect 15933 8415 15991 8421
rect 15933 8412 15945 8415
rect 15896 8384 15945 8412
rect 15896 8372 15902 8384
rect 15933 8381 15945 8384
rect 15979 8412 15991 8415
rect 16022 8412 16028 8424
rect 15979 8384 16028 8412
rect 15979 8381 15991 8384
rect 15933 8375 15991 8381
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 16666 8372 16672 8424
rect 16724 8412 16730 8424
rect 17236 8412 17264 8443
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 19058 8480 19064 8492
rect 18371 8452 19064 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 19153 8483 19211 8489
rect 19153 8449 19165 8483
rect 19199 8480 19211 8483
rect 19334 8480 19340 8492
rect 19199 8452 19340 8480
rect 19199 8449 19211 8452
rect 19153 8443 19211 8449
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 19794 8480 19800 8492
rect 19755 8452 19800 8480
rect 19794 8440 19800 8452
rect 19852 8440 19858 8492
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8480 20683 8483
rect 20990 8480 20996 8492
rect 20671 8452 20996 8480
rect 20671 8449 20683 8452
rect 20625 8443 20683 8449
rect 20990 8440 20996 8452
rect 21048 8440 21054 8492
rect 22005 8483 22063 8489
rect 22005 8449 22017 8483
rect 22051 8480 22063 8483
rect 22186 8480 22192 8492
rect 22051 8452 22192 8480
rect 22051 8449 22063 8452
rect 22005 8443 22063 8449
rect 22186 8440 22192 8452
rect 22244 8440 22250 8492
rect 23842 8480 23848 8492
rect 23803 8452 23848 8480
rect 23842 8440 23848 8452
rect 23900 8440 23906 8492
rect 24673 8483 24731 8489
rect 24673 8449 24685 8483
rect 24719 8480 24731 8483
rect 24946 8480 24952 8492
rect 24719 8452 24952 8480
rect 24719 8449 24731 8452
rect 24673 8443 24731 8449
rect 24946 8440 24952 8452
rect 25004 8440 25010 8492
rect 27893 8483 27951 8489
rect 27893 8449 27905 8483
rect 27939 8480 27951 8483
rect 28350 8480 28356 8492
rect 27939 8452 28356 8480
rect 27939 8449 27951 8452
rect 27893 8443 27951 8449
rect 28350 8440 28356 8452
rect 28408 8440 28414 8492
rect 16724 8384 17264 8412
rect 17497 8415 17555 8421
rect 16724 8372 16730 8384
rect 17497 8381 17509 8415
rect 17543 8381 17555 8415
rect 18138 8412 18144 8424
rect 18099 8384 18144 8412
rect 17497 8375 17555 8381
rect 14568 8316 15332 8344
rect 16301 8347 16359 8353
rect 14568 8276 14596 8316
rect 16301 8313 16313 8347
rect 16347 8344 16359 8347
rect 16758 8344 16764 8356
rect 16347 8316 16764 8344
rect 16347 8313 16359 8316
rect 16301 8307 16359 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 17512 8344 17540 8375
rect 18138 8372 18144 8384
rect 18196 8372 18202 8424
rect 20073 8415 20131 8421
rect 20073 8381 20085 8415
rect 20119 8412 20131 8415
rect 22738 8412 22744 8424
rect 20119 8384 22744 8412
rect 20119 8381 20131 8384
rect 20073 8375 20131 8381
rect 22738 8372 22744 8384
rect 22796 8412 22802 8424
rect 23293 8415 23351 8421
rect 23293 8412 23305 8415
rect 22796 8384 23305 8412
rect 22796 8372 22802 8384
rect 23293 8381 23305 8384
rect 23339 8381 23351 8415
rect 23293 8375 23351 8381
rect 24397 8415 24455 8421
rect 24397 8381 24409 8415
rect 24443 8381 24455 8415
rect 24578 8412 24584 8424
rect 24539 8384 24584 8412
rect 24397 8375 24455 8381
rect 18414 8344 18420 8356
rect 17512 8316 18420 8344
rect 18414 8304 18420 8316
rect 18472 8344 18478 8356
rect 18969 8347 19027 8353
rect 18969 8344 18981 8347
rect 18472 8316 18981 8344
rect 18472 8304 18478 8316
rect 18969 8313 18981 8316
rect 19015 8313 19027 8347
rect 24412 8344 24440 8375
rect 24578 8372 24584 8384
rect 24636 8372 24642 8424
rect 25130 8412 25136 8424
rect 24872 8384 25136 8412
rect 24872 8344 24900 8384
rect 25130 8372 25136 8384
rect 25188 8412 25194 8424
rect 25317 8415 25375 8421
rect 25317 8412 25329 8415
rect 25188 8384 25329 8412
rect 25188 8372 25194 8384
rect 25317 8381 25329 8384
rect 25363 8381 25375 8415
rect 25317 8375 25375 8381
rect 24412 8316 24900 8344
rect 25041 8347 25099 8353
rect 18969 8307 19027 8313
rect 25041 8313 25053 8347
rect 25087 8344 25099 8347
rect 26510 8344 26516 8356
rect 25087 8316 26516 8344
rect 25087 8313 25099 8316
rect 25041 8307 25099 8313
rect 26510 8304 26516 8316
rect 26568 8304 26574 8356
rect 18322 8276 18328 8288
rect 14384 8248 14596 8276
rect 18283 8248 18328 8276
rect 18322 8236 18328 8248
rect 18380 8236 18386 8288
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 19429 8279 19487 8285
rect 19429 8276 19441 8279
rect 19392 8248 19441 8276
rect 19392 8236 19398 8248
rect 19429 8245 19441 8248
rect 19475 8245 19487 8279
rect 20438 8276 20444 8288
rect 20399 8248 20444 8276
rect 19429 8239 19487 8245
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 22830 8276 22836 8288
rect 22791 8248 22836 8276
rect 22830 8236 22836 8248
rect 22888 8236 22894 8288
rect 28166 8276 28172 8288
rect 28127 8248 28172 8276
rect 28166 8236 28172 8248
rect 28224 8236 28230 8288
rect 1104 8186 28888 8208
rect 1104 8134 5582 8186
rect 5634 8134 5646 8186
rect 5698 8134 5710 8186
rect 5762 8134 5774 8186
rect 5826 8134 5838 8186
rect 5890 8134 14846 8186
rect 14898 8134 14910 8186
rect 14962 8134 14974 8186
rect 15026 8134 15038 8186
rect 15090 8134 15102 8186
rect 15154 8134 24110 8186
rect 24162 8134 24174 8186
rect 24226 8134 24238 8186
rect 24290 8134 24302 8186
rect 24354 8134 24366 8186
rect 24418 8134 28888 8186
rect 1104 8112 28888 8134
rect 12894 8072 12900 8084
rect 10152 8044 12900 8072
rect 10152 7945 10180 8044
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13446 8072 13452 8084
rect 13407 8044 13452 8072
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13872 8044 14105 8072
rect 13872 8032 13878 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 14608 8044 15117 8072
rect 14608 8032 14614 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 19794 8032 19800 8084
rect 19852 8072 19858 8084
rect 20073 8075 20131 8081
rect 20073 8072 20085 8075
rect 19852 8044 20085 8072
rect 19852 8032 19858 8044
rect 20073 8041 20085 8044
rect 20119 8041 20131 8075
rect 28166 8072 28172 8084
rect 20073 8035 20131 8041
rect 20180 8044 28172 8072
rect 11514 8004 11520 8016
rect 11475 7976 11520 8004
rect 11514 7964 11520 7976
rect 11572 7964 11578 8016
rect 11974 8004 11980 8016
rect 11935 7976 11980 8004
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 18322 7964 18328 8016
rect 18380 8004 18386 8016
rect 20180 8004 20208 8044
rect 28166 8032 28172 8044
rect 28224 8032 28230 8084
rect 18380 7976 20208 8004
rect 18380 7964 18386 7976
rect 21358 7964 21364 8016
rect 21416 8004 21422 8016
rect 21729 8007 21787 8013
rect 21729 8004 21741 8007
rect 21416 7976 21741 8004
rect 21416 7964 21422 7976
rect 21729 7973 21741 7976
rect 21775 7973 21787 8007
rect 24026 8004 24032 8016
rect 23939 7976 24032 8004
rect 21729 7967 21787 7973
rect 24026 7964 24032 7976
rect 24084 8004 24090 8016
rect 24578 8004 24584 8016
rect 24084 7976 24584 8004
rect 24084 7964 24090 7976
rect 24578 7964 24584 7976
rect 24636 7964 24642 8016
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7905 10195 7939
rect 12526 7936 12532 7948
rect 10137 7899 10195 7905
rect 12176 7908 12532 7936
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 10042 7868 10048 7880
rect 9723 7840 10048 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 12176 7877 12204 7908
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 12820 7908 14473 7936
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 12250 7828 12256 7880
rect 12308 7868 12314 7880
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 12308 7840 12357 7868
rect 12308 7828 12314 7840
rect 12345 7837 12357 7840
rect 12391 7868 12403 7871
rect 12820 7868 12848 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 19521 7939 19579 7945
rect 19521 7905 19533 7939
rect 19567 7936 19579 7939
rect 19978 7936 19984 7948
rect 19567 7908 19984 7936
rect 19567 7905 19579 7908
rect 19521 7899 19579 7905
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 20346 7936 20352 7948
rect 20307 7908 20352 7936
rect 20346 7896 20352 7908
rect 20404 7896 20410 7948
rect 22094 7896 22100 7948
rect 22152 7936 22158 7948
rect 22649 7939 22707 7945
rect 22649 7936 22661 7939
rect 22152 7908 22661 7936
rect 22152 7896 22158 7908
rect 22649 7905 22661 7908
rect 22695 7905 22707 7939
rect 22649 7899 22707 7905
rect 12986 7868 12992 7880
rect 12391 7840 12848 7868
rect 12947 7840 12992 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7868 14703 7871
rect 15102 7868 15108 7880
rect 14691 7840 15108 7868
rect 14691 7837 14703 7840
rect 14645 7831 14703 7837
rect 15102 7828 15108 7840
rect 15160 7828 15166 7880
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7868 16543 7871
rect 16945 7871 17003 7877
rect 16945 7868 16957 7871
rect 16531 7840 16957 7868
rect 16531 7837 16543 7840
rect 16485 7831 16543 7837
rect 16945 7837 16957 7840
rect 16991 7868 17003 7871
rect 17770 7868 17776 7880
rect 16991 7840 17776 7868
rect 16991 7837 17003 7840
rect 16945 7831 17003 7837
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19334 7868 19340 7880
rect 18923 7840 19340 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 20438 7828 20444 7880
rect 20496 7868 20502 7880
rect 20605 7871 20663 7877
rect 20605 7868 20617 7871
rect 20496 7840 20617 7868
rect 20496 7828 20502 7840
rect 20605 7837 20617 7840
rect 20651 7837 20663 7871
rect 20605 7831 20663 7837
rect 24670 7828 24676 7880
rect 24728 7868 24734 7880
rect 26053 7871 26111 7877
rect 26053 7868 26065 7871
rect 24728 7840 26065 7868
rect 24728 7828 24734 7840
rect 26053 7837 26065 7840
rect 26099 7837 26111 7871
rect 26510 7868 26516 7880
rect 26471 7840 26516 7868
rect 26053 7831 26111 7837
rect 26510 7828 26516 7840
rect 26568 7828 26574 7880
rect 10382 7803 10440 7809
rect 10382 7800 10394 7803
rect 9876 7772 10394 7800
rect 9876 7741 9904 7772
rect 10382 7769 10394 7772
rect 10428 7769 10440 7803
rect 10382 7763 10440 7769
rect 11514 7760 11520 7812
rect 11572 7800 11578 7812
rect 14274 7800 14280 7812
rect 11572 7772 14280 7800
rect 11572 7760 11578 7772
rect 14274 7760 14280 7772
rect 14332 7760 14338 7812
rect 16206 7800 16212 7812
rect 16264 7809 16270 7812
rect 16176 7772 16212 7800
rect 16206 7760 16212 7772
rect 16264 7763 16276 7809
rect 16264 7760 16270 7763
rect 17034 7760 17040 7812
rect 17092 7800 17098 7812
rect 17190 7803 17248 7809
rect 17190 7800 17202 7803
rect 17092 7772 17202 7800
rect 17092 7760 17098 7772
rect 17190 7769 17202 7772
rect 17236 7769 17248 7803
rect 19613 7803 19671 7809
rect 17190 7763 17248 7769
rect 18340 7772 18920 7800
rect 9861 7735 9919 7741
rect 9861 7701 9873 7735
rect 9907 7701 9919 7735
rect 14826 7732 14832 7744
rect 14787 7704 14832 7732
rect 9861 7695 9919 7701
rect 14826 7692 14832 7704
rect 14884 7692 14890 7744
rect 17678 7692 17684 7744
rect 17736 7732 17742 7744
rect 18340 7741 18368 7772
rect 18325 7735 18383 7741
rect 18325 7732 18337 7735
rect 17736 7704 18337 7732
rect 17736 7692 17742 7704
rect 18325 7701 18337 7704
rect 18371 7701 18383 7735
rect 18325 7695 18383 7701
rect 18693 7735 18751 7741
rect 18693 7701 18705 7735
rect 18739 7732 18751 7735
rect 18782 7732 18788 7744
rect 18739 7704 18788 7732
rect 18739 7701 18751 7704
rect 18693 7695 18751 7701
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 18892 7732 18920 7772
rect 19613 7769 19625 7803
rect 19659 7800 19671 7803
rect 19886 7800 19892 7812
rect 19659 7772 19892 7800
rect 19659 7769 19671 7772
rect 19613 7763 19671 7769
rect 19886 7760 19892 7772
rect 19944 7760 19950 7812
rect 22094 7760 22100 7812
rect 22152 7800 22158 7812
rect 22894 7803 22952 7809
rect 22894 7800 22906 7803
rect 22152 7772 22906 7800
rect 22152 7760 22158 7772
rect 22894 7769 22906 7772
rect 22940 7769 22952 7803
rect 22894 7763 22952 7769
rect 25808 7803 25866 7809
rect 25808 7769 25820 7803
rect 25854 7800 25866 7803
rect 25854 7772 26372 7800
rect 25854 7769 25866 7772
rect 25808 7763 25866 7769
rect 19705 7735 19763 7741
rect 19705 7732 19717 7735
rect 18892 7704 19717 7732
rect 19705 7701 19717 7704
rect 19751 7701 19763 7735
rect 19705 7695 19763 7701
rect 24673 7735 24731 7741
rect 24673 7701 24685 7735
rect 24719 7732 24731 7735
rect 25406 7732 25412 7744
rect 24719 7704 25412 7732
rect 24719 7701 24731 7704
rect 24673 7695 24731 7701
rect 25406 7692 25412 7704
rect 25464 7692 25470 7744
rect 26344 7741 26372 7772
rect 26329 7735 26387 7741
rect 26329 7701 26341 7735
rect 26375 7701 26387 7735
rect 26329 7695 26387 7701
rect 1104 7642 28888 7664
rect 1104 7590 10214 7642
rect 10266 7590 10278 7642
rect 10330 7590 10342 7642
rect 10394 7590 10406 7642
rect 10458 7590 10470 7642
rect 10522 7590 19478 7642
rect 19530 7590 19542 7642
rect 19594 7590 19606 7642
rect 19658 7590 19670 7642
rect 19722 7590 19734 7642
rect 19786 7590 28888 7642
rect 1104 7568 28888 7590
rect 10042 7528 10048 7540
rect 10003 7500 10048 7528
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 11606 7488 11612 7540
rect 11664 7528 11670 7540
rect 15102 7528 15108 7540
rect 11664 7500 14228 7528
rect 15063 7500 15108 7528
rect 11664 7488 11670 7500
rect 9858 7420 9864 7472
rect 9916 7460 9922 7472
rect 9916 7432 10364 7460
rect 9916 7420 9922 7432
rect 10134 7352 10140 7404
rect 10192 7392 10198 7404
rect 10336 7401 10364 7432
rect 14200 7404 14228 7500
rect 15102 7488 15108 7500
rect 15160 7488 15166 7540
rect 16206 7488 16212 7540
rect 16264 7528 16270 7540
rect 16301 7531 16359 7537
rect 16301 7528 16313 7531
rect 16264 7500 16313 7528
rect 16264 7488 16270 7500
rect 16301 7497 16313 7500
rect 16347 7497 16359 7531
rect 16301 7491 16359 7497
rect 16945 7531 17003 7537
rect 16945 7497 16957 7531
rect 16991 7528 17003 7531
rect 17034 7528 17040 7540
rect 16991 7500 17040 7528
rect 16991 7497 17003 7500
rect 16945 7491 17003 7497
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 17126 7488 17132 7540
rect 17184 7528 17190 7540
rect 17221 7531 17279 7537
rect 17221 7528 17233 7531
rect 17184 7500 17233 7528
rect 17184 7488 17190 7500
rect 17221 7497 17233 7500
rect 17267 7497 17279 7531
rect 17678 7528 17684 7540
rect 17639 7500 17684 7528
rect 17221 7491 17279 7497
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 22094 7488 22100 7540
rect 22152 7528 22158 7540
rect 22833 7531 22891 7537
rect 22152 7500 22197 7528
rect 22152 7488 22158 7500
rect 22833 7497 22845 7531
rect 22879 7528 22891 7531
rect 24026 7528 24032 7540
rect 22879 7500 24032 7528
rect 22879 7497 22891 7500
rect 22833 7491 22891 7497
rect 24026 7488 24032 7500
rect 24084 7488 24090 7540
rect 24946 7528 24952 7540
rect 24907 7500 24952 7528
rect 24946 7488 24952 7500
rect 25004 7488 25010 7540
rect 25406 7528 25412 7540
rect 25319 7500 25412 7528
rect 25406 7488 25412 7500
rect 25464 7528 25470 7540
rect 25774 7528 25780 7540
rect 25464 7500 25780 7528
rect 25464 7488 25470 7500
rect 25774 7488 25780 7500
rect 25832 7488 25838 7540
rect 14826 7420 14832 7472
rect 14884 7460 14890 7472
rect 14884 7432 16160 7460
rect 14884 7420 14890 7432
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 10192 7364 10241 7392
rect 10192 7352 10198 7364
rect 10229 7361 10241 7364
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 12250 7392 12256 7404
rect 12211 7364 12256 7392
rect 10321 7355 10379 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12345 7395 12403 7401
rect 12345 7361 12357 7395
rect 12391 7392 12403 7395
rect 13262 7392 13268 7404
rect 12391 7364 13268 7392
rect 12391 7361 12403 7364
rect 12345 7355 12403 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 13357 7395 13415 7401
rect 13357 7361 13369 7395
rect 13403 7392 13415 7395
rect 14182 7392 14188 7404
rect 13403 7364 13860 7392
rect 14143 7364 14188 7392
rect 13403 7361 13415 7364
rect 13357 7355 13415 7361
rect 12268 7324 12296 7352
rect 13173 7327 13231 7333
rect 13173 7324 13185 7327
rect 12268 7296 13185 7324
rect 13173 7293 13185 7296
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 13832 7265 13860 7364
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7392 14335 7395
rect 14458 7392 14464 7404
rect 14323 7364 14464 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 15378 7352 15384 7404
rect 15436 7392 15442 7404
rect 16132 7401 16160 7432
rect 17862 7420 17868 7472
rect 17920 7460 17926 7472
rect 20346 7460 20352 7472
rect 17920 7432 20352 7460
rect 17920 7420 17926 7432
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15436 7364 15485 7392
rect 15436 7352 15442 7364
rect 15473 7361 15485 7364
rect 15519 7392 15531 7395
rect 16117 7395 16175 7401
rect 15519 7364 16068 7392
rect 15519 7361 15531 7364
rect 15473 7355 15531 7361
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7293 14427 7327
rect 14369 7287 14427 7293
rect 13817 7259 13875 7265
rect 13817 7225 13829 7259
rect 13863 7225 13875 7259
rect 14384 7256 14412 7287
rect 14550 7284 14556 7336
rect 14608 7324 14614 7336
rect 15565 7327 15623 7333
rect 15565 7324 15577 7327
rect 14608 7296 15577 7324
rect 14608 7284 14614 7296
rect 15565 7293 15577 7296
rect 15611 7293 15623 7327
rect 15565 7287 15623 7293
rect 15657 7327 15715 7333
rect 15657 7293 15669 7327
rect 15703 7293 15715 7327
rect 16040 7324 16068 7364
rect 16117 7361 16129 7395
rect 16163 7361 16175 7395
rect 16758 7392 16764 7404
rect 16719 7364 16764 7392
rect 16117 7355 16175 7361
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 17586 7392 17592 7404
rect 17547 7364 17592 7392
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 18524 7401 18552 7432
rect 20346 7420 20352 7432
rect 20404 7420 20410 7472
rect 21358 7420 21364 7472
rect 21416 7460 21422 7472
rect 22741 7463 22799 7469
rect 22741 7460 22753 7463
rect 21416 7432 22753 7460
rect 21416 7420 21422 7432
rect 22741 7429 22753 7432
rect 22787 7429 22799 7463
rect 22741 7423 22799 7429
rect 18782 7401 18788 7404
rect 18509 7395 18567 7401
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 18776 7392 18788 7401
rect 18743 7364 18788 7392
rect 18509 7355 18567 7361
rect 18776 7355 18788 7364
rect 18782 7352 18788 7355
rect 18840 7352 18846 7404
rect 21913 7395 21971 7401
rect 21913 7361 21925 7395
rect 21959 7392 21971 7395
rect 22186 7392 22192 7404
rect 21959 7364 22192 7392
rect 21959 7361 21971 7364
rect 21913 7355 21971 7361
rect 22186 7352 22192 7364
rect 22244 7352 22250 7404
rect 24854 7352 24860 7404
rect 24912 7392 24918 7404
rect 25317 7395 25375 7401
rect 25317 7392 25329 7395
rect 24912 7364 25329 7392
rect 24912 7352 24918 7364
rect 25317 7361 25329 7364
rect 25363 7361 25375 7395
rect 25317 7355 25375 7361
rect 27801 7395 27859 7401
rect 27801 7361 27813 7395
rect 27847 7392 27859 7395
rect 28350 7392 28356 7404
rect 27847 7364 28356 7392
rect 27847 7361 27859 7364
rect 27801 7355 27859 7361
rect 28350 7352 28356 7364
rect 28408 7352 28414 7404
rect 17604 7324 17632 7352
rect 16040 7296 17632 7324
rect 17865 7327 17923 7333
rect 15657 7287 15715 7293
rect 17865 7293 17877 7327
rect 17911 7324 17923 7327
rect 18322 7324 18328 7336
rect 17911 7296 18328 7324
rect 17911 7293 17923 7296
rect 17865 7287 17923 7293
rect 15470 7256 15476 7268
rect 14384 7228 15476 7256
rect 13817 7219 13875 7225
rect 15470 7216 15476 7228
rect 15528 7256 15534 7268
rect 15672 7256 15700 7287
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 22830 7284 22836 7336
rect 22888 7324 22894 7336
rect 22925 7327 22983 7333
rect 22925 7324 22937 7327
rect 22888 7296 22937 7324
rect 22888 7284 22894 7296
rect 22925 7293 22937 7296
rect 22971 7293 22983 7327
rect 25590 7324 25596 7336
rect 25551 7296 25596 7324
rect 22925 7287 22983 7293
rect 25590 7284 25596 7296
rect 25648 7284 25654 7336
rect 15528 7228 15700 7256
rect 15528 7216 15534 7228
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12529 7191 12587 7197
rect 12529 7188 12541 7191
rect 12492 7160 12541 7188
rect 12492 7148 12498 7160
rect 12529 7157 12541 7160
rect 12575 7157 12587 7191
rect 13538 7188 13544 7200
rect 13499 7160 13544 7188
rect 12529 7151 12587 7157
rect 13538 7148 13544 7160
rect 13596 7148 13602 7200
rect 19886 7188 19892 7200
rect 19847 7160 19892 7188
rect 19886 7148 19892 7160
rect 19944 7148 19950 7200
rect 22370 7188 22376 7200
rect 22331 7160 22376 7188
rect 22370 7148 22376 7160
rect 22428 7148 22434 7200
rect 28166 7188 28172 7200
rect 28127 7160 28172 7188
rect 28166 7148 28172 7160
rect 28224 7148 28230 7200
rect 1104 7098 28888 7120
rect 1104 7046 5582 7098
rect 5634 7046 5646 7098
rect 5698 7046 5710 7098
rect 5762 7046 5774 7098
rect 5826 7046 5838 7098
rect 5890 7046 14846 7098
rect 14898 7046 14910 7098
rect 14962 7046 14974 7098
rect 15026 7046 15038 7098
rect 15090 7046 15102 7098
rect 15154 7046 24110 7098
rect 24162 7046 24174 7098
rect 24226 7046 24238 7098
rect 24290 7046 24302 7098
rect 24354 7046 24366 7098
rect 24418 7046 28888 7098
rect 1104 7024 28888 7046
rect 22186 6984 22192 6996
rect 22147 6956 22192 6984
rect 22186 6944 22192 6956
rect 22244 6944 22250 6996
rect 18322 6916 18328 6928
rect 16960 6888 18328 6916
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 13722 6848 13728 6860
rect 12952 6820 13728 6848
rect 12952 6808 12958 6820
rect 13722 6808 13728 6820
rect 13780 6848 13786 6860
rect 16960 6857 16988 6888
rect 18322 6876 18328 6888
rect 18380 6876 18386 6928
rect 22830 6916 22836 6928
rect 22066 6888 22836 6916
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13780 6820 14105 6848
rect 13780 6808 13786 6820
rect 14093 6817 14105 6820
rect 14139 6817 14151 6851
rect 14093 6811 14151 6817
rect 16945 6851 17003 6857
rect 16945 6817 16957 6851
rect 16991 6817 17003 6851
rect 16945 6811 17003 6817
rect 17586 6808 17592 6860
rect 17644 6848 17650 6860
rect 18417 6851 18475 6857
rect 18417 6848 18429 6851
rect 17644 6820 18429 6848
rect 17644 6808 17650 6820
rect 18417 6817 18429 6820
rect 18463 6848 18475 6851
rect 19150 6848 19156 6860
rect 18463 6820 19156 6848
rect 18463 6817 18475 6820
rect 18417 6811 18475 6817
rect 19150 6808 19156 6820
rect 19208 6808 19214 6860
rect 19978 6808 19984 6860
rect 20036 6848 20042 6860
rect 21545 6851 21603 6857
rect 21545 6848 21557 6851
rect 20036 6820 21557 6848
rect 20036 6808 20042 6820
rect 21545 6817 21557 6820
rect 21591 6848 21603 6851
rect 22066 6848 22094 6888
rect 22830 6876 22836 6888
rect 22888 6876 22894 6928
rect 22738 6848 22744 6860
rect 21591 6820 22094 6848
rect 22699 6820 22744 6848
rect 21591 6817 21603 6820
rect 21545 6811 21603 6817
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 24854 6848 24860 6860
rect 24815 6820 24860 6848
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 24949 6851 25007 6857
rect 24949 6817 24961 6851
rect 24995 6817 25007 6851
rect 24949 6811 25007 6817
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 12912 6780 12940 6808
rect 13538 6780 13544 6792
rect 11931 6752 12940 6780
rect 13499 6752 13544 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 17678 6740 17684 6792
rect 17736 6780 17742 6792
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 17736 6752 17877 6780
rect 17736 6740 17742 6752
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 12152 6715 12210 6721
rect 12152 6681 12164 6715
rect 12198 6712 12210 6715
rect 12250 6712 12256 6724
rect 12198 6684 12256 6712
rect 12198 6681 12210 6684
rect 12152 6675 12210 6681
rect 12250 6672 12256 6684
rect 12308 6672 12314 6724
rect 14338 6715 14396 6721
rect 14338 6712 14350 6715
rect 13740 6684 14350 6712
rect 13265 6647 13323 6653
rect 13265 6613 13277 6647
rect 13311 6644 13323 6647
rect 13354 6644 13360 6656
rect 13311 6616 13360 6644
rect 13311 6613 13323 6616
rect 13265 6607 13323 6613
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13740 6653 13768 6684
rect 14338 6681 14350 6684
rect 14384 6681 14396 6715
rect 16669 6715 16727 6721
rect 16669 6712 16681 6715
rect 14338 6675 14396 6681
rect 15948 6684 16681 6712
rect 13725 6647 13783 6653
rect 13725 6613 13737 6647
rect 13771 6613 13783 6647
rect 13725 6607 13783 6613
rect 14458 6604 14464 6656
rect 14516 6644 14522 6656
rect 15473 6647 15531 6653
rect 15473 6644 15485 6647
rect 14516 6616 15485 6644
rect 14516 6604 14522 6616
rect 15473 6613 15485 6616
rect 15519 6613 15531 6647
rect 15473 6607 15531 6613
rect 15838 6604 15844 6656
rect 15896 6644 15902 6656
rect 15948 6653 15976 6684
rect 16669 6681 16681 6684
rect 16715 6681 16727 6715
rect 18064 6712 18092 6743
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19392 6752 19441 6780
rect 19392 6740 19398 6752
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 21266 6740 21272 6792
rect 21324 6780 21330 6792
rect 21361 6783 21419 6789
rect 21361 6780 21373 6783
rect 21324 6752 21373 6780
rect 21324 6740 21330 6752
rect 21361 6749 21373 6752
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 22370 6740 22376 6792
rect 22428 6780 22434 6792
rect 22557 6783 22615 6789
rect 22557 6780 22569 6783
rect 22428 6752 22569 6780
rect 22428 6740 22434 6752
rect 22557 6749 22569 6752
rect 22603 6749 22615 6783
rect 22557 6743 22615 6749
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6780 23627 6783
rect 23658 6780 23664 6792
rect 23615 6752 23664 6780
rect 23615 6749 23627 6752
rect 23569 6743 23627 6749
rect 23584 6712 23612 6743
rect 23658 6740 23664 6752
rect 23716 6740 23722 6792
rect 23753 6783 23811 6789
rect 23753 6749 23765 6783
rect 23799 6780 23811 6783
rect 23799 6752 24440 6780
rect 23799 6749 23811 6752
rect 23753 6743 23811 6749
rect 18064 6684 23612 6712
rect 16669 6675 16727 6681
rect 15933 6647 15991 6653
rect 15933 6644 15945 6647
rect 15896 6616 15945 6644
rect 15896 6604 15902 6616
rect 15933 6613 15945 6616
rect 15979 6613 15991 6647
rect 15933 6607 15991 6613
rect 16114 6604 16120 6656
rect 16172 6644 16178 6656
rect 16301 6647 16359 6653
rect 16301 6644 16313 6647
rect 16172 6616 16313 6644
rect 16172 6604 16178 6616
rect 16301 6613 16313 6616
rect 16347 6613 16359 6647
rect 16301 6607 16359 6613
rect 16761 6647 16819 6653
rect 16761 6613 16773 6647
rect 16807 6644 16819 6647
rect 16850 6644 16856 6656
rect 16807 6616 16856 6644
rect 16807 6613 16819 6616
rect 16761 6607 16819 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 17034 6604 17040 6656
rect 17092 6644 17098 6656
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17092 6616 17693 6644
rect 17092 6604 17098 6616
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 19242 6644 19248 6656
rect 19203 6616 19248 6644
rect 17681 6607 17739 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 20806 6604 20812 6656
rect 20864 6644 20870 6656
rect 20993 6647 21051 6653
rect 20993 6644 21005 6647
rect 20864 6616 21005 6644
rect 20864 6604 20870 6616
rect 20993 6613 21005 6616
rect 21039 6613 21051 6647
rect 20993 6607 21051 6613
rect 21453 6647 21511 6653
rect 21453 6613 21465 6647
rect 21499 6644 21511 6647
rect 22094 6644 22100 6656
rect 21499 6616 22100 6644
rect 21499 6613 21511 6616
rect 21453 6607 21511 6613
rect 22094 6604 22100 6616
rect 22152 6604 22158 6656
rect 22646 6644 22652 6656
rect 22607 6616 22652 6644
rect 22646 6604 22652 6616
rect 22704 6604 22710 6656
rect 23658 6604 23664 6656
rect 23716 6644 23722 6656
rect 24412 6653 24440 6752
rect 24486 6740 24492 6792
rect 24544 6780 24550 6792
rect 24964 6780 24992 6811
rect 24544 6752 24992 6780
rect 24544 6740 24550 6752
rect 24578 6672 24584 6724
rect 24636 6712 24642 6724
rect 24765 6715 24823 6721
rect 24765 6712 24777 6715
rect 24636 6684 24777 6712
rect 24636 6672 24642 6684
rect 24765 6681 24777 6684
rect 24811 6712 24823 6715
rect 25409 6715 25467 6721
rect 25409 6712 25421 6715
rect 24811 6684 25421 6712
rect 24811 6681 24823 6684
rect 24765 6675 24823 6681
rect 25409 6681 25421 6684
rect 25455 6712 25467 6715
rect 28166 6712 28172 6724
rect 25455 6684 28172 6712
rect 25455 6681 25467 6684
rect 25409 6675 25467 6681
rect 28166 6672 28172 6684
rect 28224 6672 28230 6724
rect 23937 6647 23995 6653
rect 23937 6644 23949 6647
rect 23716 6616 23949 6644
rect 23716 6604 23722 6616
rect 23937 6613 23949 6616
rect 23983 6613 23995 6647
rect 23937 6607 23995 6613
rect 24397 6647 24455 6653
rect 24397 6613 24409 6647
rect 24443 6613 24455 6647
rect 24397 6607 24455 6613
rect 1104 6554 28888 6576
rect 1104 6502 10214 6554
rect 10266 6502 10278 6554
rect 10330 6502 10342 6554
rect 10394 6502 10406 6554
rect 10458 6502 10470 6554
rect 10522 6502 19478 6554
rect 19530 6502 19542 6554
rect 19594 6502 19606 6554
rect 19658 6502 19670 6554
rect 19722 6502 19734 6554
rect 19786 6502 28888 6554
rect 1104 6480 28888 6502
rect 12250 6440 12256 6452
rect 12211 6412 12256 6440
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 16761 6443 16819 6449
rect 16761 6409 16773 6443
rect 16807 6440 16819 6443
rect 17586 6440 17592 6452
rect 16807 6412 17592 6440
rect 16807 6409 16819 6412
rect 16761 6403 16819 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 20806 6440 20812 6452
rect 20767 6412 20812 6440
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 24486 6440 24492 6452
rect 22066 6412 24492 6440
rect 16022 6332 16028 6384
rect 16080 6372 16086 6384
rect 17862 6372 17868 6384
rect 16080 6344 16252 6372
rect 16080 6332 16086 6344
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 15473 6307 15531 6313
rect 12492 6276 12537 6304
rect 12492 6264 12498 6276
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 15933 6307 15991 6313
rect 15933 6304 15945 6307
rect 15519 6276 15945 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 15933 6273 15945 6276
rect 15979 6273 15991 6307
rect 16114 6304 16120 6316
rect 16075 6276 16120 6304
rect 15933 6267 15991 6273
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 16224 6313 16252 6344
rect 17512 6344 17868 6372
rect 17512 6316 17540 6344
rect 17862 6332 17868 6344
rect 17920 6332 17926 6384
rect 18322 6332 18328 6384
rect 18380 6372 18386 6384
rect 22066 6372 22094 6412
rect 24486 6400 24492 6412
rect 24544 6400 24550 6452
rect 24854 6400 24860 6452
rect 24912 6440 24918 6452
rect 25501 6443 25559 6449
rect 25501 6440 25513 6443
rect 24912 6412 25513 6440
rect 24912 6400 24918 6412
rect 25501 6409 25513 6412
rect 25547 6409 25559 6443
rect 25501 6403 25559 6409
rect 24670 6372 24676 6384
rect 18380 6344 22094 6372
rect 24136 6344 24676 6372
rect 18380 6332 18386 6344
rect 16209 6307 16267 6313
rect 16209 6273 16221 6307
rect 16255 6273 16267 6307
rect 17034 6304 17040 6316
rect 16995 6276 17040 6304
rect 16209 6267 16267 6273
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 17494 6304 17500 6316
rect 17407 6276 17500 6304
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 17753 6307 17811 6313
rect 17753 6304 17765 6307
rect 17604 6276 17765 6304
rect 17604 6236 17632 6276
rect 17753 6273 17765 6276
rect 17799 6273 17811 6307
rect 19794 6304 19800 6316
rect 19755 6276 19800 6304
rect 17753 6267 17811 6273
rect 19794 6264 19800 6276
rect 19852 6264 19858 6316
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6304 19947 6307
rect 20438 6304 20444 6316
rect 19935 6276 20444 6304
rect 19935 6273 19947 6276
rect 19889 6267 19947 6273
rect 20438 6264 20444 6276
rect 20496 6304 20502 6316
rect 20901 6307 20959 6313
rect 20901 6304 20913 6307
rect 20496 6276 20913 6304
rect 20496 6264 20502 6276
rect 20901 6273 20913 6276
rect 20947 6273 20959 6307
rect 22557 6307 22615 6313
rect 22557 6304 22569 6307
rect 20901 6267 20959 6273
rect 22066 6276 22569 6304
rect 19978 6236 19984 6248
rect 17236 6208 17632 6236
rect 19939 6208 19984 6236
rect 14182 6128 14188 6180
rect 14240 6168 14246 6180
rect 14737 6171 14795 6177
rect 14737 6168 14749 6171
rect 14240 6140 14749 6168
rect 14240 6128 14246 6140
rect 14737 6137 14749 6140
rect 14783 6168 14795 6171
rect 15838 6168 15844 6180
rect 14783 6140 15844 6168
rect 14783 6137 14795 6140
rect 14737 6131 14795 6137
rect 15838 6128 15844 6140
rect 15896 6128 15902 6180
rect 17236 6177 17264 6208
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 21082 6236 21088 6248
rect 21043 6208 21088 6236
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 17221 6171 17279 6177
rect 17221 6137 17233 6171
rect 17267 6137 17279 6171
rect 17221 6131 17279 6137
rect 18877 6171 18935 6177
rect 18877 6137 18889 6171
rect 18923 6168 18935 6171
rect 22066 6168 22094 6276
rect 22557 6273 22569 6276
rect 22603 6273 22615 6307
rect 23198 6304 23204 6316
rect 23159 6276 23204 6304
rect 22557 6267 22615 6273
rect 23198 6264 23204 6276
rect 23256 6264 23262 6316
rect 23658 6304 23664 6316
rect 23619 6276 23664 6304
rect 23658 6264 23664 6276
rect 23716 6264 23722 6316
rect 23750 6264 23756 6316
rect 23808 6304 23814 6316
rect 24136 6313 24164 6344
rect 24670 6332 24676 6344
rect 24728 6332 24734 6384
rect 24121 6307 24179 6313
rect 24121 6304 24133 6307
rect 23808 6276 24133 6304
rect 23808 6264 23814 6276
rect 24121 6273 24133 6276
rect 24167 6273 24179 6307
rect 24377 6307 24435 6313
rect 24377 6304 24389 6307
rect 24121 6267 24179 6273
rect 24228 6276 24389 6304
rect 22646 6236 22652 6248
rect 22607 6208 22652 6236
rect 22646 6196 22652 6208
rect 22704 6196 22710 6248
rect 22830 6236 22836 6248
rect 22791 6208 22836 6236
rect 22830 6196 22836 6208
rect 22888 6196 22894 6248
rect 24228 6236 24256 6276
rect 24377 6273 24389 6276
rect 24423 6273 24435 6307
rect 24377 6267 24435 6273
rect 23860 6208 24256 6236
rect 23860 6177 23888 6208
rect 18923 6140 22094 6168
rect 23845 6171 23903 6177
rect 18923 6137 18935 6140
rect 18877 6131 18935 6137
rect 23845 6137 23857 6171
rect 23891 6137 23903 6171
rect 23845 6131 23903 6137
rect 15654 6100 15660 6112
rect 15615 6072 15660 6100
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 18138 6060 18144 6112
rect 18196 6100 18202 6112
rect 18892 6100 18920 6131
rect 18196 6072 18920 6100
rect 19429 6103 19487 6109
rect 18196 6060 18202 6072
rect 19429 6069 19441 6103
rect 19475 6100 19487 6103
rect 19702 6100 19708 6112
rect 19475 6072 19708 6100
rect 19475 6069 19487 6072
rect 19429 6063 19487 6069
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 20441 6103 20499 6109
rect 20441 6069 20453 6103
rect 20487 6100 20499 6103
rect 20622 6100 20628 6112
rect 20487 6072 20628 6100
rect 20487 6069 20499 6072
rect 20441 6063 20499 6069
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 22186 6100 22192 6112
rect 22147 6072 22192 6100
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 23290 6060 23296 6112
rect 23348 6100 23354 6112
rect 23385 6103 23443 6109
rect 23385 6100 23397 6103
rect 23348 6072 23397 6100
rect 23348 6060 23354 6072
rect 23385 6069 23397 6072
rect 23431 6069 23443 6103
rect 23385 6063 23443 6069
rect 1104 6010 28888 6032
rect 1104 5958 5582 6010
rect 5634 5958 5646 6010
rect 5698 5958 5710 6010
rect 5762 5958 5774 6010
rect 5826 5958 5838 6010
rect 5890 5958 14846 6010
rect 14898 5958 14910 6010
rect 14962 5958 14974 6010
rect 15026 5958 15038 6010
rect 15090 5958 15102 6010
rect 15154 5958 24110 6010
rect 24162 5958 24174 6010
rect 24226 5958 24238 6010
rect 24290 5958 24302 6010
rect 24354 5958 24366 6010
rect 24418 5958 28888 6010
rect 1104 5936 28888 5958
rect 17678 5896 17684 5908
rect 17639 5868 17684 5896
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 19334 5896 19340 5908
rect 19295 5868 19340 5896
rect 19334 5856 19340 5868
rect 19392 5856 19398 5908
rect 21913 5899 21971 5905
rect 21913 5865 21925 5899
rect 21959 5896 21971 5899
rect 22094 5896 22100 5908
rect 21959 5868 22100 5896
rect 21959 5865 21971 5868
rect 21913 5859 21971 5865
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 22189 5899 22247 5905
rect 22189 5865 22201 5899
rect 22235 5896 22247 5899
rect 22646 5896 22652 5908
rect 22235 5868 22652 5896
rect 22235 5865 22247 5868
rect 22189 5859 22247 5865
rect 22646 5856 22652 5868
rect 22704 5856 22710 5908
rect 16850 5788 16856 5840
rect 16908 5828 16914 5840
rect 17221 5831 17279 5837
rect 17221 5828 17233 5831
rect 16908 5800 17233 5828
rect 16908 5788 16914 5800
rect 17221 5797 17233 5800
rect 17267 5828 17279 5831
rect 19794 5828 19800 5840
rect 17267 5800 19800 5828
rect 17267 5797 17279 5800
rect 17221 5791 17279 5797
rect 19794 5788 19800 5800
rect 19852 5788 19858 5840
rect 13722 5760 13728 5772
rect 13683 5732 13728 5760
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 18138 5760 18144 5772
rect 18099 5732 18144 5760
rect 18138 5720 18144 5732
rect 18196 5720 18202 5772
rect 18322 5760 18328 5772
rect 18283 5732 18328 5760
rect 18322 5720 18328 5732
rect 18380 5720 18386 5772
rect 19981 5763 20039 5769
rect 19981 5729 19993 5763
rect 20027 5729 20039 5763
rect 19981 5723 20039 5729
rect 13446 5692 13452 5704
rect 13504 5701 13510 5704
rect 13416 5664 13452 5692
rect 13446 5652 13452 5664
rect 13504 5655 13516 5701
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5692 15899 5695
rect 17494 5692 17500 5704
rect 15887 5664 17500 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 13504 5652 13510 5655
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 19702 5692 19708 5704
rect 19663 5664 19708 5692
rect 19702 5652 19708 5664
rect 19760 5652 19766 5704
rect 19996 5692 20024 5723
rect 20346 5720 20352 5772
rect 20404 5760 20410 5772
rect 20533 5763 20591 5769
rect 20533 5760 20545 5763
rect 20404 5732 20545 5760
rect 20404 5720 20410 5732
rect 20533 5729 20545 5732
rect 20579 5729 20591 5763
rect 20533 5723 20591 5729
rect 23569 5763 23627 5769
rect 23569 5729 23581 5763
rect 23615 5760 23627 5763
rect 23750 5760 23756 5772
rect 23615 5732 23756 5760
rect 23615 5729 23627 5732
rect 23569 5723 23627 5729
rect 23750 5720 23756 5732
rect 23808 5720 23814 5772
rect 21082 5692 21088 5704
rect 19996 5664 21088 5692
rect 21082 5652 21088 5664
rect 21140 5692 21146 5704
rect 22278 5692 22284 5704
rect 21140 5664 22284 5692
rect 21140 5652 21146 5664
rect 22278 5652 22284 5664
rect 22336 5692 22342 5704
rect 22738 5692 22744 5704
rect 22336 5664 22744 5692
rect 22336 5652 22342 5664
rect 22738 5652 22744 5664
rect 22796 5652 22802 5704
rect 23290 5652 23296 5704
rect 23348 5701 23354 5704
rect 23348 5692 23360 5701
rect 28074 5692 28080 5704
rect 23348 5664 23393 5692
rect 28035 5664 28080 5692
rect 23348 5655 23360 5664
rect 23348 5652 23354 5655
rect 28074 5652 28080 5664
rect 28132 5652 28138 5704
rect 15654 5584 15660 5636
rect 15712 5624 15718 5636
rect 16086 5627 16144 5633
rect 16086 5624 16098 5627
rect 15712 5596 16098 5624
rect 15712 5584 15718 5596
rect 16086 5593 16098 5596
rect 16132 5593 16144 5627
rect 16086 5587 16144 5593
rect 19797 5627 19855 5633
rect 19797 5593 19809 5627
rect 19843 5624 19855 5627
rect 19886 5624 19892 5636
rect 19843 5596 19892 5624
rect 19843 5593 19855 5596
rect 19797 5587 19855 5593
rect 19886 5584 19892 5596
rect 19944 5584 19950 5636
rect 20806 5633 20812 5636
rect 20800 5587 20812 5633
rect 20864 5624 20870 5636
rect 20864 5596 20900 5624
rect 20806 5584 20812 5587
rect 20864 5584 20870 5596
rect 12342 5556 12348 5568
rect 12303 5528 12348 5556
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 18012 5528 18061 5556
rect 18012 5516 18018 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 28258 5556 28264 5568
rect 28219 5528 28264 5556
rect 18049 5519 18107 5525
rect 28258 5516 28264 5528
rect 28316 5516 28322 5568
rect 1104 5466 28888 5488
rect 1104 5414 10214 5466
rect 10266 5414 10278 5466
rect 10330 5414 10342 5466
rect 10394 5414 10406 5466
rect 10458 5414 10470 5466
rect 10522 5414 19478 5466
rect 19530 5414 19542 5466
rect 19594 5414 19606 5466
rect 19658 5414 19670 5466
rect 19722 5414 19734 5466
rect 19786 5414 28888 5466
rect 1104 5392 28888 5414
rect 17589 5355 17647 5361
rect 17589 5321 17601 5355
rect 17635 5352 17647 5355
rect 17954 5352 17960 5364
rect 17635 5324 17960 5352
rect 17635 5321 17647 5324
rect 17589 5315 17647 5321
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 20806 5352 20812 5364
rect 20767 5324 20812 5352
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 22186 5352 22192 5364
rect 22147 5324 22192 5352
rect 22186 5312 22192 5324
rect 22244 5312 22250 5364
rect 22557 5355 22615 5361
rect 22557 5321 22569 5355
rect 22603 5352 22615 5355
rect 23198 5352 23204 5364
rect 22603 5324 23204 5352
rect 22603 5321 22615 5324
rect 22557 5315 22615 5321
rect 23198 5312 23204 5324
rect 23256 5312 23262 5364
rect 20346 5284 20352 5296
rect 18984 5256 20352 5284
rect 18984 5225 19012 5256
rect 20346 5244 20352 5256
rect 20404 5244 20410 5296
rect 22094 5244 22100 5296
rect 22152 5284 22158 5296
rect 22152 5256 22197 5284
rect 22152 5244 22158 5256
rect 19242 5225 19248 5228
rect 18969 5219 19027 5225
rect 18969 5185 18981 5219
rect 19015 5185 19027 5219
rect 19236 5216 19248 5225
rect 19203 5188 19248 5216
rect 18969 5179 19027 5185
rect 19236 5179 19248 5188
rect 19242 5176 19248 5179
rect 19300 5176 19306 5228
rect 20622 5216 20628 5228
rect 20583 5188 20628 5216
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 22005 5151 22063 5157
rect 22005 5117 22017 5151
rect 22051 5148 22063 5151
rect 22278 5148 22284 5160
rect 22051 5120 22284 5148
rect 22051 5117 22063 5120
rect 22005 5111 22063 5117
rect 22278 5108 22284 5120
rect 22336 5108 22342 5160
rect 20349 5083 20407 5089
rect 20349 5049 20361 5083
rect 20395 5080 20407 5083
rect 20438 5080 20444 5092
rect 20395 5052 20444 5080
rect 20395 5049 20407 5052
rect 20349 5043 20407 5049
rect 20438 5040 20444 5052
rect 20496 5040 20502 5092
rect 1104 4922 28888 4944
rect 1104 4870 5582 4922
rect 5634 4870 5646 4922
rect 5698 4870 5710 4922
rect 5762 4870 5774 4922
rect 5826 4870 5838 4922
rect 5890 4870 14846 4922
rect 14898 4870 14910 4922
rect 14962 4870 14974 4922
rect 15026 4870 15038 4922
rect 15090 4870 15102 4922
rect 15154 4870 24110 4922
rect 24162 4870 24174 4922
rect 24226 4870 24238 4922
rect 24290 4870 24302 4922
rect 24354 4870 24366 4922
rect 24418 4870 28888 4922
rect 1104 4848 28888 4870
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 27893 4607 27951 4613
rect 27893 4573 27905 4607
rect 27939 4604 27951 4607
rect 28350 4604 28356 4616
rect 27939 4576 28356 4604
rect 27939 4573 27951 4576
rect 27893 4567 27951 4573
rect 28350 4564 28356 4576
rect 28408 4564 28414 4616
rect 19058 4496 19064 4548
rect 19116 4536 19122 4548
rect 19116 4508 28212 4536
rect 19116 4496 19122 4508
rect 28184 4477 28212 4508
rect 28169 4471 28227 4477
rect 28169 4437 28181 4471
rect 28215 4437 28227 4471
rect 28169 4431 28227 4437
rect 1104 4378 28888 4400
rect 1104 4326 10214 4378
rect 10266 4326 10278 4378
rect 10330 4326 10342 4378
rect 10394 4326 10406 4378
rect 10458 4326 10470 4378
rect 10522 4326 19478 4378
rect 19530 4326 19542 4378
rect 19594 4326 19606 4378
rect 19658 4326 19670 4378
rect 19722 4326 19734 4378
rect 19786 4326 28888 4378
rect 1104 4304 28888 4326
rect 1104 3834 28888 3856
rect 1104 3782 5582 3834
rect 5634 3782 5646 3834
rect 5698 3782 5710 3834
rect 5762 3782 5774 3834
rect 5826 3782 5838 3834
rect 5890 3782 14846 3834
rect 14898 3782 14910 3834
rect 14962 3782 14974 3834
rect 15026 3782 15038 3834
rect 15090 3782 15102 3834
rect 15154 3782 24110 3834
rect 24162 3782 24174 3834
rect 24226 3782 24238 3834
rect 24290 3782 24302 3834
rect 24354 3782 24366 3834
rect 24418 3782 28888 3834
rect 1104 3760 28888 3782
rect 1104 3290 28888 3312
rect 1104 3238 10214 3290
rect 10266 3238 10278 3290
rect 10330 3238 10342 3290
rect 10394 3238 10406 3290
rect 10458 3238 10470 3290
rect 10522 3238 19478 3290
rect 19530 3238 19542 3290
rect 19594 3238 19606 3290
rect 19658 3238 19670 3290
rect 19722 3238 19734 3290
rect 19786 3238 28888 3290
rect 1104 3216 28888 3238
rect 16574 3136 16580 3188
rect 16632 3176 16638 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 16632 3148 16865 3176
rect 16632 3136 16638 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 17402 3136 17408 3188
rect 17460 3176 17466 3188
rect 17957 3179 18015 3185
rect 17957 3176 17969 3179
rect 17460 3148 17969 3176
rect 17460 3136 17466 3148
rect 17957 3145 17969 3148
rect 18003 3145 18015 3179
rect 17957 3139 18015 3145
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 12342 3040 12348 3052
rect 1719 3012 12348 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 17310 3040 17316 3052
rect 17271 3012 17316 3040
rect 17310 3000 17316 3012
rect 17368 3040 17374 3052
rect 17589 3043 17647 3049
rect 17589 3040 17601 3043
rect 17368 3012 17601 3040
rect 17368 3000 17374 3012
rect 17589 3009 17601 3012
rect 17635 3009 17647 3043
rect 17589 3003 17647 3009
rect 17773 3043 17831 3049
rect 17773 3009 17785 3043
rect 17819 3040 17831 3043
rect 24578 3040 24584 3052
rect 17819 3012 24584 3040
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 1486 2836 1492 2848
rect 1447 2808 1492 2836
rect 1486 2796 1492 2808
rect 1544 2796 1550 2848
rect 17221 2839 17279 2845
rect 17221 2805 17233 2839
rect 17267 2836 17279 2839
rect 17788 2836 17816 3003
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 28350 2836 28356 2848
rect 17267 2808 17816 2836
rect 28311 2808 28356 2836
rect 17267 2805 17279 2808
rect 17221 2799 17279 2805
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 1104 2746 28888 2768
rect 1104 2694 5582 2746
rect 5634 2694 5646 2746
rect 5698 2694 5710 2746
rect 5762 2694 5774 2746
rect 5826 2694 5838 2746
rect 5890 2694 14846 2746
rect 14898 2694 14910 2746
rect 14962 2694 14974 2746
rect 15026 2694 15038 2746
rect 15090 2694 15102 2746
rect 15154 2694 24110 2746
rect 24162 2694 24174 2746
rect 24226 2694 24238 2746
rect 24290 2694 24302 2746
rect 24354 2694 24366 2746
rect 24418 2694 28888 2746
rect 1104 2672 28888 2694
rect 5629 2635 5687 2641
rect 5629 2601 5641 2635
rect 5675 2632 5687 2635
rect 9214 2632 9220 2644
rect 5675 2604 9220 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 15657 2635 15715 2641
rect 15657 2601 15669 2635
rect 15703 2632 15715 2635
rect 15838 2632 15844 2644
rect 15703 2604 15844 2632
rect 15703 2601 15715 2604
rect 15657 2595 15715 2601
rect 15838 2592 15844 2604
rect 15896 2592 15902 2644
rect 18046 2592 18052 2644
rect 18104 2632 18110 2644
rect 18141 2635 18199 2641
rect 18141 2632 18153 2635
rect 18104 2604 18153 2632
rect 18104 2592 18110 2604
rect 18141 2601 18153 2604
rect 18187 2601 18199 2635
rect 24578 2632 24584 2644
rect 24539 2604 24584 2632
rect 18141 2595 18199 2601
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 2869 2567 2927 2573
rect 2869 2533 2881 2567
rect 2915 2564 2927 2567
rect 8021 2567 8079 2573
rect 2915 2536 6914 2564
rect 2915 2533 2927 2536
rect 2869 2527 2927 2533
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2590 2388 2596 2440
rect 2648 2428 2654 2440
rect 2685 2431 2743 2437
rect 2685 2428 2697 2431
rect 2648 2400 2697 2428
rect 2648 2388 2654 2400
rect 2685 2397 2697 2400
rect 2731 2428 2743 2431
rect 3237 2431 3295 2437
rect 3237 2428 3249 2431
rect 2731 2400 3249 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 3237 2397 3249 2400
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6512 2400 6561 2428
rect 6512 2388 6518 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 5184 2332 5365 2360
rect 5184 2304 5212 2332
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 6886 2360 6914 2536
rect 8021 2533 8033 2567
rect 8067 2533 8079 2567
rect 8021 2527 8079 2533
rect 8036 2496 8064 2527
rect 15930 2524 15936 2576
rect 15988 2564 15994 2576
rect 15988 2536 20760 2564
rect 15988 2524 15994 2536
rect 17310 2496 17316 2508
rect 8036 2468 17316 2496
rect 17310 2456 17316 2468
rect 17368 2456 17374 2508
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7800 2400 7849 2428
rect 7800 2388 7806 2400
rect 7837 2397 7849 2400
rect 7883 2428 7895 2431
rect 8297 2431 8355 2437
rect 8297 2428 8309 2431
rect 7883 2400 8309 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 8297 2397 8309 2400
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 10134 2388 10140 2440
rect 10192 2428 10198 2440
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 10192 2400 10425 2428
rect 10192 2388 10198 2400
rect 10413 2397 10425 2400
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 15841 2431 15899 2437
rect 15841 2428 15853 2431
rect 15528 2400 15853 2428
rect 15528 2388 15534 2400
rect 15841 2397 15853 2400
rect 15887 2428 15899 2431
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15887 2400 16129 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 20732 2437 20760 2536
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 18104 2400 18337 2428
rect 18104 2388 18110 2400
rect 18325 2397 18337 2400
rect 18371 2428 18383 2431
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 18371 2400 18613 2428
rect 18371 2397 18383 2400
rect 18325 2391 18383 2397
rect 18601 2397 18613 2400
rect 18647 2397 18659 2431
rect 18601 2391 18659 2397
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24544 2400 24777 2428
rect 24544 2388 24550 2400
rect 24765 2397 24777 2400
rect 24811 2428 24823 2431
rect 25041 2431 25099 2437
rect 25041 2428 25053 2431
rect 24811 2400 25053 2428
rect 24811 2397 24823 2400
rect 24765 2391 24823 2397
rect 25041 2397 25053 2400
rect 25087 2397 25099 2431
rect 25041 2391 25099 2397
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 25832 2400 25881 2428
rect 25832 2388 25838 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 27522 2388 27528 2440
rect 27580 2428 27586 2440
rect 28353 2431 28411 2437
rect 28353 2428 28365 2431
rect 27580 2400 28365 2428
rect 27580 2388 27586 2400
rect 28353 2397 28365 2400
rect 28399 2397 28411 2431
rect 28353 2391 28411 2397
rect 12618 2360 12624 2372
rect 6886 2332 12624 2360
rect 5353 2323 5411 2329
rect 12618 2320 12624 2332
rect 12676 2320 12682 2372
rect 1486 2292 1492 2304
rect 1447 2264 1492 2292
rect 1486 2252 1492 2264
rect 1544 2252 1550 2304
rect 4985 2295 5043 2301
rect 4985 2261 4997 2295
rect 5031 2292 5043 2295
rect 5166 2292 5172 2304
rect 5031 2264 5172 2292
rect 5031 2261 5043 2264
rect 4985 2255 5043 2261
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20680 2264 20913 2292
rect 20680 2252 20686 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 1104 2202 28888 2224
rect 1104 2150 10214 2202
rect 10266 2150 10278 2202
rect 10330 2150 10342 2202
rect 10394 2150 10406 2202
rect 10458 2150 10470 2202
rect 10522 2150 19478 2202
rect 19530 2150 19542 2202
rect 19594 2150 19606 2202
rect 19658 2150 19670 2202
rect 19722 2150 19734 2202
rect 19786 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 5582 27718 5634 27770
rect 5646 27718 5698 27770
rect 5710 27718 5762 27770
rect 5774 27718 5826 27770
rect 5838 27718 5890 27770
rect 14846 27718 14898 27770
rect 14910 27718 14962 27770
rect 14974 27718 15026 27770
rect 15038 27718 15090 27770
rect 15102 27718 15154 27770
rect 24110 27718 24162 27770
rect 24174 27718 24226 27770
rect 24238 27718 24290 27770
rect 24302 27718 24354 27770
rect 24366 27718 24418 27770
rect 2044 27591 2096 27600
rect 2044 27557 2053 27591
rect 2053 27557 2087 27591
rect 2087 27557 2096 27591
rect 2044 27548 2096 27557
rect 3332 27591 3384 27600
rect 3332 27557 3341 27591
rect 3341 27557 3375 27591
rect 3375 27557 3384 27591
rect 3332 27548 3384 27557
rect 6184 27548 6236 27600
rect 12348 27591 12400 27600
rect 12348 27557 12357 27591
rect 12357 27557 12391 27591
rect 12391 27557 12400 27591
rect 12348 27548 12400 27557
rect 13820 27548 13872 27600
rect 14740 27548 14792 27600
rect 16120 27548 16172 27600
rect 18696 27548 18748 27600
rect 19984 27548 20036 27600
rect 21272 27548 21324 27600
rect 25136 27548 25188 27600
rect 26516 27591 26568 27600
rect 26516 27557 26525 27591
rect 26525 27557 26559 27591
rect 26559 27557 26568 27591
rect 26516 27548 26568 27557
rect 28080 27591 28132 27600
rect 28080 27557 28089 27591
rect 28089 27557 28123 27591
rect 28123 27557 28132 27591
rect 28080 27548 28132 27557
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 21088 27480 21140 27532
rect 13728 27412 13780 27464
rect 14648 27412 14700 27464
rect 16304 27412 16356 27464
rect 18052 27412 18104 27464
rect 4436 27387 4488 27396
rect 4436 27353 4445 27387
rect 4445 27353 4479 27387
rect 4479 27353 4488 27387
rect 4436 27344 4488 27353
rect 20628 27412 20680 27464
rect 27896 27455 27948 27464
rect 27896 27421 27905 27455
rect 27905 27421 27939 27455
rect 27939 27421 27948 27455
rect 27896 27412 27948 27421
rect 20996 27344 21048 27396
rect 25872 27344 25924 27396
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 17960 27319 18012 27328
rect 17960 27285 17969 27319
rect 17969 27285 18003 27319
rect 18003 27285 18012 27319
rect 17960 27276 18012 27285
rect 20260 27276 20312 27328
rect 27344 27319 27396 27328
rect 27344 27285 27353 27319
rect 27353 27285 27387 27319
rect 27387 27285 27396 27319
rect 27344 27276 27396 27285
rect 10214 27174 10266 27226
rect 10278 27174 10330 27226
rect 10342 27174 10394 27226
rect 10406 27174 10458 27226
rect 10470 27174 10522 27226
rect 19478 27174 19530 27226
rect 19542 27174 19594 27226
rect 19606 27174 19658 27226
rect 19670 27174 19722 27226
rect 19734 27174 19786 27226
rect 1492 27072 1544 27124
rect 14648 27115 14700 27124
rect 14648 27081 14657 27115
rect 14657 27081 14691 27115
rect 14691 27081 14700 27115
rect 14648 27072 14700 27081
rect 16304 27115 16356 27124
rect 16304 27081 16313 27115
rect 16313 27081 16347 27115
rect 16347 27081 16356 27115
rect 16304 27072 16356 27081
rect 1400 26979 1452 26988
rect 1400 26945 1409 26979
rect 1409 26945 1443 26979
rect 1443 26945 1452 26979
rect 1400 26936 1452 26945
rect 14740 27004 14792 27056
rect 14004 26936 14056 26988
rect 15384 27004 15436 27056
rect 17960 27004 18012 27056
rect 23848 27072 23900 27124
rect 27896 27072 27948 27124
rect 20444 26936 20496 26988
rect 21732 26936 21784 26988
rect 17500 26911 17552 26920
rect 17500 26877 17509 26911
rect 17509 26877 17543 26911
rect 17543 26877 17552 26911
rect 17500 26868 17552 26877
rect 19524 26800 19576 26852
rect 19064 26732 19116 26784
rect 19340 26732 19392 26784
rect 23388 26868 23440 26920
rect 26148 27004 26200 27056
rect 25504 26979 25556 26988
rect 25504 26945 25538 26979
rect 25538 26945 25556 26979
rect 25504 26936 25556 26945
rect 26700 26868 26752 26920
rect 24676 26843 24728 26852
rect 24676 26809 24685 26843
rect 24685 26809 24719 26843
rect 24719 26809 24728 26843
rect 24676 26800 24728 26809
rect 22192 26732 22244 26784
rect 28356 26775 28408 26784
rect 28356 26741 28365 26775
rect 28365 26741 28399 26775
rect 28399 26741 28408 26775
rect 28356 26732 28408 26741
rect 5582 26630 5634 26682
rect 5646 26630 5698 26682
rect 5710 26630 5762 26682
rect 5774 26630 5826 26682
rect 5838 26630 5890 26682
rect 14846 26630 14898 26682
rect 14910 26630 14962 26682
rect 14974 26630 15026 26682
rect 15038 26630 15090 26682
rect 15102 26630 15154 26682
rect 24110 26630 24162 26682
rect 24174 26630 24226 26682
rect 24238 26630 24290 26682
rect 24302 26630 24354 26682
rect 24366 26630 24418 26682
rect 18052 26571 18104 26580
rect 18052 26537 18061 26571
rect 18061 26537 18095 26571
rect 18095 26537 18104 26571
rect 18052 26528 18104 26537
rect 18236 26571 18288 26580
rect 18236 26537 18245 26571
rect 18245 26537 18279 26571
rect 18279 26537 18288 26571
rect 18236 26528 18288 26537
rect 20444 26571 20496 26580
rect 20444 26537 20453 26571
rect 20453 26537 20487 26571
rect 20487 26537 20496 26571
rect 20444 26528 20496 26537
rect 27528 26528 27580 26580
rect 21732 26503 21784 26512
rect 21732 26469 21741 26503
rect 21741 26469 21775 26503
rect 21775 26469 21784 26503
rect 21732 26460 21784 26469
rect 1676 26367 1728 26376
rect 1676 26333 1685 26367
rect 1685 26333 1719 26367
rect 1719 26333 1728 26367
rect 1676 26324 1728 26333
rect 17500 26324 17552 26376
rect 19340 26324 19392 26376
rect 1768 26256 1820 26308
rect 16672 26256 16724 26308
rect 18328 26256 18380 26308
rect 18420 26299 18472 26308
rect 18420 26265 18429 26299
rect 18429 26265 18463 26299
rect 18463 26265 18472 26299
rect 19524 26367 19576 26376
rect 19524 26333 19533 26367
rect 19533 26333 19567 26367
rect 19567 26333 19576 26367
rect 19524 26324 19576 26333
rect 19984 26324 20036 26376
rect 20996 26367 21048 26376
rect 18420 26256 18472 26265
rect 19892 26256 19944 26308
rect 20260 26299 20312 26308
rect 20260 26265 20285 26299
rect 20285 26265 20312 26299
rect 20996 26333 21005 26367
rect 21005 26333 21039 26367
rect 21039 26333 21048 26367
rect 20996 26324 21048 26333
rect 22192 26324 22244 26376
rect 28356 26367 28408 26376
rect 28356 26333 28365 26367
rect 28365 26333 28399 26367
rect 28399 26333 28408 26367
rect 28356 26324 28408 26333
rect 20260 26256 20312 26265
rect 25136 26299 25188 26308
rect 25136 26265 25145 26299
rect 25145 26265 25179 26299
rect 25179 26265 25188 26299
rect 25136 26256 25188 26265
rect 26700 26256 26752 26308
rect 17592 26188 17644 26240
rect 21088 26231 21140 26240
rect 21088 26197 21097 26231
rect 21097 26197 21131 26231
rect 21131 26197 21140 26231
rect 21088 26188 21140 26197
rect 21916 26231 21968 26240
rect 21916 26197 21943 26231
rect 21943 26197 21968 26231
rect 21916 26188 21968 26197
rect 10214 26086 10266 26138
rect 10278 26086 10330 26138
rect 10342 26086 10394 26138
rect 10406 26086 10458 26138
rect 10470 26086 10522 26138
rect 19478 26086 19530 26138
rect 19542 26086 19594 26138
rect 19606 26086 19658 26138
rect 19670 26086 19722 26138
rect 19734 26086 19786 26138
rect 16672 26027 16724 26036
rect 16672 25993 16681 26027
rect 16681 25993 16715 26027
rect 16715 25993 16724 26027
rect 16672 25984 16724 25993
rect 17316 25984 17368 26036
rect 18236 25984 18288 26036
rect 18512 25984 18564 26036
rect 20260 25984 20312 26036
rect 21456 25984 21508 26036
rect 21916 25984 21968 26036
rect 15476 25891 15528 25900
rect 15476 25857 15485 25891
rect 15485 25857 15519 25891
rect 15519 25857 15528 25891
rect 15476 25848 15528 25857
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 17316 25891 17368 25900
rect 17316 25857 17325 25891
rect 17325 25857 17359 25891
rect 17359 25857 17368 25891
rect 17316 25848 17368 25857
rect 17500 25848 17552 25900
rect 17684 25848 17736 25900
rect 19156 25916 19208 25968
rect 18696 25891 18748 25900
rect 18696 25857 18706 25891
rect 18706 25857 18740 25891
rect 18740 25857 18748 25891
rect 18696 25848 18748 25857
rect 19064 25848 19116 25900
rect 20720 25916 20772 25968
rect 18328 25780 18380 25832
rect 19156 25780 19208 25832
rect 15292 25687 15344 25696
rect 15292 25653 15301 25687
rect 15301 25653 15335 25687
rect 15335 25653 15344 25687
rect 15292 25644 15344 25653
rect 17224 25644 17276 25696
rect 18696 25712 18748 25764
rect 18972 25712 19024 25764
rect 19984 25780 20036 25832
rect 20260 25780 20312 25832
rect 20996 25848 21048 25900
rect 22192 25916 22244 25968
rect 25688 25959 25740 25968
rect 22100 25891 22152 25900
rect 22100 25857 22109 25891
rect 22109 25857 22143 25891
rect 22143 25857 22152 25891
rect 22100 25848 22152 25857
rect 25688 25925 25697 25959
rect 25697 25925 25731 25959
rect 25731 25925 25740 25959
rect 25688 25916 25740 25925
rect 23756 25891 23808 25900
rect 23756 25857 23790 25891
rect 23790 25857 23808 25891
rect 25412 25891 25464 25900
rect 21088 25780 21140 25832
rect 23756 25848 23808 25857
rect 25412 25857 25421 25891
rect 25421 25857 25455 25891
rect 25455 25857 25464 25891
rect 25412 25848 25464 25857
rect 25596 25891 25648 25900
rect 25596 25857 25605 25891
rect 25605 25857 25639 25891
rect 25639 25857 25648 25891
rect 25596 25848 25648 25857
rect 25780 25891 25832 25900
rect 25780 25857 25789 25891
rect 25789 25857 25823 25891
rect 25823 25857 25832 25891
rect 25780 25848 25832 25857
rect 23388 25780 23440 25832
rect 20536 25712 20588 25764
rect 20628 25712 20680 25764
rect 22100 25712 22152 25764
rect 18604 25644 18656 25696
rect 19524 25644 19576 25696
rect 24768 25644 24820 25696
rect 25964 25687 26016 25696
rect 25964 25653 25973 25687
rect 25973 25653 26007 25687
rect 26007 25653 26016 25687
rect 25964 25644 26016 25653
rect 5582 25542 5634 25594
rect 5646 25542 5698 25594
rect 5710 25542 5762 25594
rect 5774 25542 5826 25594
rect 5838 25542 5890 25594
rect 14846 25542 14898 25594
rect 14910 25542 14962 25594
rect 14974 25542 15026 25594
rect 15038 25542 15090 25594
rect 15102 25542 15154 25594
rect 24110 25542 24162 25594
rect 24174 25542 24226 25594
rect 24238 25542 24290 25594
rect 24302 25542 24354 25594
rect 24366 25542 24418 25594
rect 17132 25483 17184 25492
rect 17132 25449 17141 25483
rect 17141 25449 17175 25483
rect 17175 25449 17184 25483
rect 17132 25440 17184 25449
rect 17224 25483 17276 25492
rect 17224 25449 17233 25483
rect 17233 25449 17267 25483
rect 17267 25449 17276 25483
rect 17224 25440 17276 25449
rect 23756 25440 23808 25492
rect 25688 25440 25740 25492
rect 16580 25415 16632 25424
rect 16580 25381 16589 25415
rect 16589 25381 16623 25415
rect 16623 25381 16632 25415
rect 16580 25372 16632 25381
rect 16856 25372 16908 25424
rect 14740 25304 14792 25356
rect 18328 25372 18380 25424
rect 19064 25372 19116 25424
rect 22008 25415 22060 25424
rect 15292 25168 15344 25220
rect 16672 25279 16724 25288
rect 16672 25245 16681 25279
rect 16681 25245 16715 25279
rect 16715 25245 16724 25279
rect 16672 25236 16724 25245
rect 17408 25236 17460 25288
rect 18512 25304 18564 25356
rect 22008 25381 22017 25415
rect 22017 25381 22051 25415
rect 22051 25381 22060 25415
rect 22008 25372 22060 25381
rect 19524 25236 19576 25288
rect 20720 25304 20772 25356
rect 20904 25236 20956 25288
rect 21088 25279 21140 25288
rect 21088 25245 21097 25279
rect 21097 25245 21131 25279
rect 21131 25245 21140 25279
rect 21088 25236 21140 25245
rect 22376 25304 22428 25356
rect 24768 25304 24820 25356
rect 25780 25304 25832 25356
rect 21456 25279 21508 25288
rect 21456 25245 21465 25279
rect 21465 25245 21499 25279
rect 21499 25245 21508 25279
rect 21456 25236 21508 25245
rect 22652 25236 22704 25288
rect 23388 25279 23440 25288
rect 23388 25245 23397 25279
rect 23397 25245 23431 25279
rect 23431 25245 23440 25279
rect 23388 25236 23440 25245
rect 24860 25279 24912 25288
rect 16212 25143 16264 25152
rect 16212 25109 16221 25143
rect 16221 25109 16255 25143
rect 16255 25109 16264 25143
rect 16212 25100 16264 25109
rect 16672 25100 16724 25152
rect 17500 25100 17552 25152
rect 19064 25100 19116 25152
rect 19248 25143 19300 25152
rect 19248 25109 19257 25143
rect 19257 25109 19291 25143
rect 19291 25109 19300 25143
rect 19248 25100 19300 25109
rect 20168 25168 20220 25220
rect 20352 25168 20404 25220
rect 21272 25100 21324 25152
rect 24860 25245 24869 25279
rect 24869 25245 24903 25279
rect 24903 25245 24912 25279
rect 24860 25236 24912 25245
rect 26148 25236 26200 25288
rect 25412 25168 25464 25220
rect 25780 25168 25832 25220
rect 25964 25168 26016 25220
rect 10214 24998 10266 25050
rect 10278 24998 10330 25050
rect 10342 24998 10394 25050
rect 10406 24998 10458 25050
rect 10470 24998 10522 25050
rect 19478 24998 19530 25050
rect 19542 24998 19594 25050
rect 19606 24998 19658 25050
rect 19670 24998 19722 25050
rect 19734 24998 19786 25050
rect 15476 24896 15528 24948
rect 19064 24939 19116 24948
rect 19064 24905 19073 24939
rect 19073 24905 19107 24939
rect 19107 24905 19116 24939
rect 19064 24896 19116 24905
rect 19156 24896 19208 24948
rect 19984 24896 20036 24948
rect 20904 24896 20956 24948
rect 21272 24939 21324 24948
rect 21272 24905 21281 24939
rect 21281 24905 21315 24939
rect 21315 24905 21324 24939
rect 21272 24896 21324 24905
rect 15476 24760 15528 24812
rect 16304 24828 16356 24880
rect 18420 24828 18472 24880
rect 16580 24760 16632 24812
rect 15752 24692 15804 24744
rect 15844 24692 15896 24744
rect 16212 24692 16264 24744
rect 17776 24760 17828 24812
rect 19708 24760 19760 24812
rect 20168 24828 20220 24880
rect 22376 24896 22428 24948
rect 25596 24896 25648 24948
rect 23020 24871 23072 24880
rect 20536 24803 20588 24812
rect 16856 24735 16908 24744
rect 16856 24701 16865 24735
rect 16865 24701 16899 24735
rect 16899 24701 16908 24735
rect 16856 24692 16908 24701
rect 16488 24624 16540 24676
rect 17408 24692 17460 24744
rect 18328 24735 18380 24744
rect 18328 24701 18337 24735
rect 18337 24701 18371 24735
rect 18371 24701 18380 24735
rect 18328 24692 18380 24701
rect 18420 24692 18472 24744
rect 20536 24769 20545 24803
rect 20545 24769 20579 24803
rect 20579 24769 20588 24803
rect 20536 24760 20588 24769
rect 20628 24803 20680 24812
rect 20628 24769 20637 24803
rect 20637 24769 20671 24803
rect 20671 24769 20680 24803
rect 20628 24760 20680 24769
rect 22192 24803 22244 24812
rect 22192 24769 22201 24803
rect 22201 24769 22235 24803
rect 22235 24769 22244 24803
rect 22192 24760 22244 24769
rect 22376 24760 22428 24812
rect 23020 24837 23029 24871
rect 23029 24837 23063 24871
rect 23063 24837 23072 24871
rect 23020 24828 23072 24837
rect 24768 24760 24820 24812
rect 25688 24760 25740 24812
rect 28264 24803 28316 24812
rect 28264 24769 28273 24803
rect 28273 24769 28307 24803
rect 28307 24769 28316 24803
rect 28264 24760 28316 24769
rect 20352 24735 20404 24744
rect 19892 24624 19944 24676
rect 15200 24599 15252 24608
rect 15200 24565 15209 24599
rect 15209 24565 15243 24599
rect 15243 24565 15252 24599
rect 15200 24556 15252 24565
rect 17040 24556 17092 24608
rect 18604 24556 18656 24608
rect 19064 24556 19116 24608
rect 20352 24701 20361 24735
rect 20361 24701 20395 24735
rect 20395 24701 20404 24735
rect 20352 24692 20404 24701
rect 22468 24624 22520 24676
rect 23020 24624 23072 24676
rect 25136 24624 25188 24676
rect 20444 24599 20496 24608
rect 20444 24565 20453 24599
rect 20453 24565 20487 24599
rect 20487 24565 20496 24599
rect 20444 24556 20496 24565
rect 21824 24599 21876 24608
rect 21824 24565 21833 24599
rect 21833 24565 21867 24599
rect 21867 24565 21876 24599
rect 21824 24556 21876 24565
rect 22008 24599 22060 24608
rect 22008 24565 22017 24599
rect 22017 24565 22051 24599
rect 22051 24565 22060 24599
rect 22008 24556 22060 24565
rect 22376 24556 22428 24608
rect 23848 24556 23900 24608
rect 5582 24454 5634 24506
rect 5646 24454 5698 24506
rect 5710 24454 5762 24506
rect 5774 24454 5826 24506
rect 5838 24454 5890 24506
rect 14846 24454 14898 24506
rect 14910 24454 14962 24506
rect 14974 24454 15026 24506
rect 15038 24454 15090 24506
rect 15102 24454 15154 24506
rect 24110 24454 24162 24506
rect 24174 24454 24226 24506
rect 24238 24454 24290 24506
rect 24302 24454 24354 24506
rect 24366 24454 24418 24506
rect 13728 24395 13780 24404
rect 13728 24361 13737 24395
rect 13737 24361 13771 24395
rect 13771 24361 13780 24395
rect 13728 24352 13780 24361
rect 15476 24352 15528 24404
rect 15200 24284 15252 24336
rect 13820 24148 13872 24200
rect 14740 24148 14792 24200
rect 15660 24148 15712 24200
rect 16672 24352 16724 24404
rect 18420 24352 18472 24404
rect 18604 24395 18656 24404
rect 18604 24361 18613 24395
rect 18613 24361 18647 24395
rect 18647 24361 18656 24395
rect 18604 24352 18656 24361
rect 20260 24352 20312 24404
rect 18236 24284 18288 24336
rect 20444 24284 20496 24336
rect 16212 24216 16264 24268
rect 19708 24259 19760 24268
rect 12808 24080 12860 24132
rect 14832 24080 14884 24132
rect 17040 24148 17092 24200
rect 15844 24123 15896 24132
rect 15844 24089 15853 24123
rect 15853 24089 15887 24123
rect 15887 24089 15896 24123
rect 15844 24080 15896 24089
rect 16672 24080 16724 24132
rect 17592 24123 17644 24132
rect 17592 24089 17601 24123
rect 17601 24089 17635 24123
rect 17635 24089 17644 24123
rect 17592 24080 17644 24089
rect 17776 24123 17828 24132
rect 17776 24089 17785 24123
rect 17785 24089 17819 24123
rect 17819 24089 17828 24123
rect 17776 24080 17828 24089
rect 19708 24225 19717 24259
rect 19717 24225 19751 24259
rect 19751 24225 19760 24259
rect 19708 24216 19760 24225
rect 21088 24352 21140 24404
rect 25688 24352 25740 24404
rect 25780 24352 25832 24404
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 19248 24148 19300 24200
rect 20260 24148 20312 24200
rect 20352 24148 20404 24200
rect 20904 24191 20956 24200
rect 20904 24157 20913 24191
rect 20913 24157 20947 24191
rect 20947 24157 20956 24191
rect 20904 24148 20956 24157
rect 21272 24191 21324 24200
rect 21272 24157 21281 24191
rect 21281 24157 21315 24191
rect 21315 24157 21324 24191
rect 21272 24148 21324 24157
rect 22008 24191 22060 24200
rect 22008 24157 22017 24191
rect 22017 24157 22051 24191
rect 22051 24157 22060 24191
rect 22008 24148 22060 24157
rect 22192 24191 22244 24200
rect 22192 24157 22201 24191
rect 22201 24157 22235 24191
rect 22235 24157 22244 24191
rect 22652 24191 22704 24200
rect 22192 24148 22244 24157
rect 22652 24157 22661 24191
rect 22661 24157 22695 24191
rect 22695 24157 22704 24191
rect 22652 24148 22704 24157
rect 25228 24216 25280 24268
rect 24860 24148 24912 24200
rect 25412 24216 25464 24268
rect 18420 24123 18472 24132
rect 18420 24089 18429 24123
rect 18429 24089 18463 24123
rect 18463 24089 18472 24123
rect 18420 24080 18472 24089
rect 18972 24080 19024 24132
rect 23296 24080 23348 24132
rect 24768 24080 24820 24132
rect 25136 24080 25188 24132
rect 14556 24012 14608 24064
rect 15476 24055 15528 24064
rect 15476 24021 15485 24055
rect 15485 24021 15519 24055
rect 15519 24021 15528 24055
rect 15476 24012 15528 24021
rect 22376 24012 22428 24064
rect 24492 24012 24544 24064
rect 25780 24055 25832 24064
rect 25780 24021 25789 24055
rect 25789 24021 25823 24055
rect 25823 24021 25832 24055
rect 25780 24012 25832 24021
rect 10214 23910 10266 23962
rect 10278 23910 10330 23962
rect 10342 23910 10394 23962
rect 10406 23910 10458 23962
rect 10470 23910 10522 23962
rect 19478 23910 19530 23962
rect 19542 23910 19594 23962
rect 19606 23910 19658 23962
rect 19670 23910 19722 23962
rect 19734 23910 19786 23962
rect 14648 23715 14700 23724
rect 14648 23681 14657 23715
rect 14657 23681 14691 23715
rect 14691 23681 14700 23715
rect 14648 23672 14700 23681
rect 14832 23715 14884 23724
rect 14832 23681 14841 23715
rect 14841 23681 14875 23715
rect 14875 23681 14884 23715
rect 14832 23672 14884 23681
rect 15568 23715 15620 23724
rect 15568 23681 15577 23715
rect 15577 23681 15611 23715
rect 15611 23681 15620 23715
rect 15568 23672 15620 23681
rect 20352 23808 20404 23860
rect 23296 23851 23348 23860
rect 23296 23817 23305 23851
rect 23305 23817 23339 23851
rect 23339 23817 23348 23851
rect 23296 23808 23348 23817
rect 25228 23808 25280 23860
rect 25964 23808 26016 23860
rect 16488 23740 16540 23792
rect 15752 23715 15804 23724
rect 15752 23681 15761 23715
rect 15761 23681 15795 23715
rect 15795 23681 15804 23715
rect 16672 23715 16724 23724
rect 15752 23672 15804 23681
rect 16672 23681 16681 23715
rect 16681 23681 16715 23715
rect 16715 23681 16724 23715
rect 16672 23672 16724 23681
rect 19340 23740 19392 23792
rect 20444 23740 20496 23792
rect 20720 23740 20772 23792
rect 22008 23740 22060 23792
rect 18144 23715 18196 23724
rect 18144 23681 18153 23715
rect 18153 23681 18187 23715
rect 18187 23681 18196 23715
rect 18144 23672 18196 23681
rect 18420 23715 18472 23724
rect 18420 23681 18454 23715
rect 18454 23681 18472 23715
rect 18420 23672 18472 23681
rect 19984 23672 20036 23724
rect 20536 23715 20588 23724
rect 15476 23604 15528 23656
rect 20536 23681 20545 23715
rect 20545 23681 20579 23715
rect 20579 23681 20588 23715
rect 20536 23672 20588 23681
rect 22192 23672 22244 23724
rect 24492 23740 24544 23792
rect 24768 23740 24820 23792
rect 24860 23783 24912 23792
rect 24860 23749 24869 23783
rect 24869 23749 24903 23783
rect 24903 23749 24912 23783
rect 24860 23740 24912 23749
rect 26148 23740 26200 23792
rect 23848 23715 23900 23724
rect 14464 23536 14516 23588
rect 21732 23604 21784 23656
rect 22100 23647 22152 23656
rect 22100 23613 22109 23647
rect 22109 23613 22143 23647
rect 22143 23613 22152 23647
rect 22100 23604 22152 23613
rect 23848 23681 23857 23715
rect 23857 23681 23891 23715
rect 23891 23681 23900 23715
rect 23848 23672 23900 23681
rect 25044 23672 25096 23724
rect 25504 23715 25556 23724
rect 25504 23681 25538 23715
rect 25538 23681 25556 23715
rect 25504 23672 25556 23681
rect 28264 23715 28316 23724
rect 28264 23681 28273 23715
rect 28273 23681 28307 23715
rect 28307 23681 28316 23715
rect 28264 23672 28316 23681
rect 23756 23604 23808 23656
rect 23940 23647 23992 23656
rect 23940 23613 23949 23647
rect 23949 23613 23983 23647
rect 23983 23613 23992 23647
rect 23940 23604 23992 23613
rect 24584 23604 24636 23656
rect 25228 23647 25280 23656
rect 25228 23613 25237 23647
rect 25237 23613 25271 23647
rect 25271 23613 25280 23647
rect 25228 23604 25280 23613
rect 20260 23536 20312 23588
rect 20352 23536 20404 23588
rect 20812 23536 20864 23588
rect 25136 23536 25188 23588
rect 27988 23536 28040 23588
rect 1400 23511 1452 23520
rect 1400 23477 1409 23511
rect 1409 23477 1443 23511
rect 1443 23477 1452 23511
rect 1400 23468 1452 23477
rect 14740 23468 14792 23520
rect 15936 23468 15988 23520
rect 16856 23468 16908 23520
rect 20076 23468 20128 23520
rect 21916 23468 21968 23520
rect 5582 23366 5634 23418
rect 5646 23366 5698 23418
rect 5710 23366 5762 23418
rect 5774 23366 5826 23418
rect 5838 23366 5890 23418
rect 14846 23366 14898 23418
rect 14910 23366 14962 23418
rect 14974 23366 15026 23418
rect 15038 23366 15090 23418
rect 15102 23366 15154 23418
rect 24110 23366 24162 23418
rect 24174 23366 24226 23418
rect 24238 23366 24290 23418
rect 24302 23366 24354 23418
rect 24366 23366 24418 23418
rect 13820 23264 13872 23316
rect 14648 23264 14700 23316
rect 15568 23264 15620 23316
rect 14464 23128 14516 23180
rect 18144 23264 18196 23316
rect 18512 23264 18564 23316
rect 18788 23307 18840 23316
rect 18788 23273 18797 23307
rect 18797 23273 18831 23307
rect 18831 23273 18840 23307
rect 18788 23264 18840 23273
rect 20536 23264 20588 23316
rect 22468 23264 22520 23316
rect 22652 23264 22704 23316
rect 25228 23264 25280 23316
rect 25504 23264 25556 23316
rect 16672 23196 16724 23248
rect 14556 23060 14608 23112
rect 13360 22992 13412 23044
rect 15752 23060 15804 23112
rect 15936 23103 15988 23112
rect 15936 23069 15970 23103
rect 15970 23069 15988 23103
rect 15936 23060 15988 23069
rect 19984 23196 20036 23248
rect 23388 23239 23440 23248
rect 23388 23205 23397 23239
rect 23397 23205 23431 23239
rect 23431 23205 23440 23239
rect 23388 23196 23440 23205
rect 18512 23128 18564 23180
rect 21824 23128 21876 23180
rect 23480 23128 23532 23180
rect 18972 23060 19024 23112
rect 20444 23060 20496 23112
rect 21272 23060 21324 23112
rect 20536 23035 20588 23044
rect 20536 23001 20545 23035
rect 20545 23001 20579 23035
rect 20579 23001 20588 23035
rect 20536 22992 20588 23001
rect 21916 23035 21968 23044
rect 21916 23001 21925 23035
rect 21925 23001 21959 23035
rect 21959 23001 21968 23035
rect 21916 22992 21968 23001
rect 22100 23060 22152 23112
rect 22468 23060 22520 23112
rect 25044 23196 25096 23248
rect 25780 23128 25832 23180
rect 23756 23060 23808 23112
rect 23940 23060 23992 23112
rect 25504 23060 25556 23112
rect 25964 23103 26016 23112
rect 22928 22992 22980 23044
rect 24492 23035 24544 23044
rect 24492 23001 24501 23035
rect 24501 23001 24535 23035
rect 24535 23001 24544 23035
rect 24492 22992 24544 23001
rect 25964 23069 25973 23103
rect 25973 23069 26007 23103
rect 26007 23069 26016 23103
rect 25964 23060 26016 23069
rect 26148 23060 26200 23112
rect 18604 22924 18656 22976
rect 19892 22967 19944 22976
rect 19892 22933 19901 22967
rect 19901 22933 19935 22967
rect 19935 22933 19944 22967
rect 19892 22924 19944 22933
rect 23480 22924 23532 22976
rect 23664 22924 23716 22976
rect 24952 22924 25004 22976
rect 10214 22822 10266 22874
rect 10278 22822 10330 22874
rect 10342 22822 10394 22874
rect 10406 22822 10458 22874
rect 10470 22822 10522 22874
rect 19478 22822 19530 22874
rect 19542 22822 19594 22874
rect 19606 22822 19658 22874
rect 19670 22822 19722 22874
rect 19734 22822 19786 22874
rect 16212 22763 16264 22772
rect 16212 22729 16221 22763
rect 16221 22729 16255 22763
rect 16255 22729 16264 22763
rect 16212 22720 16264 22729
rect 18604 22720 18656 22772
rect 19892 22720 19944 22772
rect 23756 22763 23808 22772
rect 23756 22729 23765 22763
rect 23765 22729 23799 22763
rect 23799 22729 23808 22763
rect 23756 22720 23808 22729
rect 13820 22652 13872 22704
rect 14740 22652 14792 22704
rect 17776 22584 17828 22636
rect 20168 22584 20220 22636
rect 20812 22627 20864 22636
rect 20812 22593 20821 22627
rect 20821 22593 20855 22627
rect 20855 22593 20864 22627
rect 20812 22584 20864 22593
rect 21824 22584 21876 22636
rect 22652 22652 22704 22704
rect 23388 22584 23440 22636
rect 19340 22559 19392 22568
rect 19340 22525 19349 22559
rect 19349 22525 19383 22559
rect 19383 22525 19392 22559
rect 19340 22516 19392 22525
rect 22928 22516 22980 22568
rect 23940 22652 23992 22704
rect 24584 22720 24636 22772
rect 25044 22720 25096 22772
rect 25320 22652 25372 22704
rect 24216 22584 24268 22636
rect 25596 22627 25648 22636
rect 19892 22448 19944 22500
rect 23572 22448 23624 22500
rect 23848 22448 23900 22500
rect 11980 22380 12032 22432
rect 12532 22380 12584 22432
rect 24584 22448 24636 22500
rect 24768 22448 24820 22500
rect 25596 22593 25605 22627
rect 25605 22593 25639 22627
rect 25639 22593 25648 22627
rect 25596 22584 25648 22593
rect 27252 22627 27304 22636
rect 27252 22593 27286 22627
rect 27286 22593 27304 22627
rect 27252 22584 27304 22593
rect 25228 22516 25280 22568
rect 26056 22448 26108 22500
rect 25412 22380 25464 22432
rect 25504 22423 25556 22432
rect 25504 22389 25513 22423
rect 25513 22389 25547 22423
rect 25547 22389 25556 22423
rect 25504 22380 25556 22389
rect 25872 22380 25924 22432
rect 5582 22278 5634 22330
rect 5646 22278 5698 22330
rect 5710 22278 5762 22330
rect 5774 22278 5826 22330
rect 5838 22278 5890 22330
rect 14846 22278 14898 22330
rect 14910 22278 14962 22330
rect 14974 22278 15026 22330
rect 15038 22278 15090 22330
rect 15102 22278 15154 22330
rect 24110 22278 24162 22330
rect 24174 22278 24226 22330
rect 24238 22278 24290 22330
rect 24302 22278 24354 22330
rect 24366 22278 24418 22330
rect 19064 22108 19116 22160
rect 19984 22108 20036 22160
rect 4436 22040 4488 22092
rect 14188 22040 14240 22092
rect 16396 22040 16448 22092
rect 17408 22040 17460 22092
rect 17776 22083 17828 22092
rect 17776 22049 17785 22083
rect 17785 22049 17819 22083
rect 17819 22049 17828 22083
rect 17776 22040 17828 22049
rect 18052 22083 18104 22092
rect 18052 22049 18061 22083
rect 18061 22049 18095 22083
rect 18095 22049 18104 22083
rect 18052 22040 18104 22049
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 13360 21972 13412 22024
rect 14280 22015 14332 22024
rect 11980 21947 12032 21956
rect 11980 21913 11989 21947
rect 11989 21913 12023 21947
rect 12023 21913 12032 21947
rect 11980 21904 12032 21913
rect 12716 21947 12768 21956
rect 12716 21913 12725 21947
rect 12725 21913 12759 21947
rect 12759 21913 12768 21947
rect 12716 21904 12768 21913
rect 13544 21904 13596 21956
rect 12624 21836 12676 21888
rect 14280 21981 14289 22015
rect 14289 21981 14323 22015
rect 14323 21981 14332 22015
rect 14280 21972 14332 21981
rect 15752 21972 15804 22024
rect 16212 21972 16264 22024
rect 17592 21972 17644 22024
rect 18880 21972 18932 22024
rect 23480 22176 23532 22228
rect 24768 22176 24820 22228
rect 27252 22219 27304 22228
rect 27252 22185 27261 22219
rect 27261 22185 27295 22219
rect 27295 22185 27304 22219
rect 27252 22176 27304 22185
rect 20444 22015 20496 22024
rect 14372 21836 14424 21888
rect 15660 21879 15712 21888
rect 15660 21845 15669 21879
rect 15669 21845 15703 21879
rect 15703 21845 15712 21879
rect 15660 21836 15712 21845
rect 16488 21836 16540 21888
rect 19340 21836 19392 21888
rect 19892 21836 19944 21888
rect 20444 21981 20453 22015
rect 20453 21981 20487 22015
rect 20487 21981 20496 22015
rect 20444 21972 20496 21981
rect 23572 22015 23624 22024
rect 23572 21981 23581 22015
rect 23581 21981 23615 22015
rect 23615 21981 23624 22015
rect 23572 21972 23624 21981
rect 23664 22015 23716 22024
rect 23664 21981 23673 22015
rect 23673 21981 23707 22015
rect 23707 21981 23716 22015
rect 23664 21972 23716 21981
rect 23848 21972 23900 22024
rect 24308 22040 24360 22092
rect 24584 22108 24636 22160
rect 28356 22151 28408 22160
rect 28356 22117 28365 22151
rect 28365 22117 28399 22151
rect 28399 22117 28408 22151
rect 28356 22108 28408 22117
rect 24952 22040 25004 22092
rect 26056 22083 26108 22092
rect 20720 21947 20772 21956
rect 20720 21913 20754 21947
rect 20754 21913 20772 21947
rect 20720 21904 20772 21913
rect 24308 21904 24360 21956
rect 24860 21972 24912 22024
rect 25504 21947 25556 21956
rect 25504 21913 25513 21947
rect 25513 21913 25547 21947
rect 25547 21913 25556 21947
rect 25504 21904 25556 21913
rect 26056 22049 26065 22083
rect 26065 22049 26099 22083
rect 26099 22049 26108 22083
rect 26056 22040 26108 22049
rect 25964 21972 26016 22024
rect 27068 22015 27120 22024
rect 27068 21981 27077 22015
rect 27077 21981 27111 22015
rect 27111 21981 27120 22015
rect 27068 21972 27120 21981
rect 21732 21836 21784 21888
rect 23480 21836 23532 21888
rect 24676 21836 24728 21888
rect 25964 21836 26016 21888
rect 26516 21836 26568 21888
rect 10214 21734 10266 21786
rect 10278 21734 10330 21786
rect 10342 21734 10394 21786
rect 10406 21734 10458 21786
rect 10470 21734 10522 21786
rect 19478 21734 19530 21786
rect 19542 21734 19594 21786
rect 19606 21734 19658 21786
rect 19670 21734 19722 21786
rect 19734 21734 19786 21786
rect 12716 21632 12768 21684
rect 14004 21675 14056 21684
rect 14004 21641 14013 21675
rect 14013 21641 14047 21675
rect 14047 21641 14056 21675
rect 14004 21632 14056 21641
rect 11520 21428 11572 21480
rect 13820 21564 13872 21616
rect 12348 21496 12400 21548
rect 14004 21496 14056 21548
rect 14372 21539 14424 21548
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 15660 21564 15712 21616
rect 17960 21496 18012 21548
rect 18052 21496 18104 21548
rect 19892 21632 19944 21684
rect 21180 21632 21232 21684
rect 23480 21632 23532 21684
rect 18696 21539 18748 21548
rect 18696 21505 18705 21539
rect 18705 21505 18739 21539
rect 18739 21505 18748 21539
rect 19064 21539 19116 21548
rect 18696 21496 18748 21505
rect 19064 21505 19073 21539
rect 19073 21505 19107 21539
rect 19107 21505 19116 21539
rect 19064 21496 19116 21505
rect 19156 21496 19208 21548
rect 20168 21564 20220 21616
rect 20260 21564 20312 21616
rect 17224 21360 17276 21412
rect 18880 21428 18932 21480
rect 19524 21428 19576 21480
rect 20076 21496 20128 21548
rect 20352 21539 20404 21548
rect 20352 21505 20361 21539
rect 20361 21505 20395 21539
rect 20395 21505 20404 21539
rect 20352 21496 20404 21505
rect 20812 21564 20864 21616
rect 24768 21632 24820 21684
rect 21916 21496 21968 21548
rect 22100 21539 22152 21548
rect 22100 21505 22134 21539
rect 22134 21505 22152 21539
rect 25412 21607 25464 21616
rect 22100 21496 22152 21505
rect 20444 21428 20496 21480
rect 15568 21292 15620 21344
rect 16488 21292 16540 21344
rect 17592 21335 17644 21344
rect 17592 21301 17601 21335
rect 17601 21301 17635 21335
rect 17635 21301 17644 21335
rect 17592 21292 17644 21301
rect 19892 21360 19944 21412
rect 20628 21360 20680 21412
rect 20720 21360 20772 21412
rect 21180 21292 21232 21344
rect 22192 21292 22244 21344
rect 23940 21496 23992 21548
rect 24768 21496 24820 21548
rect 25412 21573 25421 21607
rect 25421 21573 25455 21607
rect 25455 21573 25464 21607
rect 25412 21564 25464 21573
rect 25504 21564 25556 21616
rect 25044 21496 25096 21548
rect 26148 21496 26200 21548
rect 26424 21539 26476 21548
rect 26424 21505 26433 21539
rect 26433 21505 26467 21539
rect 26467 21505 26476 21539
rect 26424 21496 26476 21505
rect 23664 21403 23716 21412
rect 23664 21369 23673 21403
rect 23673 21369 23707 21403
rect 23707 21369 23716 21403
rect 23664 21360 23716 21369
rect 23848 21360 23900 21412
rect 23572 21292 23624 21344
rect 23940 21292 23992 21344
rect 24676 21335 24728 21344
rect 24676 21301 24685 21335
rect 24685 21301 24719 21335
rect 24719 21301 24728 21335
rect 24676 21292 24728 21301
rect 25872 21292 25924 21344
rect 26056 21292 26108 21344
rect 26332 21335 26384 21344
rect 26332 21301 26341 21335
rect 26341 21301 26375 21335
rect 26375 21301 26384 21335
rect 26332 21292 26384 21301
rect 28356 21335 28408 21344
rect 28356 21301 28365 21335
rect 28365 21301 28399 21335
rect 28399 21301 28408 21335
rect 28356 21292 28408 21301
rect 5582 21190 5634 21242
rect 5646 21190 5698 21242
rect 5710 21190 5762 21242
rect 5774 21190 5826 21242
rect 5838 21190 5890 21242
rect 14846 21190 14898 21242
rect 14910 21190 14962 21242
rect 14974 21190 15026 21242
rect 15038 21190 15090 21242
rect 15102 21190 15154 21242
rect 24110 21190 24162 21242
rect 24174 21190 24226 21242
rect 24238 21190 24290 21242
rect 24302 21190 24354 21242
rect 24366 21190 24418 21242
rect 12348 21088 12400 21140
rect 15752 21131 15804 21140
rect 13176 21020 13228 21072
rect 13820 21020 13872 21072
rect 15752 21097 15761 21131
rect 15761 21097 15795 21131
rect 15795 21097 15804 21131
rect 15752 21088 15804 21097
rect 12256 20816 12308 20868
rect 12624 20927 12676 20936
rect 12624 20893 12633 20927
rect 12633 20893 12667 20927
rect 12667 20893 12676 20927
rect 12624 20884 12676 20893
rect 12900 20884 12952 20936
rect 13360 20927 13412 20936
rect 13360 20893 13369 20927
rect 13369 20893 13403 20927
rect 13403 20893 13412 20927
rect 13360 20884 13412 20893
rect 14188 20884 14240 20936
rect 17224 21020 17276 21072
rect 20352 21088 20404 21140
rect 22100 21088 22152 21140
rect 23848 21088 23900 21140
rect 24676 21131 24728 21140
rect 19524 21020 19576 21072
rect 20076 21020 20128 21072
rect 20996 21020 21048 21072
rect 21824 21020 21876 21072
rect 24400 21020 24452 21072
rect 24676 21097 24685 21131
rect 24685 21097 24719 21131
rect 24719 21097 24728 21131
rect 24676 21088 24728 21097
rect 24860 21020 24912 21072
rect 14740 20927 14792 20936
rect 14740 20893 14749 20927
rect 14749 20893 14783 20927
rect 14783 20893 14792 20927
rect 20260 20952 20312 21004
rect 15936 20927 15988 20936
rect 14740 20884 14792 20893
rect 15936 20893 15945 20927
rect 15945 20893 15979 20927
rect 15979 20893 15988 20927
rect 15936 20884 15988 20893
rect 16396 20927 16448 20936
rect 15200 20859 15252 20868
rect 15200 20825 15209 20859
rect 15209 20825 15243 20859
rect 15243 20825 15252 20859
rect 15200 20816 15252 20825
rect 15292 20816 15344 20868
rect 16396 20893 16405 20927
rect 16405 20893 16439 20927
rect 16439 20893 16448 20927
rect 16396 20884 16448 20893
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 17592 20884 17644 20936
rect 19524 20927 19576 20936
rect 19524 20893 19533 20927
rect 19533 20893 19567 20927
rect 19567 20893 19576 20927
rect 19524 20884 19576 20893
rect 20628 20927 20680 20936
rect 20628 20893 20637 20927
rect 20637 20893 20671 20927
rect 20671 20893 20680 20927
rect 20628 20884 20680 20893
rect 21364 20952 21416 21004
rect 20812 20927 20864 20936
rect 20812 20893 20821 20927
rect 20821 20893 20855 20927
rect 20855 20893 20864 20927
rect 20812 20884 20864 20893
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 20996 20884 21048 20893
rect 21824 20927 21876 20936
rect 21824 20893 21833 20927
rect 21833 20893 21867 20927
rect 21867 20893 21876 20927
rect 21824 20884 21876 20893
rect 23112 20952 23164 21004
rect 22192 20884 22244 20936
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 22560 20884 22612 20893
rect 23664 20884 23716 20936
rect 23848 20927 23900 20936
rect 23848 20893 23857 20927
rect 23857 20893 23891 20927
rect 23891 20893 23900 20927
rect 23848 20884 23900 20893
rect 24676 20952 24728 21004
rect 24768 20927 24820 20936
rect 24768 20893 24777 20927
rect 24777 20893 24811 20927
rect 24811 20893 24820 20927
rect 24768 20884 24820 20893
rect 24952 20884 25004 20936
rect 18328 20816 18380 20868
rect 14096 20791 14148 20800
rect 14096 20757 14105 20791
rect 14105 20757 14139 20791
rect 14139 20757 14148 20791
rect 14096 20748 14148 20757
rect 16856 20791 16908 20800
rect 16856 20757 16865 20791
rect 16865 20757 16899 20791
rect 16899 20757 16908 20791
rect 16856 20748 16908 20757
rect 17132 20748 17184 20800
rect 18696 20748 18748 20800
rect 20444 20816 20496 20868
rect 23204 20859 23256 20868
rect 23204 20825 23213 20859
rect 23213 20825 23247 20859
rect 23247 20825 23256 20859
rect 23204 20816 23256 20825
rect 23296 20816 23348 20868
rect 25688 20995 25740 21004
rect 25688 20961 25697 20995
rect 25697 20961 25731 20995
rect 25731 20961 25740 20995
rect 25688 20952 25740 20961
rect 26332 21020 26384 21072
rect 25320 20927 25372 20936
rect 25320 20893 25329 20927
rect 25329 20893 25363 20927
rect 25363 20893 25372 20927
rect 25872 20927 25924 20936
rect 25320 20884 25372 20893
rect 25872 20893 25881 20927
rect 25881 20893 25915 20927
rect 25915 20893 25924 20927
rect 25872 20884 25924 20893
rect 26056 20884 26108 20936
rect 26608 20884 26660 20936
rect 26884 20884 26936 20936
rect 20076 20791 20128 20800
rect 20076 20757 20085 20791
rect 20085 20757 20119 20791
rect 20119 20757 20128 20791
rect 20076 20748 20128 20757
rect 20352 20791 20404 20800
rect 20352 20757 20361 20791
rect 20361 20757 20395 20791
rect 20395 20757 20404 20791
rect 20352 20748 20404 20757
rect 25228 20748 25280 20800
rect 10214 20646 10266 20698
rect 10278 20646 10330 20698
rect 10342 20646 10394 20698
rect 10406 20646 10458 20698
rect 10470 20646 10522 20698
rect 19478 20646 19530 20698
rect 19542 20646 19594 20698
rect 19606 20646 19658 20698
rect 19670 20646 19722 20698
rect 19734 20646 19786 20698
rect 13084 20544 13136 20596
rect 15292 20544 15344 20596
rect 15936 20544 15988 20596
rect 17960 20544 18012 20596
rect 20628 20544 20680 20596
rect 23664 20544 23716 20596
rect 25872 20544 25924 20596
rect 26516 20587 26568 20596
rect 26516 20553 26525 20587
rect 26525 20553 26559 20587
rect 26559 20553 26568 20587
rect 26516 20544 26568 20553
rect 13544 20519 13596 20528
rect 13544 20485 13553 20519
rect 13553 20485 13587 20519
rect 13587 20485 13596 20519
rect 13544 20476 13596 20485
rect 14096 20519 14148 20528
rect 14096 20485 14130 20519
rect 14130 20485 14148 20519
rect 14096 20476 14148 20485
rect 9680 20408 9732 20460
rect 11796 20451 11848 20460
rect 11796 20417 11830 20451
rect 11830 20417 11848 20451
rect 13820 20451 13872 20460
rect 11796 20408 11848 20417
rect 13820 20417 13829 20451
rect 13829 20417 13863 20451
rect 13863 20417 13872 20451
rect 13820 20408 13872 20417
rect 16396 20408 16448 20460
rect 16948 20408 17000 20460
rect 18696 20476 18748 20528
rect 19340 20476 19392 20528
rect 20536 20476 20588 20528
rect 8852 20340 8904 20392
rect 11520 20383 11572 20392
rect 11520 20349 11529 20383
rect 11529 20349 11563 20383
rect 11563 20349 11572 20383
rect 11520 20340 11572 20349
rect 16488 20340 16540 20392
rect 16212 20272 16264 20324
rect 17224 20340 17276 20392
rect 18328 20451 18380 20460
rect 18328 20417 18337 20451
rect 18337 20417 18371 20451
rect 18371 20417 18380 20451
rect 18328 20408 18380 20417
rect 19064 20408 19116 20460
rect 20168 20408 20220 20460
rect 20352 20451 20404 20460
rect 20352 20417 20386 20451
rect 20386 20417 20404 20451
rect 20352 20408 20404 20417
rect 23112 20451 23164 20460
rect 23112 20417 23121 20451
rect 23121 20417 23155 20451
rect 23155 20417 23164 20451
rect 23112 20408 23164 20417
rect 25504 20476 25556 20528
rect 25688 20476 25740 20528
rect 23480 20408 23532 20460
rect 23848 20408 23900 20460
rect 25320 20451 25372 20460
rect 25320 20417 25329 20451
rect 25329 20417 25363 20451
rect 25363 20417 25372 20451
rect 25320 20408 25372 20417
rect 25596 20451 25648 20460
rect 25596 20417 25605 20451
rect 25605 20417 25639 20451
rect 25639 20417 25648 20451
rect 25596 20408 25648 20417
rect 26792 20408 26844 20460
rect 19248 20272 19300 20324
rect 21088 20340 21140 20392
rect 23204 20340 23256 20392
rect 24768 20340 24820 20392
rect 21916 20272 21968 20324
rect 24584 20272 24636 20324
rect 25504 20340 25556 20392
rect 26056 20340 26108 20392
rect 26884 20340 26936 20392
rect 8392 20204 8444 20256
rect 12624 20204 12676 20256
rect 15200 20247 15252 20256
rect 15200 20213 15209 20247
rect 15209 20213 15243 20247
rect 15243 20213 15252 20247
rect 15200 20204 15252 20213
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 18420 20204 18472 20256
rect 18788 20204 18840 20256
rect 19156 20247 19208 20256
rect 19156 20213 19165 20247
rect 19165 20213 19199 20247
rect 19199 20213 19208 20247
rect 19156 20204 19208 20213
rect 24032 20204 24084 20256
rect 26424 20272 26476 20324
rect 26332 20247 26384 20256
rect 26332 20213 26341 20247
rect 26341 20213 26375 20247
rect 26375 20213 26384 20247
rect 26332 20204 26384 20213
rect 5582 20102 5634 20154
rect 5646 20102 5698 20154
rect 5710 20102 5762 20154
rect 5774 20102 5826 20154
rect 5838 20102 5890 20154
rect 14846 20102 14898 20154
rect 14910 20102 14962 20154
rect 14974 20102 15026 20154
rect 15038 20102 15090 20154
rect 15102 20102 15154 20154
rect 24110 20102 24162 20154
rect 24174 20102 24226 20154
rect 24238 20102 24290 20154
rect 24302 20102 24354 20154
rect 24366 20102 24418 20154
rect 11796 20043 11848 20052
rect 11796 20009 11805 20043
rect 11805 20009 11839 20043
rect 11839 20009 11848 20043
rect 11796 20000 11848 20009
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 8944 19839 8996 19848
rect 8944 19805 8953 19839
rect 8953 19805 8987 19839
rect 8987 19805 8996 19839
rect 8944 19796 8996 19805
rect 12072 19839 12124 19848
rect 12072 19805 12095 19839
rect 12095 19805 12124 19839
rect 12072 19796 12124 19805
rect 12256 20000 12308 20052
rect 17132 20000 17184 20052
rect 17776 20043 17828 20052
rect 17776 20009 17785 20043
rect 17785 20009 17819 20043
rect 17819 20009 17828 20043
rect 17776 20000 17828 20009
rect 20168 20000 20220 20052
rect 20352 20000 20404 20052
rect 21088 20043 21140 20052
rect 21088 20009 21097 20043
rect 21097 20009 21131 20043
rect 21131 20009 21140 20043
rect 21088 20000 21140 20009
rect 23296 20000 23348 20052
rect 23848 20000 23900 20052
rect 26792 20043 26844 20052
rect 26792 20009 26801 20043
rect 26801 20009 26835 20043
rect 26835 20009 26844 20043
rect 26792 20000 26844 20009
rect 12624 19864 12676 19916
rect 13084 19907 13136 19916
rect 13084 19873 13093 19907
rect 13093 19873 13127 19907
rect 13127 19873 13136 19907
rect 13084 19864 13136 19873
rect 12716 19839 12768 19848
rect 8852 19660 8904 19712
rect 9864 19660 9916 19712
rect 12072 19660 12124 19712
rect 12716 19805 12725 19839
rect 12725 19805 12759 19839
rect 12759 19805 12768 19839
rect 12716 19796 12768 19805
rect 14280 19932 14332 19984
rect 14924 19932 14976 19984
rect 15108 19932 15160 19984
rect 23664 19932 23716 19984
rect 19248 19907 19300 19916
rect 14740 19796 14792 19848
rect 14924 19839 14976 19848
rect 14924 19805 14933 19839
rect 14933 19805 14967 19839
rect 14967 19805 14976 19839
rect 14924 19796 14976 19805
rect 15108 19796 15160 19848
rect 14556 19728 14608 19780
rect 17500 19796 17552 19848
rect 15660 19728 15712 19780
rect 15844 19771 15896 19780
rect 15844 19737 15853 19771
rect 15853 19737 15887 19771
rect 15887 19737 15896 19771
rect 15844 19728 15896 19737
rect 17040 19728 17092 19780
rect 12900 19660 12952 19712
rect 13728 19660 13780 19712
rect 13820 19660 13872 19712
rect 18420 19839 18472 19848
rect 18420 19805 18429 19839
rect 18429 19805 18463 19839
rect 18463 19805 18472 19839
rect 18420 19796 18472 19805
rect 18604 19796 18656 19848
rect 18972 19796 19024 19848
rect 19248 19873 19257 19907
rect 19257 19873 19291 19907
rect 19291 19873 19300 19907
rect 19248 19864 19300 19873
rect 19892 19796 19944 19848
rect 21456 19839 21508 19848
rect 21456 19805 21465 19839
rect 21465 19805 21499 19839
rect 21499 19805 21508 19839
rect 21456 19796 21508 19805
rect 21548 19839 21600 19848
rect 21548 19805 21557 19839
rect 21557 19805 21591 19839
rect 21591 19805 21600 19839
rect 21548 19796 21600 19805
rect 22376 19839 22428 19848
rect 22376 19805 22385 19839
rect 22385 19805 22419 19839
rect 22419 19805 22428 19839
rect 22376 19796 22428 19805
rect 18696 19660 18748 19712
rect 19156 19660 19208 19712
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 22284 19728 22336 19780
rect 23480 19839 23532 19848
rect 23480 19805 23489 19839
rect 23489 19805 23523 19839
rect 23523 19805 23532 19839
rect 23480 19796 23532 19805
rect 23664 19796 23716 19848
rect 24032 19839 24084 19848
rect 24032 19805 24041 19839
rect 24041 19805 24075 19839
rect 24075 19805 24084 19839
rect 24032 19796 24084 19805
rect 24768 19864 24820 19916
rect 24676 19839 24728 19848
rect 24676 19805 24685 19839
rect 24685 19805 24719 19839
rect 24719 19805 24728 19839
rect 24676 19796 24728 19805
rect 24860 19839 24912 19848
rect 24860 19805 24869 19839
rect 24869 19805 24903 19839
rect 24903 19805 24912 19839
rect 24860 19796 24912 19805
rect 25596 19932 25648 19984
rect 25412 19796 25464 19848
rect 26332 19864 26384 19916
rect 26608 19796 26660 19848
rect 28356 19839 28408 19848
rect 28356 19805 28365 19839
rect 28365 19805 28399 19839
rect 28399 19805 28408 19839
rect 28356 19796 28408 19805
rect 22192 19660 22244 19712
rect 23940 19703 23992 19712
rect 23940 19669 23949 19703
rect 23949 19669 23983 19703
rect 23983 19669 23992 19703
rect 26424 19728 26476 19780
rect 23940 19660 23992 19669
rect 25412 19703 25464 19712
rect 25412 19669 25421 19703
rect 25421 19669 25455 19703
rect 25455 19669 25464 19703
rect 25412 19660 25464 19669
rect 25504 19660 25556 19712
rect 25872 19703 25924 19712
rect 25872 19669 25881 19703
rect 25881 19669 25915 19703
rect 25915 19669 25924 19703
rect 25872 19660 25924 19669
rect 26240 19660 26292 19712
rect 10214 19558 10266 19610
rect 10278 19558 10330 19610
rect 10342 19558 10394 19610
rect 10406 19558 10458 19610
rect 10470 19558 10522 19610
rect 19478 19558 19530 19610
rect 19542 19558 19594 19610
rect 19606 19558 19658 19610
rect 19670 19558 19722 19610
rect 19734 19558 19786 19610
rect 9680 19499 9732 19508
rect 9680 19465 9689 19499
rect 9689 19465 9723 19499
rect 9723 19465 9732 19499
rect 9680 19456 9732 19465
rect 13820 19456 13872 19508
rect 14924 19456 14976 19508
rect 15292 19456 15344 19508
rect 15384 19456 15436 19508
rect 17500 19456 17552 19508
rect 19248 19456 19300 19508
rect 20812 19456 20864 19508
rect 23940 19456 23992 19508
rect 25044 19456 25096 19508
rect 25504 19456 25556 19508
rect 26240 19456 26292 19508
rect 11980 19388 12032 19440
rect 8484 19363 8536 19372
rect 8484 19329 8493 19363
rect 8493 19329 8527 19363
rect 8527 19329 8536 19363
rect 8484 19320 8536 19329
rect 9036 19363 9088 19372
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 9864 19320 9916 19372
rect 11336 19320 11388 19372
rect 8852 19295 8904 19304
rect 8852 19261 8861 19295
rect 8861 19261 8895 19295
rect 8895 19261 8904 19295
rect 8852 19252 8904 19261
rect 10324 19295 10376 19304
rect 10324 19261 10333 19295
rect 10333 19261 10367 19295
rect 10367 19261 10376 19295
rect 10324 19252 10376 19261
rect 11888 19320 11940 19372
rect 14464 19388 14516 19440
rect 13636 19320 13688 19372
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 14924 19320 14976 19372
rect 17224 19388 17276 19440
rect 19340 19388 19392 19440
rect 20168 19431 20220 19440
rect 20168 19397 20177 19431
rect 20177 19397 20211 19431
rect 20211 19397 20220 19431
rect 20168 19388 20220 19397
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 17316 19363 17368 19372
rect 17316 19329 17325 19363
rect 17325 19329 17359 19363
rect 17359 19329 17368 19363
rect 17316 19320 17368 19329
rect 17868 19320 17920 19372
rect 18604 19320 18656 19372
rect 18788 19363 18840 19372
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 18788 19320 18840 19329
rect 19156 19320 19208 19372
rect 19524 19363 19576 19372
rect 19524 19329 19533 19363
rect 19533 19329 19567 19363
rect 19567 19329 19576 19363
rect 19524 19320 19576 19329
rect 8300 19227 8352 19236
rect 8300 19193 8309 19227
rect 8309 19193 8343 19227
rect 8343 19193 8352 19227
rect 8300 19184 8352 19193
rect 14740 19184 14792 19236
rect 15752 19252 15804 19304
rect 18328 19252 18380 19304
rect 19984 19295 20036 19304
rect 16304 19184 16356 19236
rect 19984 19261 19993 19295
rect 19993 19261 20027 19295
rect 20027 19261 20036 19295
rect 19984 19252 20036 19261
rect 18972 19227 19024 19236
rect 18972 19193 18981 19227
rect 18981 19193 19015 19227
rect 19015 19193 19024 19227
rect 18972 19184 19024 19193
rect 20720 19320 20772 19372
rect 21456 19363 21508 19372
rect 21456 19329 21465 19363
rect 21465 19329 21499 19363
rect 21499 19329 21508 19363
rect 21824 19363 21876 19372
rect 21456 19320 21508 19329
rect 21824 19329 21833 19363
rect 21833 19329 21867 19363
rect 21867 19329 21876 19363
rect 21824 19320 21876 19329
rect 22284 19320 22336 19372
rect 23664 19320 23716 19372
rect 23940 19363 23992 19372
rect 23940 19329 23949 19363
rect 23949 19329 23983 19363
rect 23983 19329 23992 19363
rect 23940 19320 23992 19329
rect 24492 19388 24544 19440
rect 25136 19388 25188 19440
rect 27068 19456 27120 19508
rect 26332 19320 26384 19372
rect 26516 19320 26568 19372
rect 24492 19252 24544 19304
rect 25964 19252 26016 19304
rect 22652 19184 22704 19236
rect 26884 19184 26936 19236
rect 9496 19116 9548 19168
rect 11980 19116 12032 19168
rect 12624 19116 12676 19168
rect 12900 19116 12952 19168
rect 17592 19116 17644 19168
rect 17684 19116 17736 19168
rect 20628 19116 20680 19168
rect 23756 19159 23808 19168
rect 23756 19125 23765 19159
rect 23765 19125 23799 19159
rect 23799 19125 23808 19159
rect 23756 19116 23808 19125
rect 24584 19116 24636 19168
rect 26240 19159 26292 19168
rect 26240 19125 26249 19159
rect 26249 19125 26283 19159
rect 26283 19125 26292 19159
rect 26240 19116 26292 19125
rect 28172 19116 28224 19168
rect 5582 19014 5634 19066
rect 5646 19014 5698 19066
rect 5710 19014 5762 19066
rect 5774 19014 5826 19066
rect 5838 19014 5890 19066
rect 14846 19014 14898 19066
rect 14910 19014 14962 19066
rect 14974 19014 15026 19066
rect 15038 19014 15090 19066
rect 15102 19014 15154 19066
rect 24110 19014 24162 19066
rect 24174 19014 24226 19066
rect 24238 19014 24290 19066
rect 24302 19014 24354 19066
rect 24366 19014 24418 19066
rect 9036 18912 9088 18964
rect 11888 18955 11940 18964
rect 11888 18921 11897 18955
rect 11897 18921 11931 18955
rect 11931 18921 11940 18955
rect 11888 18912 11940 18921
rect 13636 18912 13688 18964
rect 14556 18955 14608 18964
rect 9036 18776 9088 18828
rect 10324 18776 10376 18828
rect 11520 18776 11572 18828
rect 14556 18921 14565 18955
rect 14565 18921 14599 18955
rect 14599 18921 14608 18955
rect 14556 18912 14608 18921
rect 15752 18955 15804 18964
rect 15752 18921 15761 18955
rect 15761 18921 15795 18955
rect 15795 18921 15804 18955
rect 15752 18912 15804 18921
rect 16120 18912 16172 18964
rect 17040 18955 17092 18964
rect 17040 18921 17049 18955
rect 17049 18921 17083 18955
rect 17083 18921 17092 18955
rect 17040 18912 17092 18921
rect 19340 18912 19392 18964
rect 19524 18912 19576 18964
rect 20536 18912 20588 18964
rect 22284 18912 22336 18964
rect 22560 18912 22612 18964
rect 24032 18955 24084 18964
rect 24032 18921 24041 18955
rect 24041 18921 24075 18955
rect 24075 18921 24084 18955
rect 24032 18912 24084 18921
rect 24492 18912 24544 18964
rect 25964 18955 26016 18964
rect 25964 18921 25973 18955
rect 25973 18921 26007 18955
rect 26007 18921 26016 18955
rect 25964 18912 26016 18921
rect 26240 18955 26292 18964
rect 26240 18921 26249 18955
rect 26249 18921 26283 18955
rect 26283 18921 26292 18955
rect 26240 18912 26292 18921
rect 27804 18955 27856 18964
rect 27804 18921 27813 18955
rect 27813 18921 27847 18955
rect 27847 18921 27856 18955
rect 27804 18912 27856 18921
rect 28172 18955 28224 18964
rect 28172 18921 28181 18955
rect 28181 18921 28215 18955
rect 28215 18921 28224 18955
rect 28172 18912 28224 18921
rect 13820 18844 13872 18896
rect 14004 18844 14056 18896
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 8300 18708 8352 18760
rect 9864 18708 9916 18760
rect 15200 18776 15252 18828
rect 16212 18776 16264 18828
rect 16580 18819 16632 18828
rect 16580 18785 16589 18819
rect 16589 18785 16623 18819
rect 16623 18785 16632 18819
rect 16580 18776 16632 18785
rect 6644 18640 6696 18692
rect 8944 18640 8996 18692
rect 9404 18640 9456 18692
rect 11520 18640 11572 18692
rect 13084 18640 13136 18692
rect 14188 18683 14240 18692
rect 14188 18649 14197 18683
rect 14197 18649 14231 18683
rect 14231 18649 14240 18683
rect 14188 18640 14240 18649
rect 14280 18640 14332 18692
rect 14740 18640 14792 18692
rect 16120 18708 16172 18760
rect 15936 18640 15988 18692
rect 16304 18640 16356 18692
rect 19984 18844 20036 18896
rect 17500 18819 17552 18828
rect 17500 18785 17509 18819
rect 17509 18785 17543 18819
rect 17543 18785 17552 18819
rect 17500 18776 17552 18785
rect 20168 18776 20220 18828
rect 17224 18751 17276 18760
rect 17224 18717 17233 18751
rect 17233 18717 17267 18751
rect 17267 18717 17276 18751
rect 17224 18708 17276 18717
rect 17592 18708 17644 18760
rect 19984 18708 20036 18760
rect 20444 18751 20496 18760
rect 20444 18717 20453 18751
rect 20453 18717 20487 18751
rect 20487 18717 20496 18751
rect 20444 18708 20496 18717
rect 20720 18751 20772 18760
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 19248 18640 19300 18692
rect 22468 18844 22520 18896
rect 24676 18844 24728 18896
rect 22100 18776 22152 18828
rect 22652 18819 22704 18828
rect 22652 18785 22661 18819
rect 22661 18785 22695 18819
rect 22695 18785 22704 18819
rect 22652 18776 22704 18785
rect 23756 18708 23808 18760
rect 25504 18776 25556 18828
rect 27068 18844 27120 18896
rect 25044 18751 25096 18760
rect 6920 18615 6972 18624
rect 6920 18581 6929 18615
rect 6929 18581 6963 18615
rect 6963 18581 6972 18615
rect 6920 18572 6972 18581
rect 9956 18572 10008 18624
rect 14372 18572 14424 18624
rect 15200 18615 15252 18624
rect 15200 18581 15209 18615
rect 15209 18581 15243 18615
rect 15243 18581 15252 18615
rect 15200 18572 15252 18581
rect 16396 18615 16448 18624
rect 16396 18581 16405 18615
rect 16405 18581 16439 18615
rect 16439 18581 16448 18615
rect 16396 18572 16448 18581
rect 16672 18572 16724 18624
rect 21364 18572 21416 18624
rect 22376 18572 22428 18624
rect 25044 18717 25053 18751
rect 25053 18717 25087 18751
rect 25087 18717 25096 18751
rect 25044 18708 25096 18717
rect 25872 18708 25924 18760
rect 26332 18708 26384 18760
rect 28080 18751 28132 18760
rect 25136 18640 25188 18692
rect 28080 18717 28089 18751
rect 28089 18717 28123 18751
rect 28123 18717 28132 18751
rect 28080 18708 28132 18717
rect 28264 18708 28316 18760
rect 26424 18572 26476 18624
rect 10214 18470 10266 18522
rect 10278 18470 10330 18522
rect 10342 18470 10394 18522
rect 10406 18470 10458 18522
rect 10470 18470 10522 18522
rect 19478 18470 19530 18522
rect 19542 18470 19594 18522
rect 19606 18470 19658 18522
rect 19670 18470 19722 18522
rect 19734 18470 19786 18522
rect 7380 18368 7432 18420
rect 11520 18411 11572 18420
rect 11520 18377 11529 18411
rect 11529 18377 11563 18411
rect 11563 18377 11572 18411
rect 11520 18368 11572 18377
rect 13084 18411 13136 18420
rect 13084 18377 13093 18411
rect 13093 18377 13127 18411
rect 13127 18377 13136 18411
rect 13084 18368 13136 18377
rect 6920 18343 6972 18352
rect 6920 18309 6954 18343
rect 6954 18309 6972 18343
rect 6920 18300 6972 18309
rect 9496 18275 9548 18284
rect 5172 18164 5224 18216
rect 6644 18207 6696 18216
rect 6644 18173 6653 18207
rect 6653 18173 6687 18207
rect 6687 18173 6696 18207
rect 6644 18164 6696 18173
rect 9036 18164 9088 18216
rect 9496 18241 9505 18275
rect 9505 18241 9539 18275
rect 9539 18241 9548 18275
rect 9496 18232 9548 18241
rect 11520 18232 11572 18284
rect 9404 18164 9456 18216
rect 11704 18232 11756 18284
rect 11980 18275 12032 18284
rect 11980 18241 11994 18275
rect 11994 18241 12028 18275
rect 12028 18241 12032 18275
rect 12164 18275 12216 18284
rect 11980 18232 12032 18241
rect 12164 18241 12173 18275
rect 12173 18241 12207 18275
rect 12207 18241 12216 18275
rect 12164 18232 12216 18241
rect 12624 18275 12676 18284
rect 12624 18241 12633 18275
rect 12633 18241 12667 18275
rect 12667 18241 12676 18275
rect 12624 18232 12676 18241
rect 12348 18164 12400 18216
rect 12992 18232 13044 18284
rect 13820 18300 13872 18352
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 15384 18368 15436 18420
rect 15568 18368 15620 18420
rect 16120 18368 16172 18420
rect 16856 18411 16908 18420
rect 16856 18377 16865 18411
rect 16865 18377 16899 18411
rect 16899 18377 16908 18411
rect 16856 18368 16908 18377
rect 17316 18368 17368 18420
rect 17408 18368 17460 18420
rect 17684 18411 17736 18420
rect 17684 18377 17693 18411
rect 17693 18377 17727 18411
rect 17727 18377 17736 18411
rect 17684 18368 17736 18377
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14740 18275 14792 18284
rect 14556 18232 14608 18241
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 16028 18300 16080 18352
rect 19248 18343 19300 18352
rect 19248 18309 19257 18343
rect 19257 18309 19291 18343
rect 19291 18309 19300 18343
rect 19248 18300 19300 18309
rect 1676 18028 1728 18080
rect 8392 18028 8444 18080
rect 9220 18028 9272 18080
rect 13544 18096 13596 18148
rect 9956 18028 10008 18080
rect 11060 18028 11112 18080
rect 11888 18028 11940 18080
rect 12164 18028 12216 18080
rect 14372 18028 14424 18080
rect 15752 18232 15804 18284
rect 16672 18232 16724 18284
rect 17592 18275 17644 18284
rect 17592 18241 17601 18275
rect 17601 18241 17635 18275
rect 17635 18241 17644 18275
rect 17592 18232 17644 18241
rect 18880 18232 18932 18284
rect 19892 18232 19944 18284
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20168 18232 20220 18241
rect 20444 18275 20496 18284
rect 20444 18241 20453 18275
rect 20453 18241 20487 18275
rect 20487 18241 20496 18275
rect 20444 18232 20496 18241
rect 16948 18164 17000 18216
rect 17868 18207 17920 18216
rect 17868 18173 17877 18207
rect 17877 18173 17911 18207
rect 17911 18173 17920 18207
rect 17868 18164 17920 18173
rect 18512 18164 18564 18216
rect 15384 18096 15436 18148
rect 19064 18096 19116 18148
rect 16764 18028 16816 18080
rect 17132 18028 17184 18080
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 18880 18028 18932 18080
rect 19340 18071 19392 18080
rect 19340 18037 19349 18071
rect 19349 18037 19383 18071
rect 19383 18037 19392 18071
rect 19340 18028 19392 18037
rect 20260 18207 20312 18216
rect 20260 18173 20269 18207
rect 20269 18173 20303 18207
rect 20303 18173 20312 18207
rect 21640 18368 21692 18420
rect 22928 18411 22980 18420
rect 22928 18377 22937 18411
rect 22937 18377 22971 18411
rect 22971 18377 22980 18411
rect 22928 18368 22980 18377
rect 24584 18411 24636 18420
rect 24584 18377 24593 18411
rect 24593 18377 24627 18411
rect 24627 18377 24636 18411
rect 24584 18368 24636 18377
rect 25412 18368 25464 18420
rect 27344 18300 27396 18352
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 22928 18232 22980 18284
rect 24032 18232 24084 18284
rect 25872 18232 25924 18284
rect 26056 18232 26108 18284
rect 26332 18275 26384 18284
rect 26332 18241 26341 18275
rect 26341 18241 26375 18275
rect 26375 18241 26384 18275
rect 26332 18232 26384 18241
rect 28080 18232 28132 18284
rect 28448 18232 28500 18284
rect 20260 18164 20312 18173
rect 21180 18164 21232 18216
rect 22008 18207 22060 18216
rect 21364 18096 21416 18148
rect 22008 18173 22017 18207
rect 22017 18173 22051 18207
rect 22051 18173 22060 18207
rect 22008 18164 22060 18173
rect 22928 18096 22980 18148
rect 23296 18139 23348 18148
rect 23296 18105 23305 18139
rect 23305 18105 23339 18139
rect 23339 18105 23348 18139
rect 23296 18096 23348 18105
rect 20720 18028 20772 18080
rect 21180 18071 21232 18080
rect 21180 18037 21189 18071
rect 21189 18037 21223 18071
rect 21223 18037 21232 18071
rect 21180 18028 21232 18037
rect 25964 18071 26016 18080
rect 25964 18037 25973 18071
rect 25973 18037 26007 18071
rect 26007 18037 26016 18071
rect 25964 18028 26016 18037
rect 26424 18028 26476 18080
rect 28172 18071 28224 18080
rect 28172 18037 28181 18071
rect 28181 18037 28215 18071
rect 28215 18037 28224 18071
rect 28172 18028 28224 18037
rect 5582 17926 5634 17978
rect 5646 17926 5698 17978
rect 5710 17926 5762 17978
rect 5774 17926 5826 17978
rect 5838 17926 5890 17978
rect 14846 17926 14898 17978
rect 14910 17926 14962 17978
rect 14974 17926 15026 17978
rect 15038 17926 15090 17978
rect 15102 17926 15154 17978
rect 24110 17926 24162 17978
rect 24174 17926 24226 17978
rect 24238 17926 24290 17978
rect 24302 17926 24354 17978
rect 24366 17926 24418 17978
rect 7104 17824 7156 17876
rect 7196 17824 7248 17876
rect 8852 17824 8904 17876
rect 1400 17799 1452 17808
rect 1400 17765 1409 17799
rect 1409 17765 1443 17799
rect 1443 17765 1452 17799
rect 1400 17756 1452 17765
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 8944 17756 8996 17808
rect 7196 17620 7248 17629
rect 8392 17688 8444 17740
rect 11980 17824 12032 17876
rect 15200 17867 15252 17876
rect 15200 17833 15209 17867
rect 15209 17833 15243 17867
rect 15243 17833 15252 17867
rect 15200 17824 15252 17833
rect 15660 17824 15712 17876
rect 16396 17756 16448 17808
rect 12164 17688 12216 17740
rect 14096 17688 14148 17740
rect 8300 17620 8352 17672
rect 9220 17663 9272 17672
rect 9220 17629 9254 17663
rect 9254 17629 9272 17663
rect 9220 17620 9272 17629
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 12440 17620 12492 17672
rect 13728 17663 13780 17672
rect 11336 17552 11388 17604
rect 12624 17552 12676 17604
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 14280 17552 14332 17604
rect 7656 17484 7708 17536
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 9956 17484 10008 17536
rect 10784 17527 10836 17536
rect 10784 17493 10793 17527
rect 10793 17493 10827 17527
rect 10827 17493 10836 17527
rect 10784 17484 10836 17493
rect 11888 17484 11940 17536
rect 12348 17484 12400 17536
rect 13360 17527 13412 17536
rect 13360 17493 13369 17527
rect 13369 17493 13403 17527
rect 13403 17493 13412 17527
rect 13360 17484 13412 17493
rect 13452 17484 13504 17536
rect 14556 17663 14608 17672
rect 14556 17629 14565 17663
rect 14565 17629 14599 17663
rect 14599 17629 14608 17663
rect 14832 17688 14884 17740
rect 15568 17731 15620 17740
rect 14556 17620 14608 17629
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 15568 17697 15577 17731
rect 15577 17697 15611 17731
rect 15611 17697 15620 17731
rect 15568 17688 15620 17697
rect 17500 17824 17552 17876
rect 18512 17867 18564 17876
rect 18512 17833 18521 17867
rect 18521 17833 18555 17867
rect 18555 17833 18564 17867
rect 18512 17824 18564 17833
rect 15844 17620 15896 17672
rect 16212 17663 16264 17672
rect 16212 17629 16221 17663
rect 16221 17629 16255 17663
rect 16255 17629 16264 17663
rect 16212 17620 16264 17629
rect 16396 17620 16448 17672
rect 16488 17552 16540 17604
rect 16856 17595 16908 17604
rect 15936 17484 15988 17536
rect 16028 17484 16080 17536
rect 16856 17561 16865 17595
rect 16865 17561 16899 17595
rect 16899 17561 16908 17595
rect 16856 17552 16908 17561
rect 17040 17552 17092 17604
rect 17224 17552 17276 17604
rect 18604 17484 18656 17536
rect 19248 17552 19300 17604
rect 21916 17824 21968 17876
rect 23848 17824 23900 17876
rect 25504 17824 25556 17876
rect 28080 17824 28132 17876
rect 21916 17688 21968 17740
rect 19892 17620 19944 17672
rect 20168 17620 20220 17672
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 20812 17620 20864 17672
rect 22008 17663 22060 17672
rect 22008 17629 22017 17663
rect 22017 17629 22051 17663
rect 22051 17629 22060 17663
rect 22008 17620 22060 17629
rect 22100 17620 22152 17672
rect 23664 17688 23716 17740
rect 24492 17688 24544 17740
rect 23112 17663 23164 17672
rect 23112 17629 23121 17663
rect 23121 17629 23155 17663
rect 23155 17629 23164 17663
rect 23112 17620 23164 17629
rect 24860 17663 24912 17672
rect 20996 17484 21048 17536
rect 21548 17484 21600 17536
rect 23204 17484 23256 17536
rect 24860 17629 24869 17663
rect 24869 17629 24903 17663
rect 24903 17629 24912 17663
rect 24860 17620 24912 17629
rect 25964 17620 26016 17672
rect 25136 17552 25188 17604
rect 25504 17595 25556 17604
rect 25504 17561 25513 17595
rect 25513 17561 25547 17595
rect 25547 17561 25556 17595
rect 25504 17552 25556 17561
rect 25688 17552 25740 17604
rect 26240 17620 26292 17672
rect 26424 17620 26476 17672
rect 26884 17620 26936 17672
rect 25872 17484 25924 17536
rect 26332 17527 26384 17536
rect 26332 17493 26341 17527
rect 26341 17493 26375 17527
rect 26375 17493 26384 17527
rect 26332 17484 26384 17493
rect 10214 17382 10266 17434
rect 10278 17382 10330 17434
rect 10342 17382 10394 17434
rect 10406 17382 10458 17434
rect 10470 17382 10522 17434
rect 19478 17382 19530 17434
rect 19542 17382 19594 17434
rect 19606 17382 19658 17434
rect 19670 17382 19722 17434
rect 19734 17382 19786 17434
rect 7380 17323 7432 17332
rect 7380 17289 7389 17323
rect 7389 17289 7423 17323
rect 7423 17289 7432 17323
rect 7380 17280 7432 17289
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 7196 17144 7248 17196
rect 8944 17144 8996 17196
rect 11060 17144 11112 17196
rect 11336 17144 11388 17196
rect 12624 17280 12676 17332
rect 13084 17280 13136 17332
rect 14832 17280 14884 17332
rect 15108 17280 15160 17332
rect 16672 17323 16724 17332
rect 16672 17289 16681 17323
rect 16681 17289 16715 17323
rect 16715 17289 16724 17323
rect 16672 17280 16724 17289
rect 14556 17212 14608 17264
rect 7104 17076 7156 17128
rect 7656 17119 7708 17128
rect 7656 17085 7665 17119
rect 7665 17085 7699 17119
rect 7699 17085 7708 17119
rect 7656 17076 7708 17085
rect 8392 17119 8444 17128
rect 8392 17085 8401 17119
rect 8401 17085 8435 17119
rect 8435 17085 8444 17119
rect 8392 17076 8444 17085
rect 6000 16940 6052 16992
rect 6736 16940 6788 16992
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 12072 17144 12124 17196
rect 12716 17144 12768 17196
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 13452 17144 13504 17196
rect 13728 17144 13780 17196
rect 14280 17144 14332 17196
rect 14648 17187 14700 17196
rect 14648 17153 14657 17187
rect 14657 17153 14691 17187
rect 14691 17153 14700 17187
rect 14648 17144 14700 17153
rect 15752 17212 15804 17264
rect 12440 17076 12492 17128
rect 13912 17076 13964 17128
rect 15476 17144 15528 17196
rect 16212 17187 16264 17196
rect 16212 17153 16221 17187
rect 16221 17153 16255 17187
rect 16255 17153 16264 17187
rect 16212 17144 16264 17153
rect 17408 17280 17460 17332
rect 17132 17212 17184 17264
rect 20720 17280 20772 17332
rect 26424 17280 26476 17332
rect 28172 17323 28224 17332
rect 28172 17289 28181 17323
rect 28181 17289 28215 17323
rect 28215 17289 28224 17323
rect 28172 17280 28224 17289
rect 17776 17076 17828 17128
rect 11888 17008 11940 17060
rect 11980 16940 12032 16992
rect 14004 16983 14056 16992
rect 14004 16949 14013 16983
rect 14013 16949 14047 16983
rect 14047 16949 14056 16983
rect 14004 16940 14056 16949
rect 14280 16983 14332 16992
rect 14280 16949 14289 16983
rect 14289 16949 14323 16983
rect 14323 16949 14332 16983
rect 14280 16940 14332 16949
rect 14464 16940 14516 16992
rect 16212 16940 16264 16992
rect 17960 17187 18012 17196
rect 17960 17153 17969 17187
rect 17969 17153 18003 17187
rect 18003 17153 18012 17187
rect 17960 17144 18012 17153
rect 19800 17212 19852 17264
rect 19340 17187 19392 17196
rect 19340 17153 19349 17187
rect 19349 17153 19383 17187
rect 19383 17153 19392 17187
rect 19340 17144 19392 17153
rect 19708 17144 19760 17196
rect 19984 17212 20036 17264
rect 20260 17255 20312 17264
rect 20260 17221 20269 17255
rect 20269 17221 20303 17255
rect 20303 17221 20312 17255
rect 20260 17212 20312 17221
rect 22468 17212 22520 17264
rect 20076 17187 20128 17196
rect 20076 17153 20085 17187
rect 20085 17153 20119 17187
rect 20119 17153 20128 17187
rect 20076 17144 20128 17153
rect 20720 17187 20772 17196
rect 20720 17153 20729 17187
rect 20729 17153 20763 17187
rect 20763 17153 20772 17187
rect 20720 17144 20772 17153
rect 19892 17076 19944 17128
rect 21916 17144 21968 17196
rect 21364 17076 21416 17128
rect 23112 17144 23164 17196
rect 24584 17187 24636 17196
rect 24584 17153 24593 17187
rect 24593 17153 24627 17187
rect 24627 17153 24636 17187
rect 24584 17144 24636 17153
rect 25780 17212 25832 17264
rect 28264 17212 28316 17264
rect 24952 17144 25004 17196
rect 25320 17144 25372 17196
rect 24492 17076 24544 17128
rect 21916 17008 21968 17060
rect 22376 17008 22428 17060
rect 25136 17076 25188 17128
rect 28356 17187 28408 17196
rect 28356 17153 28365 17187
rect 28365 17153 28399 17187
rect 28399 17153 28408 17187
rect 28356 17144 28408 17153
rect 26056 17076 26108 17128
rect 26424 17008 26476 17060
rect 18696 16940 18748 16992
rect 18880 16940 18932 16992
rect 20720 16940 20772 16992
rect 21088 16940 21140 16992
rect 23388 16940 23440 16992
rect 24952 16940 25004 16992
rect 25412 16940 25464 16992
rect 25688 16940 25740 16992
rect 26148 16940 26200 16992
rect 5582 16838 5634 16890
rect 5646 16838 5698 16890
rect 5710 16838 5762 16890
rect 5774 16838 5826 16890
rect 5838 16838 5890 16890
rect 14846 16838 14898 16890
rect 14910 16838 14962 16890
rect 14974 16838 15026 16890
rect 15038 16838 15090 16890
rect 15102 16838 15154 16890
rect 24110 16838 24162 16890
rect 24174 16838 24226 16890
rect 24238 16838 24290 16890
rect 24302 16838 24354 16890
rect 24366 16838 24418 16890
rect 8392 16736 8444 16788
rect 8944 16779 8996 16788
rect 8944 16745 8953 16779
rect 8953 16745 8987 16779
rect 8987 16745 8996 16779
rect 8944 16736 8996 16745
rect 11428 16736 11480 16788
rect 12808 16736 12860 16788
rect 13360 16736 13412 16788
rect 15292 16736 15344 16788
rect 16212 16736 16264 16788
rect 20444 16736 20496 16788
rect 23848 16736 23900 16788
rect 25412 16736 25464 16788
rect 28264 16779 28316 16788
rect 28264 16745 28273 16779
rect 28273 16745 28307 16779
rect 28307 16745 28316 16779
rect 28264 16736 28316 16745
rect 8576 16668 8628 16720
rect 7380 16600 7432 16652
rect 11704 16668 11756 16720
rect 6000 16575 6052 16584
rect 6000 16541 6034 16575
rect 6034 16541 6052 16575
rect 6000 16532 6052 16541
rect 8208 16532 8260 16584
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 12716 16668 12768 16720
rect 13636 16668 13688 16720
rect 14188 16668 14240 16720
rect 14556 16668 14608 16720
rect 16304 16711 16356 16720
rect 16304 16677 16313 16711
rect 16313 16677 16347 16711
rect 16347 16677 16356 16711
rect 16304 16668 16356 16677
rect 17224 16711 17276 16720
rect 17224 16677 17233 16711
rect 17233 16677 17267 16711
rect 17267 16677 17276 16711
rect 17224 16668 17276 16677
rect 20904 16668 20956 16720
rect 21824 16668 21876 16720
rect 22008 16711 22060 16720
rect 22008 16677 22017 16711
rect 22017 16677 22051 16711
rect 22051 16677 22060 16711
rect 22008 16668 22060 16677
rect 25136 16668 25188 16720
rect 26240 16668 26292 16720
rect 12808 16643 12860 16652
rect 12808 16609 12817 16643
rect 12817 16609 12851 16643
rect 12851 16609 12860 16643
rect 12808 16600 12860 16609
rect 12992 16600 13044 16652
rect 17500 16643 17552 16652
rect 12348 16532 12400 16584
rect 13084 16532 13136 16584
rect 1492 16396 1544 16448
rect 7104 16439 7156 16448
rect 7104 16405 7113 16439
rect 7113 16405 7147 16439
rect 7147 16405 7156 16439
rect 7104 16396 7156 16405
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 9772 16396 9824 16448
rect 11888 16464 11940 16516
rect 11796 16396 11848 16448
rect 12440 16464 12492 16516
rect 13820 16396 13872 16448
rect 14556 16575 14608 16584
rect 14556 16541 14565 16575
rect 14565 16541 14599 16575
rect 14599 16541 14608 16575
rect 17500 16609 17509 16643
rect 17509 16609 17543 16643
rect 17543 16609 17552 16643
rect 17500 16600 17552 16609
rect 19248 16643 19300 16652
rect 19248 16609 19257 16643
rect 19257 16609 19291 16643
rect 19291 16609 19300 16643
rect 19248 16600 19300 16609
rect 19708 16600 19760 16652
rect 19892 16600 19944 16652
rect 20260 16600 20312 16652
rect 14556 16532 14608 16541
rect 16764 16532 16816 16584
rect 19340 16532 19392 16584
rect 19800 16532 19852 16584
rect 21640 16532 21692 16584
rect 15016 16507 15068 16516
rect 15016 16473 15025 16507
rect 15025 16473 15059 16507
rect 15059 16473 15068 16507
rect 15016 16464 15068 16473
rect 18788 16464 18840 16516
rect 15200 16396 15252 16448
rect 15752 16396 15804 16448
rect 21180 16464 21232 16516
rect 20720 16396 20772 16448
rect 21456 16396 21508 16448
rect 23480 16396 23532 16448
rect 25044 16532 25096 16584
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 26148 16575 26200 16584
rect 26148 16541 26157 16575
rect 26157 16541 26191 16575
rect 26191 16541 26200 16575
rect 26148 16532 26200 16541
rect 26332 16532 26384 16584
rect 26884 16575 26936 16584
rect 26424 16507 26476 16516
rect 26424 16473 26433 16507
rect 26433 16473 26467 16507
rect 26467 16473 26476 16507
rect 26424 16464 26476 16473
rect 26884 16541 26893 16575
rect 26893 16541 26927 16575
rect 26927 16541 26936 16575
rect 26884 16532 26936 16541
rect 25504 16396 25556 16448
rect 10214 16294 10266 16346
rect 10278 16294 10330 16346
rect 10342 16294 10394 16346
rect 10406 16294 10458 16346
rect 10470 16294 10522 16346
rect 19478 16294 19530 16346
rect 19542 16294 19594 16346
rect 19606 16294 19658 16346
rect 19670 16294 19722 16346
rect 19734 16294 19786 16346
rect 9128 16192 9180 16244
rect 9956 16235 10008 16244
rect 9956 16201 9965 16235
rect 9965 16201 9999 16235
rect 9999 16201 10008 16235
rect 9956 16192 10008 16201
rect 11152 16235 11204 16244
rect 11152 16201 11161 16235
rect 11161 16201 11195 16235
rect 11195 16201 11204 16235
rect 11152 16192 11204 16201
rect 13728 16192 13780 16244
rect 13820 16192 13872 16244
rect 10692 16124 10744 16176
rect 15016 16124 15068 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 5908 16056 5960 16108
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 7840 16056 7892 16108
rect 9220 15988 9272 16040
rect 11060 16056 11112 16108
rect 11796 16099 11848 16108
rect 11796 16065 11830 16099
rect 11830 16065 11848 16099
rect 11796 16056 11848 16065
rect 13084 16056 13136 16108
rect 14280 16056 14332 16108
rect 14464 16056 14516 16108
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 16028 16099 16080 16108
rect 16028 16065 16037 16099
rect 16037 16065 16071 16099
rect 16071 16065 16080 16099
rect 16028 16056 16080 16065
rect 9956 15988 10008 16040
rect 13636 16031 13688 16040
rect 9588 15920 9640 15972
rect 13636 15997 13645 16031
rect 13645 15997 13679 16031
rect 13679 15997 13688 16031
rect 13636 15988 13688 15997
rect 17684 16124 17736 16176
rect 17868 16192 17920 16244
rect 18788 16192 18840 16244
rect 20076 16192 20128 16244
rect 21456 16235 21508 16244
rect 21456 16201 21465 16235
rect 21465 16201 21499 16235
rect 21499 16201 21508 16235
rect 21456 16192 21508 16201
rect 21088 16124 21140 16176
rect 22008 16124 22060 16176
rect 17132 16056 17184 16108
rect 14372 15920 14424 15972
rect 14648 15920 14700 15972
rect 17684 16031 17736 16040
rect 17684 15997 17693 16031
rect 17693 15997 17727 16031
rect 17727 15997 17736 16031
rect 17684 15988 17736 15997
rect 17868 15920 17920 15972
rect 19340 16056 19392 16108
rect 20812 16099 20864 16108
rect 19984 15988 20036 16040
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 20904 16099 20956 16108
rect 20904 16065 20913 16099
rect 20913 16065 20947 16099
rect 20947 16065 20956 16099
rect 21272 16099 21324 16108
rect 20904 16056 20956 16065
rect 21272 16065 21281 16099
rect 21281 16065 21315 16099
rect 21315 16065 21324 16099
rect 21272 16056 21324 16065
rect 23480 16099 23532 16108
rect 23480 16065 23489 16099
rect 23489 16065 23523 16099
rect 23523 16065 23532 16099
rect 23480 16056 23532 16065
rect 23572 16099 23624 16108
rect 23572 16065 23581 16099
rect 23581 16065 23615 16099
rect 23615 16065 23624 16099
rect 23572 16056 23624 16065
rect 23848 16056 23900 16108
rect 26884 16124 26936 16176
rect 25780 16099 25832 16108
rect 25780 16065 25789 16099
rect 25789 16065 25823 16099
rect 25823 16065 25832 16099
rect 25780 16056 25832 16065
rect 26148 16099 26200 16108
rect 5448 15895 5500 15904
rect 5448 15861 5457 15895
rect 5457 15861 5491 15895
rect 5491 15861 5500 15895
rect 5448 15852 5500 15861
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 10140 15852 10192 15904
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 12256 15852 12308 15904
rect 12992 15852 13044 15904
rect 13176 15895 13228 15904
rect 13176 15861 13185 15895
rect 13185 15861 13219 15895
rect 13219 15861 13228 15895
rect 13176 15852 13228 15861
rect 15292 15852 15344 15904
rect 16948 15852 17000 15904
rect 17316 15852 17368 15904
rect 20444 15895 20496 15904
rect 20444 15861 20453 15895
rect 20453 15861 20487 15895
rect 20487 15861 20496 15895
rect 20444 15852 20496 15861
rect 25412 15988 25464 16040
rect 26148 16065 26157 16099
rect 26157 16065 26191 16099
rect 26191 16065 26200 16099
rect 26148 16056 26200 16065
rect 26240 16099 26292 16108
rect 26240 16065 26249 16099
rect 26249 16065 26283 16099
rect 26283 16065 26292 16099
rect 26240 16056 26292 16065
rect 26884 15988 26936 16040
rect 22284 15852 22336 15904
rect 25228 15852 25280 15904
rect 28356 15895 28408 15904
rect 28356 15861 28365 15895
rect 28365 15861 28399 15895
rect 28399 15861 28408 15895
rect 28356 15852 28408 15861
rect 5582 15750 5634 15802
rect 5646 15750 5698 15802
rect 5710 15750 5762 15802
rect 5774 15750 5826 15802
rect 5838 15750 5890 15802
rect 14846 15750 14898 15802
rect 14910 15750 14962 15802
rect 14974 15750 15026 15802
rect 15038 15750 15090 15802
rect 15102 15750 15154 15802
rect 24110 15750 24162 15802
rect 24174 15750 24226 15802
rect 24238 15750 24290 15802
rect 24302 15750 24354 15802
rect 24366 15750 24418 15802
rect 11060 15691 11112 15700
rect 11060 15657 11069 15691
rect 11069 15657 11103 15691
rect 11103 15657 11112 15691
rect 11060 15648 11112 15657
rect 11796 15648 11848 15700
rect 5172 15555 5224 15564
rect 5172 15521 5181 15555
rect 5181 15521 5215 15555
rect 5215 15521 5224 15555
rect 5172 15512 5224 15521
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 9588 15512 9640 15564
rect 5448 15487 5500 15496
rect 5448 15453 5482 15487
rect 5482 15453 5500 15487
rect 5448 15444 5500 15453
rect 7748 15444 7800 15496
rect 6828 15308 6880 15360
rect 7196 15351 7248 15360
rect 7196 15317 7205 15351
rect 7205 15317 7239 15351
rect 7239 15317 7248 15351
rect 7196 15308 7248 15317
rect 10048 15376 10100 15428
rect 11704 15623 11756 15632
rect 11704 15589 11713 15623
rect 11713 15589 11747 15623
rect 11747 15589 11756 15623
rect 11704 15580 11756 15589
rect 12440 15648 12492 15700
rect 13636 15648 13688 15700
rect 16212 15648 16264 15700
rect 17776 15648 17828 15700
rect 21640 15691 21692 15700
rect 21640 15657 21649 15691
rect 21649 15657 21683 15691
rect 21683 15657 21692 15691
rect 21640 15648 21692 15657
rect 23572 15648 23624 15700
rect 24860 15691 24912 15700
rect 24860 15657 24869 15691
rect 24869 15657 24903 15691
rect 24903 15657 24912 15691
rect 24860 15648 24912 15657
rect 25044 15648 25096 15700
rect 25504 15691 25556 15700
rect 25504 15657 25513 15691
rect 25513 15657 25547 15691
rect 25547 15657 25556 15691
rect 25504 15648 25556 15657
rect 12256 15580 12308 15632
rect 12808 15580 12860 15632
rect 12992 15580 13044 15632
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 11428 15444 11480 15496
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 14004 15512 14056 15564
rect 12532 15444 12584 15496
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 13452 15487 13504 15496
rect 13452 15453 13461 15487
rect 13461 15453 13495 15487
rect 13495 15453 13504 15487
rect 13452 15444 13504 15453
rect 13728 15444 13780 15496
rect 14372 15487 14424 15496
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 14464 15444 14516 15496
rect 15200 15512 15252 15564
rect 15292 15444 15344 15496
rect 15384 15444 15436 15496
rect 15936 15512 15988 15564
rect 16856 15580 16908 15632
rect 16948 15580 17000 15632
rect 16580 15487 16632 15496
rect 16580 15453 16589 15487
rect 16589 15453 16623 15487
rect 16623 15453 16632 15487
rect 16580 15444 16632 15453
rect 17316 15487 17368 15496
rect 17316 15453 17325 15487
rect 17325 15453 17359 15487
rect 17359 15453 17368 15487
rect 17868 15512 17920 15564
rect 17316 15444 17368 15453
rect 19892 15512 19944 15564
rect 21272 15512 21324 15564
rect 21732 15512 21784 15564
rect 18788 15487 18840 15496
rect 18788 15453 18797 15487
rect 18797 15453 18831 15487
rect 18831 15453 18840 15487
rect 18788 15444 18840 15453
rect 19984 15487 20036 15496
rect 12716 15308 12768 15360
rect 15200 15376 15252 15428
rect 15660 15419 15712 15428
rect 15660 15385 15669 15419
rect 15669 15385 15703 15419
rect 15703 15385 15712 15419
rect 15660 15376 15712 15385
rect 16396 15376 16448 15428
rect 16856 15419 16908 15428
rect 16856 15385 16865 15419
rect 16865 15385 16899 15419
rect 16899 15385 16908 15419
rect 16856 15376 16908 15385
rect 17224 15376 17276 15428
rect 13452 15308 13504 15360
rect 13544 15308 13596 15360
rect 16764 15308 16816 15360
rect 17408 15376 17460 15428
rect 17960 15419 18012 15428
rect 17592 15351 17644 15360
rect 17592 15317 17601 15351
rect 17601 15317 17635 15351
rect 17635 15317 17644 15351
rect 17592 15308 17644 15317
rect 17960 15385 17969 15419
rect 17969 15385 18003 15419
rect 18003 15385 18012 15419
rect 17960 15376 18012 15385
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 20996 15444 21048 15496
rect 26148 15512 26200 15564
rect 18604 15351 18656 15360
rect 18604 15317 18613 15351
rect 18613 15317 18647 15351
rect 18647 15317 18656 15351
rect 18604 15308 18656 15317
rect 19892 15376 19944 15428
rect 20260 15419 20312 15428
rect 20260 15385 20294 15419
rect 20294 15385 20312 15419
rect 20260 15376 20312 15385
rect 20812 15376 20864 15428
rect 22284 15444 22336 15496
rect 24952 15487 25004 15496
rect 24952 15453 24961 15487
rect 24961 15453 24995 15487
rect 24995 15453 25004 15487
rect 24952 15444 25004 15453
rect 26516 15487 26568 15496
rect 22560 15376 22612 15428
rect 24860 15376 24912 15428
rect 25596 15376 25648 15428
rect 26516 15453 26525 15487
rect 26525 15453 26559 15487
rect 26559 15453 26568 15487
rect 26516 15444 26568 15453
rect 26884 15648 26936 15700
rect 26792 15580 26844 15632
rect 26056 15376 26108 15428
rect 28356 15512 28408 15564
rect 20536 15308 20588 15360
rect 21364 15351 21416 15360
rect 21364 15317 21373 15351
rect 21373 15317 21407 15351
rect 21407 15317 21416 15351
rect 21364 15308 21416 15317
rect 26792 15308 26844 15360
rect 26976 15308 27028 15360
rect 28264 15351 28316 15360
rect 28264 15317 28273 15351
rect 28273 15317 28307 15351
rect 28307 15317 28316 15351
rect 28264 15308 28316 15317
rect 10214 15206 10266 15258
rect 10278 15206 10330 15258
rect 10342 15206 10394 15258
rect 10406 15206 10458 15258
rect 10470 15206 10522 15258
rect 19478 15206 19530 15258
rect 19542 15206 19594 15258
rect 19606 15206 19658 15258
rect 19670 15206 19722 15258
rect 19734 15206 19786 15258
rect 4068 15104 4120 15156
rect 10692 15104 10744 15156
rect 12256 15104 12308 15156
rect 13728 15104 13780 15156
rect 14372 15104 14424 15156
rect 14740 15104 14792 15156
rect 15660 15104 15712 15156
rect 16672 15104 16724 15156
rect 17868 15104 17920 15156
rect 5908 15036 5960 15088
rect 7196 15036 7248 15088
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 7104 14968 7156 15020
rect 9404 15011 9456 15020
rect 9404 14977 9413 15011
rect 9413 14977 9447 15011
rect 9447 14977 9456 15011
rect 9404 14968 9456 14977
rect 10140 14968 10192 15020
rect 12072 15011 12124 15020
rect 12072 14977 12081 15011
rect 12081 14977 12115 15011
rect 12115 14977 12124 15011
rect 12072 14968 12124 14977
rect 12624 15036 12676 15088
rect 12716 15011 12768 15020
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 8208 14943 8260 14952
rect 6736 14832 6788 14884
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 9220 14943 9272 14952
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 11796 14900 11848 14952
rect 12348 14900 12400 14952
rect 12716 14977 12725 15011
rect 12725 14977 12759 15011
rect 12759 14977 12768 15011
rect 12716 14968 12768 14977
rect 13084 14968 13136 15020
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 13452 15011 13504 15020
rect 13452 14977 13462 15011
rect 13462 14977 13496 15011
rect 13496 14977 13504 15011
rect 13636 15011 13688 15020
rect 13452 14968 13504 14977
rect 13636 14977 13645 15011
rect 13645 14977 13679 15011
rect 13679 14977 13688 15011
rect 13636 14968 13688 14977
rect 13820 15011 13872 15020
rect 13820 14977 13834 15011
rect 13834 14977 13868 15011
rect 13868 14977 13872 15011
rect 13820 14968 13872 14977
rect 14188 14968 14240 15020
rect 14372 15011 14424 15020
rect 14372 14977 14382 15011
rect 14382 14977 14416 15011
rect 14416 14977 14424 15011
rect 14372 14968 14424 14977
rect 14004 14900 14056 14952
rect 7564 14875 7616 14884
rect 7564 14841 7573 14875
rect 7573 14841 7607 14875
rect 7607 14841 7616 14875
rect 7564 14832 7616 14841
rect 10048 14832 10100 14884
rect 13084 14875 13136 14884
rect 10140 14807 10192 14816
rect 10140 14773 10149 14807
rect 10149 14773 10183 14807
rect 10183 14773 10192 14807
rect 10140 14764 10192 14773
rect 11796 14764 11848 14816
rect 13084 14841 13093 14875
rect 13093 14841 13127 14875
rect 13127 14841 13136 14875
rect 13084 14832 13136 14841
rect 12900 14764 12952 14816
rect 13636 14764 13688 14816
rect 15200 14968 15252 15020
rect 16764 14968 16816 15020
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 17316 14968 17368 15020
rect 15384 14943 15436 14952
rect 15384 14909 15393 14943
rect 15393 14909 15427 14943
rect 15427 14909 15436 14943
rect 15384 14900 15436 14909
rect 17776 14900 17828 14952
rect 16580 14832 16632 14884
rect 14280 14764 14332 14816
rect 14372 14764 14424 14816
rect 15292 14764 15344 14816
rect 19892 15104 19944 15156
rect 21732 15104 21784 15156
rect 22560 15147 22612 15156
rect 22560 15113 22569 15147
rect 22569 15113 22603 15147
rect 22603 15113 22612 15147
rect 22560 15104 22612 15113
rect 19984 15036 20036 15088
rect 20628 15036 20680 15088
rect 18604 15011 18656 15020
rect 18604 14977 18638 15011
rect 18638 14977 18656 15011
rect 18604 14968 18656 14977
rect 20352 14968 20404 15020
rect 20444 15011 20496 15020
rect 20444 14977 20453 15011
rect 20453 14977 20487 15011
rect 20487 14977 20496 15011
rect 21364 15036 21416 15088
rect 22100 15036 22152 15088
rect 20444 14968 20496 14977
rect 18328 14943 18380 14952
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 18328 14900 18380 14909
rect 19708 14900 19760 14952
rect 20076 14900 20128 14952
rect 21732 14968 21784 15020
rect 22560 14900 22612 14952
rect 18512 14764 18564 14816
rect 19708 14807 19760 14816
rect 19708 14773 19717 14807
rect 19717 14773 19751 14807
rect 19751 14773 19760 14807
rect 19708 14764 19760 14773
rect 20260 14832 20312 14884
rect 20536 14832 20588 14884
rect 26792 15036 26844 15088
rect 23664 14968 23716 15020
rect 20904 14764 20956 14816
rect 23388 14764 23440 14816
rect 24032 14764 24084 14816
rect 26056 14968 26108 15020
rect 27252 15011 27304 15020
rect 27252 14977 27286 15011
rect 27286 14977 27304 15011
rect 27252 14968 27304 14977
rect 25596 14943 25648 14952
rect 25228 14832 25280 14884
rect 25596 14909 25605 14943
rect 25605 14909 25639 14943
rect 25639 14909 25648 14943
rect 25596 14900 25648 14909
rect 26148 14900 26200 14952
rect 25872 14832 25924 14884
rect 25044 14807 25096 14816
rect 25044 14773 25053 14807
rect 25053 14773 25087 14807
rect 25087 14773 25096 14807
rect 25044 14764 25096 14773
rect 28356 14807 28408 14816
rect 28356 14773 28365 14807
rect 28365 14773 28399 14807
rect 28399 14773 28408 14807
rect 28356 14764 28408 14773
rect 5582 14662 5634 14714
rect 5646 14662 5698 14714
rect 5710 14662 5762 14714
rect 5774 14662 5826 14714
rect 5838 14662 5890 14714
rect 14846 14662 14898 14714
rect 14910 14662 14962 14714
rect 14974 14662 15026 14714
rect 15038 14662 15090 14714
rect 15102 14662 15154 14714
rect 24110 14662 24162 14714
rect 24174 14662 24226 14714
rect 24238 14662 24290 14714
rect 24302 14662 24354 14714
rect 24366 14662 24418 14714
rect 11612 14560 11664 14612
rect 13452 14560 13504 14612
rect 17224 14560 17276 14612
rect 18788 14560 18840 14612
rect 9220 14424 9272 14476
rect 9772 14424 9824 14476
rect 7564 14399 7616 14408
rect 7564 14365 7573 14399
rect 7573 14365 7607 14399
rect 7607 14365 7616 14399
rect 7564 14356 7616 14365
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 10140 14356 10192 14408
rect 12164 14492 12216 14544
rect 13820 14492 13872 14544
rect 12072 14424 12124 14476
rect 15292 14492 15344 14544
rect 15384 14492 15436 14544
rect 18420 14492 18472 14544
rect 19156 14492 19208 14544
rect 14188 14424 14240 14476
rect 14464 14424 14516 14476
rect 13360 14356 13412 14408
rect 14096 14399 14148 14408
rect 9312 14288 9364 14340
rect 5908 14220 5960 14272
rect 6552 14220 6604 14272
rect 8024 14263 8076 14272
rect 8024 14229 8033 14263
rect 8033 14229 8067 14263
rect 8067 14229 8076 14263
rect 8024 14220 8076 14229
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 11612 14220 11664 14229
rect 12900 14288 12952 14340
rect 13452 14331 13504 14340
rect 13084 14220 13136 14272
rect 13452 14297 13461 14331
rect 13461 14297 13495 14331
rect 13495 14297 13504 14331
rect 13452 14288 13504 14297
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 15200 14356 15252 14408
rect 16120 14424 16172 14476
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 16580 14424 16632 14476
rect 16856 14356 16908 14408
rect 19340 14424 19392 14476
rect 14648 14288 14700 14340
rect 15292 14263 15344 14272
rect 15292 14229 15301 14263
rect 15301 14229 15335 14263
rect 15335 14229 15344 14263
rect 15292 14220 15344 14229
rect 17592 14356 17644 14408
rect 18512 14399 18564 14408
rect 17500 14288 17552 14340
rect 18512 14365 18521 14399
rect 18521 14365 18555 14399
rect 18555 14365 18564 14399
rect 18512 14356 18564 14365
rect 18696 14399 18748 14408
rect 18696 14365 18705 14399
rect 18705 14365 18739 14399
rect 18739 14365 18748 14399
rect 18696 14356 18748 14365
rect 19340 14288 19392 14340
rect 21916 14492 21968 14544
rect 24032 14560 24084 14612
rect 25136 14560 25188 14612
rect 26056 14603 26108 14612
rect 23664 14535 23716 14544
rect 23664 14501 23673 14535
rect 23673 14501 23707 14535
rect 23707 14501 23716 14535
rect 23664 14492 23716 14501
rect 26056 14569 26065 14603
rect 26065 14569 26099 14603
rect 26099 14569 26108 14603
rect 26056 14560 26108 14569
rect 27252 14560 27304 14612
rect 20260 14356 20312 14408
rect 20444 14399 20496 14408
rect 20444 14365 20453 14399
rect 20453 14365 20487 14399
rect 20487 14365 20496 14399
rect 20444 14356 20496 14365
rect 20996 14356 21048 14408
rect 22008 14399 22060 14408
rect 22008 14365 22017 14399
rect 22017 14365 22051 14399
rect 22051 14365 22060 14399
rect 22008 14356 22060 14365
rect 22100 14356 22152 14408
rect 22468 14356 22520 14408
rect 23296 14399 23348 14408
rect 23296 14365 23305 14399
rect 23305 14365 23339 14399
rect 23339 14365 23348 14399
rect 23296 14356 23348 14365
rect 24584 14424 24636 14476
rect 25504 14424 25556 14476
rect 25044 14399 25096 14408
rect 23020 14288 23072 14340
rect 23204 14288 23256 14340
rect 25044 14365 25053 14399
rect 25053 14365 25087 14399
rect 25087 14365 25096 14399
rect 25044 14356 25096 14365
rect 17132 14220 17184 14272
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 20904 14220 20956 14272
rect 21640 14220 21692 14272
rect 22100 14220 22152 14272
rect 22560 14220 22612 14272
rect 24860 14288 24912 14340
rect 26516 14356 26568 14408
rect 26792 14399 26844 14408
rect 26792 14365 26801 14399
rect 26801 14365 26835 14399
rect 26835 14365 26844 14399
rect 26792 14356 26844 14365
rect 26976 14399 27028 14408
rect 26976 14365 26985 14399
rect 26985 14365 27019 14399
rect 27019 14365 27028 14399
rect 26976 14356 27028 14365
rect 27068 14399 27120 14408
rect 27068 14365 27077 14399
rect 27077 14365 27111 14399
rect 27111 14365 27120 14399
rect 27068 14356 27120 14365
rect 25872 14331 25924 14340
rect 25872 14297 25881 14331
rect 25881 14297 25915 14331
rect 25915 14297 25924 14331
rect 25872 14288 25924 14297
rect 28356 14356 28408 14408
rect 27896 14331 27948 14340
rect 27896 14297 27905 14331
rect 27905 14297 27939 14331
rect 27939 14297 27948 14331
rect 27896 14288 27948 14297
rect 23848 14220 23900 14272
rect 24216 14220 24268 14272
rect 25044 14220 25096 14272
rect 25504 14263 25556 14272
rect 25504 14229 25513 14263
rect 25513 14229 25547 14263
rect 25547 14229 25556 14263
rect 25504 14220 25556 14229
rect 26332 14263 26384 14272
rect 26332 14229 26341 14263
rect 26341 14229 26375 14263
rect 26375 14229 26384 14263
rect 26332 14220 26384 14229
rect 10214 14118 10266 14170
rect 10278 14118 10330 14170
rect 10342 14118 10394 14170
rect 10406 14118 10458 14170
rect 10470 14118 10522 14170
rect 19478 14118 19530 14170
rect 19542 14118 19594 14170
rect 19606 14118 19658 14170
rect 19670 14118 19722 14170
rect 19734 14118 19786 14170
rect 5908 14016 5960 14068
rect 8944 14059 8996 14068
rect 8944 14025 8953 14059
rect 8953 14025 8987 14059
rect 8987 14025 8996 14059
rect 8944 14016 8996 14025
rect 9404 14016 9456 14068
rect 11612 14016 11664 14068
rect 6828 13948 6880 14000
rect 8024 13948 8076 14000
rect 8208 13948 8260 14000
rect 6552 13812 6604 13864
rect 10048 13948 10100 14000
rect 10600 13948 10652 14000
rect 12532 14016 12584 14068
rect 12992 14016 13044 14068
rect 13360 14016 13412 14068
rect 13452 14016 13504 14068
rect 18420 14016 18472 14068
rect 20260 14016 20312 14068
rect 11704 13880 11756 13932
rect 14096 13948 14148 14000
rect 14464 13948 14516 14000
rect 15936 13948 15988 14000
rect 16212 13948 16264 14000
rect 17500 13948 17552 14000
rect 18328 13948 18380 14000
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 13084 13923 13136 13932
rect 13084 13889 13094 13923
rect 13094 13889 13128 13923
rect 13128 13889 13136 13923
rect 13084 13880 13136 13889
rect 6736 13744 6788 13796
rect 6644 13676 6696 13728
rect 7196 13676 7248 13728
rect 12348 13812 12400 13864
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 13728 13880 13780 13932
rect 13636 13812 13688 13864
rect 14372 13812 14424 13864
rect 16764 13880 16816 13932
rect 18420 13923 18472 13932
rect 18420 13889 18429 13923
rect 18429 13889 18463 13923
rect 18463 13889 18472 13923
rect 18420 13880 18472 13889
rect 19248 13948 19300 14000
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 20536 13923 20588 13932
rect 20536 13889 20545 13923
rect 20545 13889 20579 13923
rect 20579 13889 20588 13923
rect 21088 13948 21140 14000
rect 20536 13880 20588 13889
rect 20812 13923 20864 13932
rect 20812 13889 20821 13923
rect 20821 13889 20855 13923
rect 20855 13889 20864 13923
rect 20812 13880 20864 13889
rect 11152 13787 11204 13796
rect 7840 13676 7892 13728
rect 11152 13753 11161 13787
rect 11161 13753 11195 13787
rect 11195 13753 11204 13787
rect 11152 13744 11204 13753
rect 14096 13744 14148 13796
rect 16580 13744 16632 13796
rect 17040 13812 17092 13864
rect 21088 13812 21140 13864
rect 21640 14016 21692 14068
rect 22560 14059 22612 14068
rect 22560 14025 22569 14059
rect 22569 14025 22603 14059
rect 22603 14025 22612 14059
rect 23296 14059 23348 14068
rect 22560 14016 22612 14025
rect 23296 14025 23305 14059
rect 23305 14025 23339 14059
rect 23339 14025 23348 14059
rect 23296 14016 23348 14025
rect 23664 14016 23716 14068
rect 21548 13880 21600 13932
rect 21640 13880 21692 13932
rect 22284 13880 22336 13932
rect 23204 13880 23256 13932
rect 24124 14016 24176 14068
rect 24032 13948 24084 14000
rect 24584 13948 24636 14000
rect 24216 13923 24268 13932
rect 23020 13812 23072 13864
rect 23572 13855 23624 13864
rect 23572 13821 23581 13855
rect 23581 13821 23615 13855
rect 23615 13821 23624 13855
rect 23572 13812 23624 13821
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 24676 13880 24728 13932
rect 25872 14016 25924 14068
rect 26792 14016 26844 14068
rect 26332 13991 26384 14000
rect 26332 13957 26341 13991
rect 26341 13957 26375 13991
rect 26375 13957 26384 13991
rect 26332 13948 26384 13957
rect 9772 13676 9824 13728
rect 13912 13676 13964 13728
rect 15292 13676 15344 13728
rect 17132 13676 17184 13728
rect 23296 13744 23348 13796
rect 24584 13812 24636 13864
rect 24860 13855 24912 13864
rect 24860 13821 24869 13855
rect 24869 13821 24903 13855
rect 24903 13821 24912 13855
rect 24860 13812 24912 13821
rect 26240 13923 26292 13932
rect 26240 13889 26249 13923
rect 26249 13889 26283 13923
rect 26283 13889 26292 13923
rect 27896 13948 27948 14000
rect 26240 13880 26292 13889
rect 26976 13923 27028 13932
rect 26976 13889 26985 13923
rect 26985 13889 27019 13923
rect 27019 13889 27028 13923
rect 26976 13880 27028 13889
rect 28264 13923 28316 13932
rect 28264 13889 28273 13923
rect 28273 13889 28307 13923
rect 28307 13889 28316 13923
rect 28264 13880 28316 13889
rect 27068 13812 27120 13864
rect 25688 13744 25740 13796
rect 20628 13676 20680 13728
rect 21456 13719 21508 13728
rect 21456 13685 21465 13719
rect 21465 13685 21499 13719
rect 21499 13685 21508 13719
rect 21456 13676 21508 13685
rect 21732 13676 21784 13728
rect 22284 13719 22336 13728
rect 22284 13685 22293 13719
rect 22293 13685 22327 13719
rect 22327 13685 22336 13719
rect 22284 13676 22336 13685
rect 22376 13676 22428 13728
rect 24492 13676 24544 13728
rect 25044 13719 25096 13728
rect 25044 13685 25053 13719
rect 25053 13685 25087 13719
rect 25087 13685 25096 13719
rect 25044 13676 25096 13685
rect 25964 13719 26016 13728
rect 25964 13685 25973 13719
rect 25973 13685 26007 13719
rect 26007 13685 26016 13719
rect 25964 13676 26016 13685
rect 27160 13719 27212 13728
rect 27160 13685 27169 13719
rect 27169 13685 27203 13719
rect 27203 13685 27212 13719
rect 27160 13676 27212 13685
rect 5582 13574 5634 13626
rect 5646 13574 5698 13626
rect 5710 13574 5762 13626
rect 5774 13574 5826 13626
rect 5838 13574 5890 13626
rect 14846 13574 14898 13626
rect 14910 13574 14962 13626
rect 14974 13574 15026 13626
rect 15038 13574 15090 13626
rect 15102 13574 15154 13626
rect 24110 13574 24162 13626
rect 24174 13574 24226 13626
rect 24238 13574 24290 13626
rect 24302 13574 24354 13626
rect 24366 13574 24418 13626
rect 7196 13515 7248 13524
rect 5172 13336 5224 13388
rect 7196 13481 7205 13515
rect 7205 13481 7239 13515
rect 7239 13481 7248 13515
rect 7196 13472 7248 13481
rect 7564 13472 7616 13524
rect 15844 13472 15896 13524
rect 17132 13472 17184 13524
rect 18604 13472 18656 13524
rect 6736 13336 6788 13388
rect 8208 13379 8260 13388
rect 8208 13345 8217 13379
rect 8217 13345 8251 13379
rect 8251 13345 8260 13379
rect 9680 13404 9732 13456
rect 8208 13336 8260 13345
rect 5908 13268 5960 13320
rect 8944 13268 8996 13320
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 9772 13268 9824 13320
rect 11152 13268 11204 13320
rect 14464 13404 14516 13456
rect 16580 13404 16632 13456
rect 20260 13472 20312 13524
rect 21088 13472 21140 13524
rect 21640 13472 21692 13524
rect 21824 13472 21876 13524
rect 21916 13472 21968 13524
rect 14372 13379 14424 13388
rect 9128 13200 9180 13252
rect 10876 13200 10928 13252
rect 11612 13243 11664 13252
rect 11612 13209 11646 13243
rect 11646 13209 11664 13243
rect 14004 13268 14056 13320
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 15936 13336 15988 13388
rect 16764 13336 16816 13388
rect 11612 13200 11664 13209
rect 10968 13132 11020 13184
rect 11060 13175 11112 13184
rect 11060 13141 11069 13175
rect 11069 13141 11103 13175
rect 11103 13141 11112 13175
rect 13452 13243 13504 13252
rect 13452 13209 13461 13243
rect 13461 13209 13495 13243
rect 13495 13209 13504 13243
rect 14188 13268 14240 13320
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 19892 13404 19944 13456
rect 20076 13404 20128 13456
rect 18420 13336 18472 13388
rect 19800 13336 19852 13388
rect 19984 13336 20036 13388
rect 22284 13472 22336 13524
rect 23664 13472 23716 13524
rect 24032 13472 24084 13524
rect 23572 13404 23624 13456
rect 24676 13472 24728 13524
rect 26976 13472 27028 13524
rect 28448 13472 28500 13524
rect 17132 13268 17184 13277
rect 16212 13243 16264 13252
rect 13452 13200 13504 13209
rect 16212 13209 16221 13243
rect 16221 13209 16255 13243
rect 16255 13209 16264 13243
rect 16212 13200 16264 13209
rect 19340 13268 19392 13320
rect 19892 13268 19944 13320
rect 18512 13200 18564 13252
rect 20444 13200 20496 13252
rect 22744 13268 22796 13320
rect 23204 13268 23256 13320
rect 25044 13336 25096 13388
rect 26148 13336 26200 13388
rect 24400 13311 24452 13320
rect 24400 13277 24409 13311
rect 24409 13277 24443 13311
rect 24443 13277 24452 13311
rect 24400 13268 24452 13277
rect 12716 13175 12768 13184
rect 11060 13132 11112 13141
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 14832 13132 14884 13184
rect 16028 13132 16080 13184
rect 18052 13175 18104 13184
rect 18052 13141 18061 13175
rect 18061 13141 18095 13175
rect 18095 13141 18104 13175
rect 18052 13132 18104 13141
rect 20352 13132 20404 13184
rect 21088 13132 21140 13184
rect 21824 13132 21876 13184
rect 22376 13132 22428 13184
rect 22468 13132 22520 13184
rect 23296 13132 23348 13184
rect 25872 13268 25924 13320
rect 25320 13200 25372 13252
rect 25688 13243 25740 13252
rect 25688 13209 25697 13243
rect 25697 13209 25731 13243
rect 25731 13209 25740 13243
rect 25688 13200 25740 13209
rect 25964 13200 26016 13252
rect 27252 13243 27304 13252
rect 27252 13209 27286 13243
rect 27286 13209 27304 13243
rect 27252 13200 27304 13209
rect 10214 13030 10266 13082
rect 10278 13030 10330 13082
rect 10342 13030 10394 13082
rect 10406 13030 10458 13082
rect 10470 13030 10522 13082
rect 19478 13030 19530 13082
rect 19542 13030 19594 13082
rect 19606 13030 19658 13082
rect 19670 13030 19722 13082
rect 19734 13030 19786 13082
rect 6736 12971 6788 12980
rect 6736 12937 6745 12971
rect 6745 12937 6779 12971
rect 6779 12937 6788 12971
rect 6736 12928 6788 12937
rect 9220 12928 9272 12980
rect 10876 12928 10928 12980
rect 11612 12928 11664 12980
rect 12440 12928 12492 12980
rect 12716 12971 12768 12980
rect 12716 12937 12725 12971
rect 12725 12937 12759 12971
rect 12759 12937 12768 12971
rect 12716 12928 12768 12937
rect 5816 12860 5868 12912
rect 6000 12860 6052 12912
rect 6552 12860 6604 12912
rect 11060 12860 11112 12912
rect 5816 12767 5868 12776
rect 5816 12733 5825 12767
rect 5825 12733 5859 12767
rect 5859 12733 5868 12767
rect 5816 12724 5868 12733
rect 6644 12792 6696 12844
rect 7840 12835 7892 12844
rect 6552 12724 6604 12776
rect 7840 12801 7849 12835
rect 7849 12801 7883 12835
rect 7883 12801 7892 12835
rect 7840 12792 7892 12801
rect 7932 12792 7984 12844
rect 9956 12792 10008 12844
rect 10968 12792 11020 12844
rect 11796 12792 11848 12844
rect 9864 12724 9916 12776
rect 10600 12767 10652 12776
rect 10600 12733 10609 12767
rect 10609 12733 10643 12767
rect 10643 12733 10652 12767
rect 10600 12724 10652 12733
rect 11060 12724 11112 12776
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 9312 12656 9364 12708
rect 9588 12656 9640 12708
rect 14556 12928 14608 12980
rect 15476 12928 15528 12980
rect 14832 12903 14884 12912
rect 14832 12869 14841 12903
rect 14841 12869 14875 12903
rect 14875 12869 14884 12903
rect 14832 12860 14884 12869
rect 14004 12835 14056 12844
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 14004 12801 14013 12835
rect 14013 12801 14047 12835
rect 14047 12801 14056 12835
rect 14004 12792 14056 12801
rect 14096 12835 14148 12844
rect 14096 12801 14110 12835
rect 14110 12801 14144 12835
rect 14144 12801 14148 12835
rect 14096 12792 14148 12801
rect 14464 12792 14516 12844
rect 14648 12835 14700 12844
rect 14648 12801 14658 12835
rect 14658 12801 14692 12835
rect 14692 12801 14700 12835
rect 14648 12792 14700 12801
rect 5264 12588 5316 12640
rect 9404 12588 9456 12640
rect 12808 12588 12860 12640
rect 14188 12656 14240 12708
rect 15108 12656 15160 12708
rect 16580 12928 16632 12980
rect 17868 12928 17920 12980
rect 19984 12928 20036 12980
rect 20444 12971 20496 12980
rect 20444 12937 20459 12971
rect 20459 12937 20493 12971
rect 20493 12937 20496 12971
rect 21364 12971 21416 12980
rect 20444 12928 20496 12937
rect 21364 12937 21373 12971
rect 21373 12937 21407 12971
rect 21407 12937 21416 12971
rect 21364 12928 21416 12937
rect 22560 12971 22612 12980
rect 22560 12937 22569 12971
rect 22569 12937 22603 12971
rect 22603 12937 22612 12971
rect 22560 12928 22612 12937
rect 25044 12928 25096 12980
rect 25872 12971 25924 12980
rect 25872 12937 25881 12971
rect 25881 12937 25915 12971
rect 25915 12937 25924 12971
rect 25872 12928 25924 12937
rect 27896 12928 27948 12980
rect 16948 12860 17000 12912
rect 16212 12792 16264 12844
rect 16672 12792 16724 12844
rect 17776 12792 17828 12844
rect 15752 12767 15804 12776
rect 15752 12733 15761 12767
rect 15761 12733 15795 12767
rect 15795 12733 15804 12767
rect 15752 12724 15804 12733
rect 16028 12724 16080 12776
rect 17960 12767 18012 12776
rect 17960 12733 17969 12767
rect 17969 12733 18003 12767
rect 18003 12733 18012 12767
rect 19064 12792 19116 12844
rect 20076 12860 20128 12912
rect 20352 12903 20404 12912
rect 20352 12869 20361 12903
rect 20361 12869 20395 12903
rect 20395 12869 20404 12903
rect 20352 12860 20404 12869
rect 23204 12860 23256 12912
rect 19340 12792 19392 12844
rect 20628 12835 20680 12844
rect 20628 12801 20637 12835
rect 20637 12801 20671 12835
rect 20671 12801 20680 12835
rect 20628 12792 20680 12801
rect 21088 12835 21140 12844
rect 18972 12767 19024 12776
rect 17960 12724 18012 12733
rect 18972 12733 18981 12767
rect 18981 12733 19015 12767
rect 19015 12733 19024 12767
rect 18972 12724 19024 12733
rect 19432 12724 19484 12776
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 21824 12835 21876 12844
rect 21824 12801 21833 12835
rect 21833 12801 21867 12835
rect 21867 12801 21876 12835
rect 21824 12792 21876 12801
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 23756 12860 23808 12912
rect 24492 12903 24544 12912
rect 24492 12869 24526 12903
rect 24526 12869 24544 12903
rect 24492 12860 24544 12869
rect 27160 12860 27212 12912
rect 22008 12792 22060 12801
rect 14096 12588 14148 12640
rect 15936 12588 15988 12640
rect 16212 12588 16264 12640
rect 18144 12656 18196 12708
rect 20628 12656 20680 12708
rect 22652 12724 22704 12776
rect 23480 12792 23532 12844
rect 23572 12724 23624 12776
rect 25228 12724 25280 12776
rect 26148 12724 26200 12776
rect 18052 12631 18104 12640
rect 18052 12597 18061 12631
rect 18061 12597 18095 12631
rect 18095 12597 18104 12631
rect 18052 12588 18104 12597
rect 18236 12631 18288 12640
rect 18236 12597 18245 12631
rect 18245 12597 18279 12631
rect 18279 12597 18288 12631
rect 18236 12588 18288 12597
rect 20076 12588 20128 12640
rect 20260 12588 20312 12640
rect 20720 12588 20772 12640
rect 23664 12656 23716 12708
rect 22744 12588 22796 12640
rect 23112 12588 23164 12640
rect 24860 12588 24912 12640
rect 5582 12486 5634 12538
rect 5646 12486 5698 12538
rect 5710 12486 5762 12538
rect 5774 12486 5826 12538
rect 5838 12486 5890 12538
rect 14846 12486 14898 12538
rect 14910 12486 14962 12538
rect 14974 12486 15026 12538
rect 15038 12486 15090 12538
rect 15102 12486 15154 12538
rect 24110 12486 24162 12538
rect 24174 12486 24226 12538
rect 24238 12486 24290 12538
rect 24302 12486 24354 12538
rect 24366 12486 24418 12538
rect 8852 12384 8904 12436
rect 9404 12384 9456 12436
rect 11152 12384 11204 12436
rect 14188 12384 14240 12436
rect 16396 12427 16448 12436
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 18144 12427 18196 12436
rect 18144 12393 18153 12427
rect 18153 12393 18187 12427
rect 18187 12393 18196 12427
rect 18144 12384 18196 12393
rect 18512 12384 18564 12436
rect 6552 12359 6604 12368
rect 6552 12325 6561 12359
rect 6561 12325 6595 12359
rect 6595 12325 6604 12359
rect 6552 12316 6604 12325
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 5264 12180 5316 12232
rect 6644 12248 6696 12300
rect 8208 12180 8260 12232
rect 9128 12248 9180 12300
rect 12072 12248 12124 12300
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 9956 12112 10008 12164
rect 12348 12112 12400 12164
rect 1584 12044 1636 12096
rect 1768 12044 1820 12096
rect 6644 12044 6696 12096
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 7748 12044 7800 12096
rect 9680 12044 9732 12096
rect 11520 12087 11572 12096
rect 11520 12053 11529 12087
rect 11529 12053 11563 12087
rect 11563 12053 11572 12087
rect 11520 12044 11572 12053
rect 12164 12087 12216 12096
rect 12164 12053 12173 12087
rect 12173 12053 12207 12087
rect 12207 12053 12216 12087
rect 12164 12044 12216 12053
rect 12992 12248 13044 12300
rect 12900 12180 12952 12232
rect 14280 12223 14332 12232
rect 12716 12044 12768 12096
rect 12900 12087 12952 12096
rect 12900 12053 12909 12087
rect 12909 12053 12943 12087
rect 12943 12053 12952 12087
rect 13544 12155 13596 12164
rect 13544 12121 13553 12155
rect 13553 12121 13587 12155
rect 13587 12121 13596 12155
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 18052 12248 18104 12300
rect 13544 12112 13596 12121
rect 15844 12180 15896 12232
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 16580 12223 16632 12232
rect 14648 12112 14700 12164
rect 16580 12189 16589 12223
rect 16589 12189 16623 12223
rect 16623 12189 16632 12223
rect 16580 12180 16632 12189
rect 16856 12180 16908 12232
rect 17776 12180 17828 12232
rect 17960 12112 18012 12164
rect 14740 12087 14792 12096
rect 12900 12044 12952 12053
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 17776 12044 17828 12096
rect 17868 12044 17920 12096
rect 19432 12384 19484 12436
rect 19892 12384 19944 12436
rect 20260 12384 20312 12436
rect 23204 12384 23256 12436
rect 23296 12384 23348 12436
rect 25228 12384 25280 12436
rect 27252 12427 27304 12436
rect 27252 12393 27261 12427
rect 27261 12393 27295 12427
rect 27295 12393 27304 12427
rect 27252 12384 27304 12393
rect 24584 12316 24636 12368
rect 19892 12180 19944 12232
rect 20628 12180 20680 12232
rect 21732 12223 21784 12232
rect 20720 12112 20772 12164
rect 21732 12189 21741 12223
rect 21741 12189 21775 12223
rect 21775 12189 21784 12223
rect 21732 12180 21784 12189
rect 19248 12044 19300 12096
rect 20168 12044 20220 12096
rect 20996 12044 21048 12096
rect 22100 12180 22152 12232
rect 22008 12112 22060 12164
rect 22468 12180 22520 12232
rect 22928 12180 22980 12232
rect 23204 12248 23256 12300
rect 22744 12155 22796 12164
rect 22744 12121 22753 12155
rect 22753 12121 22787 12155
rect 22787 12121 22796 12155
rect 22744 12112 22796 12121
rect 22560 12044 22612 12096
rect 22928 12044 22980 12096
rect 23204 12112 23256 12164
rect 25044 12248 25096 12300
rect 28356 12291 28408 12300
rect 28356 12257 28365 12291
rect 28365 12257 28399 12291
rect 28399 12257 28408 12291
rect 28356 12248 28408 12257
rect 23756 12180 23808 12232
rect 24676 12223 24728 12232
rect 24676 12189 24685 12223
rect 24685 12189 24719 12223
rect 24719 12189 24728 12223
rect 24676 12180 24728 12189
rect 25688 12223 25740 12232
rect 25688 12189 25697 12223
rect 25697 12189 25731 12223
rect 25731 12189 25740 12223
rect 25688 12180 25740 12189
rect 27068 12223 27120 12232
rect 27068 12189 27077 12223
rect 27077 12189 27111 12223
rect 27111 12189 27120 12223
rect 27068 12180 27120 12189
rect 23664 12112 23716 12164
rect 24492 12112 24544 12164
rect 24768 12112 24820 12164
rect 25228 12155 25280 12164
rect 25228 12121 25237 12155
rect 25237 12121 25271 12155
rect 25271 12121 25280 12155
rect 25228 12112 25280 12121
rect 23572 12044 23624 12096
rect 23848 12087 23900 12096
rect 23848 12053 23857 12087
rect 23857 12053 23891 12087
rect 23891 12053 23900 12087
rect 23848 12044 23900 12053
rect 24952 12044 25004 12096
rect 26148 12044 26200 12096
rect 10214 11942 10266 11994
rect 10278 11942 10330 11994
rect 10342 11942 10394 11994
rect 10406 11942 10458 11994
rect 10470 11942 10522 11994
rect 19478 11942 19530 11994
rect 19542 11942 19594 11994
rect 19606 11942 19658 11994
rect 19670 11942 19722 11994
rect 19734 11942 19786 11994
rect 6000 11883 6052 11892
rect 6000 11849 6009 11883
rect 6009 11849 6043 11883
rect 6043 11849 6052 11883
rect 6000 11840 6052 11849
rect 7932 11883 7984 11892
rect 7932 11849 7941 11883
rect 7941 11849 7975 11883
rect 7975 11849 7984 11883
rect 7932 11840 7984 11849
rect 8576 11840 8628 11892
rect 10876 11840 10928 11892
rect 11244 11840 11296 11892
rect 12072 11840 12124 11892
rect 15660 11883 15712 11892
rect 6644 11747 6696 11756
rect 6644 11713 6653 11747
rect 6653 11713 6687 11747
rect 6687 11713 6696 11747
rect 6644 11704 6696 11713
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 8852 11704 8904 11756
rect 9496 11704 9548 11756
rect 12532 11704 12584 11756
rect 7288 11636 7340 11688
rect 9128 11636 9180 11688
rect 9312 11636 9364 11688
rect 11152 11636 11204 11688
rect 12900 11636 12952 11688
rect 14188 11704 14240 11756
rect 9220 11611 9272 11620
rect 9220 11577 9229 11611
rect 9229 11577 9263 11611
rect 9263 11577 9272 11611
rect 9220 11568 9272 11577
rect 13728 11636 13780 11688
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 16396 11840 16448 11892
rect 16672 11883 16724 11892
rect 16672 11849 16681 11883
rect 16681 11849 16715 11883
rect 16715 11849 16724 11883
rect 16672 11840 16724 11849
rect 19248 11883 19300 11892
rect 19248 11849 19257 11883
rect 19257 11849 19291 11883
rect 19291 11849 19300 11883
rect 19248 11840 19300 11849
rect 16580 11772 16632 11824
rect 14556 11747 14608 11756
rect 14556 11713 14590 11747
rect 14590 11713 14608 11747
rect 16120 11747 16172 11756
rect 14556 11704 14608 11713
rect 16120 11713 16129 11747
rect 16129 11713 16163 11747
rect 16163 11713 16172 11747
rect 16120 11704 16172 11713
rect 16212 11704 16264 11756
rect 17868 11704 17920 11756
rect 18236 11772 18288 11824
rect 19064 11704 19116 11756
rect 20628 11840 20680 11892
rect 23848 11840 23900 11892
rect 24860 11840 24912 11892
rect 19800 11704 19852 11756
rect 24768 11772 24820 11824
rect 20996 11747 21048 11756
rect 20996 11713 21005 11747
rect 21005 11713 21039 11747
rect 21039 11713 21048 11747
rect 20996 11704 21048 11713
rect 21732 11704 21784 11756
rect 22376 11704 22428 11756
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22836 11747 22888 11756
rect 22560 11704 22612 11713
rect 22836 11713 22845 11747
rect 22845 11713 22879 11747
rect 22879 11713 22888 11747
rect 22836 11704 22888 11713
rect 23020 11747 23072 11756
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 23756 11704 23808 11756
rect 24032 11704 24084 11756
rect 17132 11679 17184 11688
rect 7380 11500 7432 11552
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 11244 11500 11296 11552
rect 13452 11568 13504 11620
rect 17132 11645 17141 11679
rect 17141 11645 17175 11679
rect 17175 11645 17184 11679
rect 17132 11636 17184 11645
rect 17408 11679 17460 11688
rect 17408 11645 17417 11679
rect 17417 11645 17451 11679
rect 17451 11645 17460 11679
rect 17408 11636 17460 11645
rect 17776 11636 17828 11688
rect 20536 11636 20588 11688
rect 23388 11636 23440 11688
rect 23480 11636 23532 11688
rect 25504 11747 25556 11756
rect 25504 11713 25513 11747
rect 25513 11713 25547 11747
rect 25547 11713 25556 11747
rect 25504 11704 25556 11713
rect 25688 11636 25740 11688
rect 13360 11500 13412 11552
rect 16212 11568 16264 11620
rect 18972 11568 19024 11620
rect 14280 11500 14332 11552
rect 18788 11543 18840 11552
rect 18788 11509 18797 11543
rect 18797 11509 18831 11543
rect 18831 11509 18840 11543
rect 18788 11500 18840 11509
rect 19524 11568 19576 11620
rect 22008 11568 22060 11620
rect 20812 11543 20864 11552
rect 20812 11509 20821 11543
rect 20821 11509 20855 11543
rect 20855 11509 20864 11543
rect 20812 11500 20864 11509
rect 22376 11543 22428 11552
rect 22376 11509 22385 11543
rect 22385 11509 22419 11543
rect 22419 11509 22428 11543
rect 22376 11500 22428 11509
rect 22652 11611 22704 11620
rect 22652 11577 22661 11611
rect 22661 11577 22695 11611
rect 22695 11577 22704 11611
rect 22652 11568 22704 11577
rect 23204 11568 23256 11620
rect 24032 11500 24084 11552
rect 24952 11500 25004 11552
rect 5582 11398 5634 11450
rect 5646 11398 5698 11450
rect 5710 11398 5762 11450
rect 5774 11398 5826 11450
rect 5838 11398 5890 11450
rect 14846 11398 14898 11450
rect 14910 11398 14962 11450
rect 14974 11398 15026 11450
rect 15038 11398 15090 11450
rect 15102 11398 15154 11450
rect 24110 11398 24162 11450
rect 24174 11398 24226 11450
rect 24238 11398 24290 11450
rect 24302 11398 24354 11450
rect 24366 11398 24418 11450
rect 7288 11296 7340 11348
rect 8576 11296 8628 11348
rect 10140 11296 10192 11348
rect 12164 11296 12216 11348
rect 12716 11296 12768 11348
rect 13452 11296 13504 11348
rect 14464 11296 14516 11348
rect 14556 11296 14608 11348
rect 17224 11339 17276 11348
rect 17224 11305 17233 11339
rect 17233 11305 17267 11339
rect 17267 11305 17276 11339
rect 17224 11296 17276 11305
rect 18604 11296 18656 11348
rect 22008 11339 22060 11348
rect 9496 11271 9548 11280
rect 9496 11237 9505 11271
rect 9505 11237 9539 11271
rect 9539 11237 9548 11271
rect 9496 11228 9548 11237
rect 8300 11160 8352 11212
rect 13176 11228 13228 11280
rect 16212 11271 16264 11280
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 7380 11135 7432 11144
rect 7380 11101 7398 11135
rect 7398 11101 7432 11135
rect 8024 11135 8076 11144
rect 7380 11092 7432 11101
rect 8024 11101 8033 11135
rect 8033 11101 8067 11135
rect 8067 11101 8076 11135
rect 8024 11092 8076 11101
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 12440 11160 12492 11212
rect 10876 11135 10928 11144
rect 8760 11024 8812 11076
rect 9864 11024 9916 11076
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 11888 11092 11940 11144
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 13360 11092 13412 11144
rect 14188 11135 14240 11144
rect 14188 11101 14197 11135
rect 14197 11101 14231 11135
rect 14231 11101 14240 11135
rect 14188 11092 14240 11101
rect 14280 11092 14332 11144
rect 14740 11160 14792 11212
rect 16212 11237 16221 11271
rect 16221 11237 16255 11271
rect 16255 11237 16264 11271
rect 16212 11228 16264 11237
rect 17132 11228 17184 11280
rect 19248 11228 19300 11280
rect 20076 11228 20128 11280
rect 17868 11160 17920 11212
rect 15292 11135 15344 11144
rect 13268 11024 13320 11076
rect 13728 11024 13780 11076
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 15660 11135 15712 11144
rect 15200 11024 15252 11076
rect 15660 11101 15669 11135
rect 15669 11101 15703 11135
rect 15703 11101 15712 11135
rect 15660 11092 15712 11101
rect 15752 11135 15804 11144
rect 15752 11101 15766 11135
rect 15766 11101 15800 11135
rect 15800 11101 15804 11135
rect 18236 11135 18288 11144
rect 15752 11092 15804 11101
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 20168 11160 20220 11212
rect 19984 11092 20036 11144
rect 22008 11305 22017 11339
rect 22017 11305 22051 11339
rect 22051 11305 22060 11339
rect 22008 11296 22060 11305
rect 22284 11339 22336 11348
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 22836 11296 22888 11348
rect 23204 11228 23256 11280
rect 23848 11296 23900 11348
rect 24676 11339 24728 11348
rect 24676 11305 24685 11339
rect 24685 11305 24719 11339
rect 24719 11305 24728 11339
rect 24676 11296 24728 11305
rect 25504 11296 25556 11348
rect 22468 11160 22520 11212
rect 23388 11203 23440 11212
rect 23388 11169 23397 11203
rect 23397 11169 23431 11203
rect 23431 11169 23440 11203
rect 23388 11160 23440 11169
rect 22652 11135 22704 11144
rect 11244 10956 11296 11008
rect 13912 10956 13964 11008
rect 14648 10956 14700 11008
rect 15108 10956 15160 11008
rect 17408 11067 17460 11076
rect 17408 11033 17417 11067
rect 17417 11033 17451 11067
rect 17451 11033 17460 11067
rect 17408 11024 17460 11033
rect 17960 11024 18012 11076
rect 18512 11024 18564 11076
rect 18604 11024 18656 11076
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 20720 11024 20772 11076
rect 20812 11024 20864 11076
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 23112 11092 23164 11144
rect 23296 11092 23348 11144
rect 24032 11228 24084 11280
rect 24676 11160 24728 11212
rect 22284 11024 22336 11076
rect 24032 11024 24084 11076
rect 20260 10956 20312 11008
rect 25228 11092 25280 11144
rect 28356 11135 28408 11144
rect 28356 11101 28365 11135
rect 28365 11101 28399 11135
rect 28399 11101 28408 11135
rect 28356 11092 28408 11101
rect 24492 11024 24544 11076
rect 25320 11067 25372 11076
rect 25320 11033 25329 11067
rect 25329 11033 25363 11067
rect 25363 11033 25372 11067
rect 25320 11024 25372 11033
rect 26148 11024 26200 11076
rect 24860 10956 24912 11008
rect 10214 10854 10266 10906
rect 10278 10854 10330 10906
rect 10342 10854 10394 10906
rect 10406 10854 10458 10906
rect 10470 10854 10522 10906
rect 19478 10854 19530 10906
rect 19542 10854 19594 10906
rect 19606 10854 19658 10906
rect 19670 10854 19722 10906
rect 19734 10854 19786 10906
rect 8852 10752 8904 10804
rect 10140 10752 10192 10804
rect 8300 10684 8352 10736
rect 10876 10684 10928 10736
rect 16304 10752 16356 10804
rect 16856 10795 16908 10804
rect 16856 10761 16865 10795
rect 16865 10761 16899 10795
rect 16899 10761 16908 10795
rect 16856 10752 16908 10761
rect 23388 10752 23440 10804
rect 8576 10616 8628 10668
rect 10048 10616 10100 10668
rect 9864 10548 9916 10600
rect 12992 10684 13044 10736
rect 13544 10684 13596 10736
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 12532 10523 12584 10532
rect 9772 10412 9824 10464
rect 11428 10412 11480 10464
rect 12532 10489 12541 10523
rect 12541 10489 12575 10523
rect 12575 10489 12584 10523
rect 12532 10480 12584 10489
rect 12716 10412 12768 10464
rect 13360 10591 13412 10600
rect 13360 10557 13369 10591
rect 13369 10557 13403 10591
rect 13403 10557 13412 10591
rect 13360 10548 13412 10557
rect 13268 10480 13320 10532
rect 14280 10616 14332 10668
rect 15476 10684 15528 10736
rect 14740 10616 14792 10668
rect 15384 10412 15436 10464
rect 15752 10591 15804 10600
rect 15752 10557 15761 10591
rect 15761 10557 15795 10591
rect 15795 10557 15804 10591
rect 15752 10548 15804 10557
rect 18604 10684 18656 10736
rect 22376 10684 22428 10736
rect 17684 10659 17736 10668
rect 15568 10480 15620 10532
rect 17684 10625 17693 10659
rect 17693 10625 17727 10659
rect 17727 10625 17736 10659
rect 17684 10616 17736 10625
rect 19064 10659 19116 10668
rect 19064 10625 19082 10659
rect 19082 10625 19116 10659
rect 19064 10616 19116 10625
rect 20628 10616 20680 10668
rect 24492 10752 24544 10804
rect 24676 10752 24728 10804
rect 24952 10752 25004 10804
rect 26240 10752 26292 10804
rect 25228 10684 25280 10736
rect 25320 10684 25372 10736
rect 19432 10548 19484 10600
rect 19892 10548 19944 10600
rect 18328 10480 18380 10532
rect 17316 10455 17368 10464
rect 17316 10421 17325 10455
rect 17325 10421 17359 10455
rect 17359 10421 17368 10455
rect 17316 10412 17368 10421
rect 17960 10455 18012 10464
rect 17960 10421 17969 10455
rect 17969 10421 18003 10455
rect 18003 10421 18012 10455
rect 17960 10412 18012 10421
rect 18052 10412 18104 10464
rect 18972 10412 19024 10464
rect 24584 10616 24636 10668
rect 25780 10616 25832 10668
rect 26792 10616 26844 10668
rect 21272 10412 21324 10464
rect 22100 10412 22152 10464
rect 23296 10412 23348 10464
rect 26240 10412 26292 10464
rect 27344 10412 27396 10464
rect 5582 10310 5634 10362
rect 5646 10310 5698 10362
rect 5710 10310 5762 10362
rect 5774 10310 5826 10362
rect 5838 10310 5890 10362
rect 14846 10310 14898 10362
rect 14910 10310 14962 10362
rect 14974 10310 15026 10362
rect 15038 10310 15090 10362
rect 15102 10310 15154 10362
rect 24110 10310 24162 10362
rect 24174 10310 24226 10362
rect 24238 10310 24290 10362
rect 24302 10310 24354 10362
rect 24366 10310 24418 10362
rect 9680 10208 9732 10260
rect 13084 10208 13136 10260
rect 12716 10140 12768 10192
rect 14188 10208 14240 10260
rect 15292 10208 15344 10260
rect 15568 10251 15620 10260
rect 15568 10217 15577 10251
rect 15577 10217 15611 10251
rect 15611 10217 15620 10251
rect 15568 10208 15620 10217
rect 15752 10208 15804 10260
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 19064 10208 19116 10260
rect 19984 10208 20036 10260
rect 20628 10251 20680 10260
rect 20628 10217 20637 10251
rect 20637 10217 20671 10251
rect 20671 10217 20680 10251
rect 20628 10208 20680 10217
rect 25780 10251 25832 10260
rect 25780 10217 25789 10251
rect 25789 10217 25823 10251
rect 25823 10217 25832 10251
rect 25780 10208 25832 10217
rect 13268 10140 13320 10192
rect 8300 10072 8352 10124
rect 8944 10072 8996 10124
rect 9312 10115 9364 10124
rect 9312 10081 9321 10115
rect 9321 10081 9355 10115
rect 9355 10081 9364 10115
rect 9312 10072 9364 10081
rect 11152 10115 11204 10124
rect 11152 10081 11161 10115
rect 11161 10081 11195 10115
rect 11195 10081 11204 10115
rect 11152 10072 11204 10081
rect 12440 10072 12492 10124
rect 14004 10072 14056 10124
rect 9220 10004 9272 10056
rect 11428 10047 11480 10056
rect 11428 10013 11462 10047
rect 11462 10013 11480 10047
rect 11428 10004 11480 10013
rect 1584 9936 1636 9988
rect 9588 9979 9640 9988
rect 9588 9945 9622 9979
rect 9622 9945 9640 9979
rect 9588 9936 9640 9945
rect 10692 9911 10744 9920
rect 10692 9877 10701 9911
rect 10701 9877 10735 9911
rect 10735 9877 10744 9911
rect 11796 9936 11848 9988
rect 13084 10004 13136 10056
rect 13820 10004 13872 10056
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 14280 10047 14332 10056
rect 14280 10013 14290 10047
rect 14290 10013 14324 10047
rect 14324 10013 14332 10047
rect 16212 10072 16264 10124
rect 19432 10140 19484 10192
rect 18236 10072 18288 10124
rect 18788 10072 18840 10124
rect 21272 10140 21324 10192
rect 23572 10140 23624 10192
rect 20168 10115 20220 10124
rect 20168 10081 20177 10115
rect 20177 10081 20211 10115
rect 20211 10081 20220 10115
rect 20168 10072 20220 10081
rect 14280 10004 14332 10013
rect 15384 10047 15436 10056
rect 10692 9868 10744 9877
rect 13452 9868 13504 9920
rect 13912 9936 13964 9988
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 16856 10004 16908 10056
rect 17316 10004 17368 10056
rect 19984 10047 20036 10056
rect 19984 10013 19993 10047
rect 19993 10013 20027 10047
rect 20027 10013 20036 10047
rect 23296 10072 23348 10124
rect 24676 10072 24728 10124
rect 26792 10140 26844 10192
rect 19984 10004 20036 10013
rect 20720 10004 20772 10056
rect 17960 9936 18012 9988
rect 18420 9936 18472 9988
rect 23940 10004 23992 10056
rect 25136 10004 25188 10056
rect 25320 10047 25372 10056
rect 25320 10013 25329 10047
rect 25329 10013 25363 10047
rect 25363 10013 25372 10047
rect 25320 10004 25372 10013
rect 27344 10004 27396 10056
rect 23572 9979 23624 9988
rect 23572 9945 23581 9979
rect 23581 9945 23615 9979
rect 23615 9945 23624 9979
rect 23572 9936 23624 9945
rect 24032 9936 24084 9988
rect 24860 9979 24912 9988
rect 24860 9945 24869 9979
rect 24869 9945 24903 9979
rect 24903 9945 24912 9979
rect 24860 9936 24912 9945
rect 14648 9868 14700 9920
rect 18052 9911 18104 9920
rect 18052 9877 18061 9911
rect 18061 9877 18095 9911
rect 18095 9877 18104 9911
rect 18052 9868 18104 9877
rect 19892 9868 19944 9920
rect 21180 9868 21232 9920
rect 22192 9868 22244 9920
rect 22468 9911 22520 9920
rect 22468 9877 22477 9911
rect 22477 9877 22511 9911
rect 22511 9877 22520 9911
rect 22468 9868 22520 9877
rect 23480 9868 23532 9920
rect 23848 9868 23900 9920
rect 25504 9911 25556 9920
rect 25504 9877 25513 9911
rect 25513 9877 25547 9911
rect 25547 9877 25556 9911
rect 25504 9868 25556 9877
rect 26516 9868 26568 9920
rect 28080 9868 28132 9920
rect 10214 9766 10266 9818
rect 10278 9766 10330 9818
rect 10342 9766 10394 9818
rect 10406 9766 10458 9818
rect 10470 9766 10522 9818
rect 19478 9766 19530 9818
rect 19542 9766 19594 9818
rect 19606 9766 19658 9818
rect 19670 9766 19722 9818
rect 19734 9766 19786 9818
rect 8576 9707 8628 9716
rect 8576 9673 8585 9707
rect 8585 9673 8619 9707
rect 8619 9673 8628 9707
rect 8576 9664 8628 9673
rect 9588 9707 9640 9716
rect 9588 9673 9597 9707
rect 9597 9673 9631 9707
rect 9631 9673 9640 9707
rect 9588 9664 9640 9673
rect 10048 9707 10100 9716
rect 10048 9673 10057 9707
rect 10057 9673 10091 9707
rect 10091 9673 10100 9707
rect 10048 9664 10100 9673
rect 10692 9664 10744 9716
rect 11704 9664 11756 9716
rect 11980 9664 12032 9716
rect 14280 9707 14332 9716
rect 14280 9673 14289 9707
rect 14289 9673 14323 9707
rect 14323 9673 14332 9707
rect 14280 9664 14332 9673
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 11244 9596 11296 9648
rect 12440 9596 12492 9648
rect 12716 9596 12768 9648
rect 13176 9639 13228 9648
rect 13176 9605 13210 9639
rect 13210 9605 13228 9639
rect 13176 9596 13228 9605
rect 13268 9596 13320 9648
rect 13452 9596 13504 9648
rect 11796 9528 11848 9580
rect 15568 9596 15620 9648
rect 15752 9596 15804 9648
rect 17960 9596 18012 9648
rect 22468 9664 22520 9716
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 15200 9503 15252 9512
rect 9220 9367 9272 9376
rect 9220 9333 9229 9367
rect 9229 9333 9263 9367
rect 9263 9333 9272 9367
rect 10784 9392 10836 9444
rect 12716 9392 12768 9444
rect 15200 9469 15209 9503
rect 15209 9469 15243 9503
rect 15243 9469 15252 9503
rect 15200 9460 15252 9469
rect 16212 9571 16264 9580
rect 16212 9537 16221 9571
rect 16221 9537 16255 9571
rect 16255 9537 16264 9571
rect 16212 9528 16264 9537
rect 17040 9528 17092 9580
rect 18420 9571 18472 9580
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 18604 9571 18656 9580
rect 18604 9537 18613 9571
rect 18613 9537 18647 9571
rect 18647 9537 18656 9571
rect 18604 9528 18656 9537
rect 20076 9596 20128 9648
rect 19340 9528 19392 9580
rect 15476 9392 15528 9444
rect 17868 9435 17920 9444
rect 17868 9401 17877 9435
rect 17877 9401 17911 9435
rect 17911 9401 17920 9435
rect 17868 9392 17920 9401
rect 19892 9528 19944 9580
rect 21180 9571 21232 9580
rect 21180 9537 21198 9571
rect 21198 9537 21232 9571
rect 21180 9528 21232 9537
rect 22100 9528 22152 9580
rect 19708 9503 19760 9512
rect 19708 9469 19717 9503
rect 19717 9469 19751 9503
rect 19751 9469 19760 9503
rect 19708 9460 19760 9469
rect 20168 9460 20220 9512
rect 22284 9528 22336 9580
rect 22376 9503 22428 9512
rect 22376 9469 22385 9503
rect 22385 9469 22419 9503
rect 22419 9469 22428 9503
rect 22376 9460 22428 9469
rect 9220 9324 9272 9333
rect 13544 9324 13596 9376
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 16672 9324 16724 9333
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 24032 9528 24084 9580
rect 25504 9596 25556 9648
rect 28264 9571 28316 9580
rect 28264 9537 28273 9571
rect 28273 9537 28307 9571
rect 28307 9537 28316 9571
rect 28264 9528 28316 9537
rect 23480 9435 23532 9444
rect 23480 9401 23489 9435
rect 23489 9401 23523 9435
rect 23523 9401 23532 9435
rect 23480 9392 23532 9401
rect 24676 9324 24728 9376
rect 26516 9435 26568 9444
rect 26516 9401 26525 9435
rect 26525 9401 26559 9435
rect 26559 9401 26568 9435
rect 26516 9392 26568 9401
rect 5582 9222 5634 9274
rect 5646 9222 5698 9274
rect 5710 9222 5762 9274
rect 5774 9222 5826 9274
rect 5838 9222 5890 9274
rect 14846 9222 14898 9274
rect 14910 9222 14962 9274
rect 14974 9222 15026 9274
rect 15038 9222 15090 9274
rect 15102 9222 15154 9274
rect 24110 9222 24162 9274
rect 24174 9222 24226 9274
rect 24238 9222 24290 9274
rect 24302 9222 24354 9274
rect 24366 9222 24418 9274
rect 14556 9120 14608 9172
rect 15200 9120 15252 9172
rect 17040 9163 17092 9172
rect 17040 9129 17049 9163
rect 17049 9129 17083 9163
rect 17083 9129 17092 9163
rect 17040 9120 17092 9129
rect 17316 9120 17368 9172
rect 8944 9027 8996 9036
rect 8944 8993 8953 9027
rect 8953 8993 8987 9027
rect 8987 8993 8996 9027
rect 8944 8984 8996 8993
rect 12624 9052 12676 9104
rect 12900 9052 12952 9104
rect 11244 9027 11296 9036
rect 11244 8993 11253 9027
rect 11253 8993 11287 9027
rect 11287 8993 11296 9027
rect 11244 8984 11296 8993
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 13820 8984 13872 9036
rect 18604 9052 18656 9104
rect 20812 9052 20864 9104
rect 22376 9052 22428 9104
rect 8392 8959 8444 8968
rect 8392 8925 8401 8959
rect 8401 8925 8435 8959
rect 8435 8925 8444 8959
rect 8392 8916 8444 8925
rect 11612 8916 11664 8968
rect 11888 8916 11940 8968
rect 11980 8916 12032 8968
rect 13452 8916 13504 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 19340 8984 19392 9036
rect 19708 9027 19760 9036
rect 19708 8993 19717 9027
rect 19717 8993 19751 9027
rect 19751 8993 19760 9027
rect 19708 8984 19760 8993
rect 13544 8916 13596 8925
rect 13084 8848 13136 8900
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 15844 8916 15896 8968
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 14372 8891 14424 8900
rect 14372 8857 14381 8891
rect 14381 8857 14415 8891
rect 14415 8857 14424 8891
rect 14372 8848 14424 8857
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 12532 8823 12584 8832
rect 12532 8789 12541 8823
rect 12541 8789 12575 8823
rect 12575 8789 12584 8823
rect 12532 8780 12584 8789
rect 14924 8780 14976 8832
rect 17500 8848 17552 8900
rect 20352 8916 20404 8968
rect 21364 8916 21416 8968
rect 23572 9120 23624 9172
rect 25320 9163 25372 9172
rect 25320 9129 25329 9163
rect 25329 9129 25363 9163
rect 25363 9129 25372 9163
rect 25320 9120 25372 9129
rect 26516 9052 26568 9104
rect 23480 8984 23532 9036
rect 24860 8984 24912 9036
rect 25136 8984 25188 9036
rect 24768 8916 24820 8968
rect 25596 8916 25648 8968
rect 18328 8848 18380 8900
rect 20812 8891 20864 8900
rect 17868 8780 17920 8832
rect 18144 8780 18196 8832
rect 19984 8823 20036 8832
rect 19984 8789 19993 8823
rect 19993 8789 20027 8823
rect 20027 8789 20036 8823
rect 19984 8780 20036 8789
rect 20812 8857 20821 8891
rect 20821 8857 20855 8891
rect 20855 8857 20864 8891
rect 20812 8848 20864 8857
rect 21824 8848 21876 8900
rect 22100 8848 22152 8900
rect 24676 8848 24728 8900
rect 20996 8823 21048 8832
rect 20996 8789 21005 8823
rect 21005 8789 21039 8823
rect 21039 8789 21048 8823
rect 20996 8780 21048 8789
rect 21088 8780 21140 8832
rect 22376 8780 22428 8832
rect 25780 8823 25832 8832
rect 25780 8789 25789 8823
rect 25789 8789 25823 8823
rect 25823 8789 25832 8823
rect 25780 8780 25832 8789
rect 10214 8678 10266 8730
rect 10278 8678 10330 8730
rect 10342 8678 10394 8730
rect 10406 8678 10458 8730
rect 10470 8678 10522 8730
rect 19478 8678 19530 8730
rect 19542 8678 19594 8730
rect 19606 8678 19658 8730
rect 19670 8678 19722 8730
rect 19734 8678 19786 8730
rect 8392 8576 8444 8628
rect 13084 8576 13136 8628
rect 13636 8619 13688 8628
rect 13636 8585 13645 8619
rect 13645 8585 13679 8619
rect 13679 8585 13688 8619
rect 13636 8576 13688 8585
rect 14188 8576 14240 8628
rect 14372 8576 14424 8628
rect 14556 8576 14608 8628
rect 16856 8619 16908 8628
rect 1492 8440 1544 8492
rect 10600 8440 10652 8492
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 11520 8440 11572 8492
rect 12900 8508 12952 8560
rect 16856 8585 16865 8619
rect 16865 8585 16899 8619
rect 16899 8585 16908 8619
rect 16856 8576 16908 8585
rect 17316 8619 17368 8628
rect 17316 8585 17325 8619
rect 17325 8585 17359 8619
rect 17359 8585 17368 8619
rect 17316 8576 17368 8585
rect 18512 8619 18564 8628
rect 18512 8585 18521 8619
rect 18521 8585 18555 8619
rect 18555 8585 18564 8619
rect 18512 8576 18564 8585
rect 21088 8576 21140 8628
rect 21824 8619 21876 8628
rect 21824 8585 21833 8619
rect 21833 8585 21867 8619
rect 21867 8585 21876 8619
rect 21824 8576 21876 8585
rect 24032 8619 24084 8628
rect 24032 8585 24041 8619
rect 24041 8585 24075 8619
rect 24075 8585 24084 8619
rect 24032 8576 24084 8585
rect 11888 8483 11940 8492
rect 11888 8449 11922 8483
rect 11922 8449 11940 8483
rect 11888 8440 11940 8449
rect 9864 8372 9916 8424
rect 11244 8372 11296 8424
rect 13360 8372 13412 8424
rect 15476 8551 15528 8560
rect 15476 8517 15485 8551
rect 15485 8517 15519 8551
rect 15519 8517 15528 8551
rect 15476 8508 15528 8517
rect 14280 8440 14332 8492
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 14924 8483 14976 8492
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 18236 8508 18288 8560
rect 19984 8508 20036 8560
rect 22284 8508 22336 8560
rect 23296 8508 23348 8560
rect 1584 8347 1636 8356
rect 1584 8313 1593 8347
rect 1593 8313 1627 8347
rect 1627 8313 1636 8347
rect 1584 8304 1636 8313
rect 13176 8304 13228 8356
rect 10140 8236 10192 8288
rect 13268 8279 13320 8288
rect 13268 8245 13277 8279
rect 13277 8245 13311 8279
rect 13311 8245 13320 8279
rect 13268 8236 13320 8245
rect 14464 8304 14516 8356
rect 17132 8440 17184 8492
rect 18052 8483 18104 8492
rect 15844 8372 15896 8424
rect 16028 8372 16080 8424
rect 16672 8372 16724 8424
rect 18052 8449 18061 8483
rect 18061 8449 18095 8483
rect 18095 8449 18104 8483
rect 18052 8440 18104 8449
rect 19064 8440 19116 8492
rect 19340 8440 19392 8492
rect 19800 8483 19852 8492
rect 19800 8449 19809 8483
rect 19809 8449 19843 8483
rect 19843 8449 19852 8483
rect 19800 8440 19852 8449
rect 20996 8440 21048 8492
rect 22192 8440 22244 8492
rect 23848 8483 23900 8492
rect 23848 8449 23857 8483
rect 23857 8449 23891 8483
rect 23891 8449 23900 8483
rect 23848 8440 23900 8449
rect 24952 8440 25004 8492
rect 28356 8483 28408 8492
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 18144 8415 18196 8424
rect 16764 8304 16816 8356
rect 18144 8381 18153 8415
rect 18153 8381 18187 8415
rect 18187 8381 18196 8415
rect 18144 8372 18196 8381
rect 22744 8372 22796 8424
rect 24584 8415 24636 8424
rect 18420 8304 18472 8356
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 24584 8372 24636 8381
rect 25136 8372 25188 8424
rect 26516 8304 26568 8356
rect 18328 8279 18380 8288
rect 18328 8245 18337 8279
rect 18337 8245 18371 8279
rect 18371 8245 18380 8279
rect 18328 8236 18380 8245
rect 19340 8236 19392 8288
rect 20444 8279 20496 8288
rect 20444 8245 20453 8279
rect 20453 8245 20487 8279
rect 20487 8245 20496 8279
rect 20444 8236 20496 8245
rect 22836 8279 22888 8288
rect 22836 8245 22845 8279
rect 22845 8245 22879 8279
rect 22879 8245 22888 8279
rect 22836 8236 22888 8245
rect 28172 8279 28224 8288
rect 28172 8245 28181 8279
rect 28181 8245 28215 8279
rect 28215 8245 28224 8279
rect 28172 8236 28224 8245
rect 5582 8134 5634 8186
rect 5646 8134 5698 8186
rect 5710 8134 5762 8186
rect 5774 8134 5826 8186
rect 5838 8134 5890 8186
rect 14846 8134 14898 8186
rect 14910 8134 14962 8186
rect 14974 8134 15026 8186
rect 15038 8134 15090 8186
rect 15102 8134 15154 8186
rect 24110 8134 24162 8186
rect 24174 8134 24226 8186
rect 24238 8134 24290 8186
rect 24302 8134 24354 8186
rect 24366 8134 24418 8186
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 13452 8075 13504 8084
rect 13452 8041 13461 8075
rect 13461 8041 13495 8075
rect 13495 8041 13504 8075
rect 13452 8032 13504 8041
rect 13820 8032 13872 8084
rect 14556 8032 14608 8084
rect 19800 8032 19852 8084
rect 11520 8007 11572 8016
rect 11520 7973 11529 8007
rect 11529 7973 11563 8007
rect 11563 7973 11572 8007
rect 11520 7964 11572 7973
rect 11980 8007 12032 8016
rect 11980 7973 11989 8007
rect 11989 7973 12023 8007
rect 12023 7973 12032 8007
rect 11980 7964 12032 7973
rect 18328 7964 18380 8016
rect 28172 8032 28224 8084
rect 21364 7964 21416 8016
rect 24032 8007 24084 8016
rect 24032 7973 24041 8007
rect 24041 7973 24075 8007
rect 24075 7973 24084 8007
rect 24032 7964 24084 7973
rect 24584 7964 24636 8016
rect 10048 7828 10100 7880
rect 12532 7896 12584 7948
rect 12256 7828 12308 7880
rect 19984 7896 20036 7948
rect 20352 7939 20404 7948
rect 20352 7905 20361 7939
rect 20361 7905 20395 7939
rect 20395 7905 20404 7939
rect 20352 7896 20404 7905
rect 22100 7896 22152 7948
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 15108 7828 15160 7880
rect 17776 7828 17828 7880
rect 19340 7828 19392 7880
rect 20444 7828 20496 7880
rect 24676 7828 24728 7880
rect 26516 7871 26568 7880
rect 26516 7837 26525 7871
rect 26525 7837 26559 7871
rect 26559 7837 26568 7871
rect 26516 7828 26568 7837
rect 11520 7760 11572 7812
rect 14280 7760 14332 7812
rect 16212 7803 16264 7812
rect 16212 7769 16230 7803
rect 16230 7769 16264 7803
rect 16212 7760 16264 7769
rect 17040 7760 17092 7812
rect 14832 7735 14884 7744
rect 14832 7701 14841 7735
rect 14841 7701 14875 7735
rect 14875 7701 14884 7735
rect 14832 7692 14884 7701
rect 17684 7692 17736 7744
rect 18788 7692 18840 7744
rect 19892 7760 19944 7812
rect 22100 7760 22152 7812
rect 25412 7692 25464 7744
rect 10214 7590 10266 7642
rect 10278 7590 10330 7642
rect 10342 7590 10394 7642
rect 10406 7590 10458 7642
rect 10470 7590 10522 7642
rect 19478 7590 19530 7642
rect 19542 7590 19594 7642
rect 19606 7590 19658 7642
rect 19670 7590 19722 7642
rect 19734 7590 19786 7642
rect 10048 7531 10100 7540
rect 10048 7497 10057 7531
rect 10057 7497 10091 7531
rect 10091 7497 10100 7531
rect 10048 7488 10100 7497
rect 11612 7488 11664 7540
rect 15108 7531 15160 7540
rect 9864 7420 9916 7472
rect 10140 7352 10192 7404
rect 15108 7497 15117 7531
rect 15117 7497 15151 7531
rect 15151 7497 15160 7531
rect 15108 7488 15160 7497
rect 16212 7488 16264 7540
rect 17040 7488 17092 7540
rect 17132 7488 17184 7540
rect 17684 7531 17736 7540
rect 17684 7497 17693 7531
rect 17693 7497 17727 7531
rect 17727 7497 17736 7531
rect 17684 7488 17736 7497
rect 22100 7531 22152 7540
rect 22100 7497 22109 7531
rect 22109 7497 22143 7531
rect 22143 7497 22152 7531
rect 22100 7488 22152 7497
rect 24032 7488 24084 7540
rect 24952 7531 25004 7540
rect 24952 7497 24961 7531
rect 24961 7497 24995 7531
rect 24995 7497 25004 7531
rect 24952 7488 25004 7497
rect 25412 7531 25464 7540
rect 25412 7497 25421 7531
rect 25421 7497 25455 7531
rect 25455 7497 25464 7531
rect 25412 7488 25464 7497
rect 25780 7488 25832 7540
rect 14832 7420 14884 7472
rect 12256 7395 12308 7404
rect 12256 7361 12265 7395
rect 12265 7361 12299 7395
rect 12299 7361 12308 7395
rect 12256 7352 12308 7361
rect 13268 7352 13320 7404
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 14464 7352 14516 7404
rect 15384 7352 15436 7404
rect 17868 7420 17920 7472
rect 14556 7284 14608 7336
rect 16764 7395 16816 7404
rect 16764 7361 16773 7395
rect 16773 7361 16807 7395
rect 16807 7361 16816 7395
rect 16764 7352 16816 7361
rect 17592 7395 17644 7404
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 20352 7420 20404 7472
rect 21364 7420 21416 7472
rect 18788 7395 18840 7404
rect 18788 7361 18822 7395
rect 18822 7361 18840 7395
rect 18788 7352 18840 7361
rect 22192 7352 22244 7404
rect 24860 7352 24912 7404
rect 28356 7395 28408 7404
rect 28356 7361 28365 7395
rect 28365 7361 28399 7395
rect 28399 7361 28408 7395
rect 28356 7352 28408 7361
rect 15476 7216 15528 7268
rect 18328 7284 18380 7336
rect 22836 7284 22888 7336
rect 25596 7327 25648 7336
rect 25596 7293 25605 7327
rect 25605 7293 25639 7327
rect 25639 7293 25648 7327
rect 25596 7284 25648 7293
rect 12440 7148 12492 7200
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 19892 7191 19944 7200
rect 19892 7157 19901 7191
rect 19901 7157 19935 7191
rect 19935 7157 19944 7191
rect 19892 7148 19944 7157
rect 22376 7191 22428 7200
rect 22376 7157 22385 7191
rect 22385 7157 22419 7191
rect 22419 7157 22428 7191
rect 22376 7148 22428 7157
rect 28172 7191 28224 7200
rect 28172 7157 28181 7191
rect 28181 7157 28215 7191
rect 28215 7157 28224 7191
rect 28172 7148 28224 7157
rect 5582 7046 5634 7098
rect 5646 7046 5698 7098
rect 5710 7046 5762 7098
rect 5774 7046 5826 7098
rect 5838 7046 5890 7098
rect 14846 7046 14898 7098
rect 14910 7046 14962 7098
rect 14974 7046 15026 7098
rect 15038 7046 15090 7098
rect 15102 7046 15154 7098
rect 24110 7046 24162 7098
rect 24174 7046 24226 7098
rect 24238 7046 24290 7098
rect 24302 7046 24354 7098
rect 24366 7046 24418 7098
rect 22192 6987 22244 6996
rect 22192 6953 22201 6987
rect 22201 6953 22235 6987
rect 22235 6953 22244 6987
rect 22192 6944 22244 6953
rect 12900 6808 12952 6860
rect 13728 6808 13780 6860
rect 18328 6876 18380 6928
rect 17592 6808 17644 6860
rect 19156 6808 19208 6860
rect 19984 6808 20036 6860
rect 22836 6876 22888 6928
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 22744 6808 22796 6817
rect 24860 6851 24912 6860
rect 24860 6817 24869 6851
rect 24869 6817 24903 6851
rect 24903 6817 24912 6851
rect 24860 6808 24912 6817
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 17684 6740 17736 6792
rect 12256 6672 12308 6724
rect 13360 6604 13412 6656
rect 14464 6604 14516 6656
rect 15844 6604 15896 6656
rect 19340 6740 19392 6792
rect 21272 6740 21324 6792
rect 22376 6740 22428 6792
rect 23664 6740 23716 6792
rect 16120 6604 16172 6656
rect 16856 6604 16908 6656
rect 17040 6604 17092 6656
rect 19248 6647 19300 6656
rect 19248 6613 19257 6647
rect 19257 6613 19291 6647
rect 19291 6613 19300 6647
rect 19248 6604 19300 6613
rect 20812 6604 20864 6656
rect 22100 6604 22152 6656
rect 22652 6647 22704 6656
rect 22652 6613 22661 6647
rect 22661 6613 22695 6647
rect 22695 6613 22704 6647
rect 22652 6604 22704 6613
rect 23664 6604 23716 6656
rect 24492 6740 24544 6792
rect 24584 6672 24636 6724
rect 28172 6672 28224 6724
rect 10214 6502 10266 6554
rect 10278 6502 10330 6554
rect 10342 6502 10394 6554
rect 10406 6502 10458 6554
rect 10470 6502 10522 6554
rect 19478 6502 19530 6554
rect 19542 6502 19594 6554
rect 19606 6502 19658 6554
rect 19670 6502 19722 6554
rect 19734 6502 19786 6554
rect 12256 6443 12308 6452
rect 12256 6409 12265 6443
rect 12265 6409 12299 6443
rect 12299 6409 12308 6443
rect 12256 6400 12308 6409
rect 17592 6400 17644 6452
rect 20812 6443 20864 6452
rect 20812 6409 20821 6443
rect 20821 6409 20855 6443
rect 20855 6409 20864 6443
rect 20812 6400 20864 6409
rect 16028 6332 16080 6384
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 17868 6332 17920 6384
rect 18328 6332 18380 6384
rect 24492 6400 24544 6452
rect 24860 6400 24912 6452
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 19800 6307 19852 6316
rect 19800 6273 19809 6307
rect 19809 6273 19843 6307
rect 19843 6273 19852 6307
rect 19800 6264 19852 6273
rect 20444 6264 20496 6316
rect 19984 6239 20036 6248
rect 14188 6128 14240 6180
rect 15844 6128 15896 6180
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 21088 6239 21140 6248
rect 21088 6205 21097 6239
rect 21097 6205 21131 6239
rect 21131 6205 21140 6239
rect 21088 6196 21140 6205
rect 23204 6307 23256 6316
rect 23204 6273 23213 6307
rect 23213 6273 23247 6307
rect 23247 6273 23256 6307
rect 23204 6264 23256 6273
rect 23664 6307 23716 6316
rect 23664 6273 23673 6307
rect 23673 6273 23707 6307
rect 23707 6273 23716 6307
rect 23664 6264 23716 6273
rect 23756 6264 23808 6316
rect 24676 6332 24728 6384
rect 22652 6239 22704 6248
rect 22652 6205 22661 6239
rect 22661 6205 22695 6239
rect 22695 6205 22704 6239
rect 22652 6196 22704 6205
rect 22836 6239 22888 6248
rect 22836 6205 22845 6239
rect 22845 6205 22879 6239
rect 22879 6205 22888 6239
rect 22836 6196 22888 6205
rect 15660 6103 15712 6112
rect 15660 6069 15669 6103
rect 15669 6069 15703 6103
rect 15703 6069 15712 6103
rect 15660 6060 15712 6069
rect 18144 6060 18196 6112
rect 19708 6060 19760 6112
rect 20628 6060 20680 6112
rect 22192 6103 22244 6112
rect 22192 6069 22201 6103
rect 22201 6069 22235 6103
rect 22235 6069 22244 6103
rect 22192 6060 22244 6069
rect 23296 6060 23348 6112
rect 5582 5958 5634 6010
rect 5646 5958 5698 6010
rect 5710 5958 5762 6010
rect 5774 5958 5826 6010
rect 5838 5958 5890 6010
rect 14846 5958 14898 6010
rect 14910 5958 14962 6010
rect 14974 5958 15026 6010
rect 15038 5958 15090 6010
rect 15102 5958 15154 6010
rect 24110 5958 24162 6010
rect 24174 5958 24226 6010
rect 24238 5958 24290 6010
rect 24302 5958 24354 6010
rect 24366 5958 24418 6010
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 19340 5899 19392 5908
rect 19340 5865 19349 5899
rect 19349 5865 19383 5899
rect 19383 5865 19392 5899
rect 19340 5856 19392 5865
rect 22100 5856 22152 5908
rect 22652 5856 22704 5908
rect 16856 5788 16908 5840
rect 19800 5788 19852 5840
rect 13728 5763 13780 5772
rect 13728 5729 13737 5763
rect 13737 5729 13771 5763
rect 13771 5729 13780 5763
rect 13728 5720 13780 5729
rect 18144 5763 18196 5772
rect 18144 5729 18153 5763
rect 18153 5729 18187 5763
rect 18187 5729 18196 5763
rect 18144 5720 18196 5729
rect 18328 5763 18380 5772
rect 18328 5729 18337 5763
rect 18337 5729 18371 5763
rect 18371 5729 18380 5763
rect 18328 5720 18380 5729
rect 13452 5695 13504 5704
rect 13452 5661 13470 5695
rect 13470 5661 13504 5695
rect 13452 5652 13504 5661
rect 17500 5652 17552 5704
rect 19708 5695 19760 5704
rect 19708 5661 19717 5695
rect 19717 5661 19751 5695
rect 19751 5661 19760 5695
rect 19708 5652 19760 5661
rect 20352 5720 20404 5772
rect 23756 5720 23808 5772
rect 21088 5652 21140 5704
rect 22284 5652 22336 5704
rect 22744 5652 22796 5704
rect 23296 5695 23348 5704
rect 23296 5661 23314 5695
rect 23314 5661 23348 5695
rect 28080 5695 28132 5704
rect 23296 5652 23348 5661
rect 28080 5661 28089 5695
rect 28089 5661 28123 5695
rect 28123 5661 28132 5695
rect 28080 5652 28132 5661
rect 15660 5584 15712 5636
rect 19892 5584 19944 5636
rect 20812 5627 20864 5636
rect 20812 5593 20846 5627
rect 20846 5593 20864 5627
rect 20812 5584 20864 5593
rect 12348 5559 12400 5568
rect 12348 5525 12357 5559
rect 12357 5525 12391 5559
rect 12391 5525 12400 5559
rect 12348 5516 12400 5525
rect 17960 5516 18012 5568
rect 28264 5559 28316 5568
rect 28264 5525 28273 5559
rect 28273 5525 28307 5559
rect 28307 5525 28316 5559
rect 28264 5516 28316 5525
rect 10214 5414 10266 5466
rect 10278 5414 10330 5466
rect 10342 5414 10394 5466
rect 10406 5414 10458 5466
rect 10470 5414 10522 5466
rect 19478 5414 19530 5466
rect 19542 5414 19594 5466
rect 19606 5414 19658 5466
rect 19670 5414 19722 5466
rect 19734 5414 19786 5466
rect 17960 5312 18012 5364
rect 20812 5355 20864 5364
rect 20812 5321 20821 5355
rect 20821 5321 20855 5355
rect 20855 5321 20864 5355
rect 20812 5312 20864 5321
rect 22192 5355 22244 5364
rect 22192 5321 22201 5355
rect 22201 5321 22235 5355
rect 22235 5321 22244 5355
rect 22192 5312 22244 5321
rect 23204 5312 23256 5364
rect 20352 5244 20404 5296
rect 22100 5287 22152 5296
rect 22100 5253 22109 5287
rect 22109 5253 22143 5287
rect 22143 5253 22152 5287
rect 22100 5244 22152 5253
rect 19248 5219 19300 5228
rect 19248 5185 19282 5219
rect 19282 5185 19300 5219
rect 19248 5176 19300 5185
rect 20628 5219 20680 5228
rect 20628 5185 20637 5219
rect 20637 5185 20671 5219
rect 20671 5185 20680 5219
rect 20628 5176 20680 5185
rect 22284 5108 22336 5160
rect 20444 5040 20496 5092
rect 5582 4870 5634 4922
rect 5646 4870 5698 4922
rect 5710 4870 5762 4922
rect 5774 4870 5826 4922
rect 5838 4870 5890 4922
rect 14846 4870 14898 4922
rect 14910 4870 14962 4922
rect 14974 4870 15026 4922
rect 15038 4870 15090 4922
rect 15102 4870 15154 4922
rect 24110 4870 24162 4922
rect 24174 4870 24226 4922
rect 24238 4870 24290 4922
rect 24302 4870 24354 4922
rect 24366 4870 24418 4922
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 28356 4607 28408 4616
rect 28356 4573 28365 4607
rect 28365 4573 28399 4607
rect 28399 4573 28408 4607
rect 28356 4564 28408 4573
rect 19064 4496 19116 4548
rect 10214 4326 10266 4378
rect 10278 4326 10330 4378
rect 10342 4326 10394 4378
rect 10406 4326 10458 4378
rect 10470 4326 10522 4378
rect 19478 4326 19530 4378
rect 19542 4326 19594 4378
rect 19606 4326 19658 4378
rect 19670 4326 19722 4378
rect 19734 4326 19786 4378
rect 5582 3782 5634 3834
rect 5646 3782 5698 3834
rect 5710 3782 5762 3834
rect 5774 3782 5826 3834
rect 5838 3782 5890 3834
rect 14846 3782 14898 3834
rect 14910 3782 14962 3834
rect 14974 3782 15026 3834
rect 15038 3782 15090 3834
rect 15102 3782 15154 3834
rect 24110 3782 24162 3834
rect 24174 3782 24226 3834
rect 24238 3782 24290 3834
rect 24302 3782 24354 3834
rect 24366 3782 24418 3834
rect 10214 3238 10266 3290
rect 10278 3238 10330 3290
rect 10342 3238 10394 3290
rect 10406 3238 10458 3290
rect 10470 3238 10522 3290
rect 19478 3238 19530 3290
rect 19542 3238 19594 3290
rect 19606 3238 19658 3290
rect 19670 3238 19722 3290
rect 19734 3238 19786 3290
rect 16580 3136 16632 3188
rect 17408 3136 17460 3188
rect 12348 3000 12400 3052
rect 17316 3043 17368 3052
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 24584 3000 24636 3052
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 5582 2694 5634 2746
rect 5646 2694 5698 2746
rect 5710 2694 5762 2746
rect 5774 2694 5826 2746
rect 5838 2694 5890 2746
rect 14846 2694 14898 2746
rect 14910 2694 14962 2746
rect 14974 2694 15026 2746
rect 15038 2694 15090 2746
rect 15102 2694 15154 2746
rect 24110 2694 24162 2746
rect 24174 2694 24226 2746
rect 24238 2694 24290 2746
rect 24302 2694 24354 2746
rect 24366 2694 24418 2746
rect 9220 2592 9272 2644
rect 15844 2592 15896 2644
rect 18052 2592 18104 2644
rect 24584 2635 24636 2644
rect 24584 2601 24593 2635
rect 24593 2601 24627 2635
rect 24627 2601 24636 2635
rect 24584 2592 24636 2601
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2596 2388 2648 2440
rect 6460 2388 6512 2440
rect 15936 2524 15988 2576
rect 17316 2456 17368 2508
rect 7748 2388 7800 2440
rect 10140 2388 10192 2440
rect 15476 2388 15528 2440
rect 18052 2388 18104 2440
rect 24492 2388 24544 2440
rect 25780 2388 25832 2440
rect 27068 2388 27120 2440
rect 27528 2388 27580 2440
rect 12624 2320 12676 2372
rect 1492 2295 1544 2304
rect 1492 2261 1501 2295
rect 1501 2261 1535 2295
rect 1535 2261 1544 2295
rect 1492 2252 1544 2261
rect 5172 2252 5224 2304
rect 20628 2252 20680 2304
rect 10214 2150 10266 2202
rect 10278 2150 10330 2202
rect 10342 2150 10394 2202
rect 10406 2150 10458 2202
rect 10470 2150 10522 2202
rect 19478 2150 19530 2202
rect 19542 2150 19594 2202
rect 19606 2150 19658 2202
rect 19670 2150 19722 2202
rect 19734 2150 19786 2202
<< metal2 >>
rect 18 29200 74 30000
rect 1950 29322 2006 30000
rect 3238 29322 3294 30000
rect 1950 29294 2084 29322
rect 1950 29200 2006 29294
rect 1398 28656 1454 28665
rect 1398 28591 1454 28600
rect 1412 27470 1440 28591
rect 2056 27606 2084 29294
rect 3238 29294 3372 29322
rect 3238 29200 3294 29294
rect 3344 27606 3372 29294
rect 4526 29200 4582 30000
rect 5814 29322 5870 30000
rect 5814 29294 6224 29322
rect 5814 29200 5870 29294
rect 5582 27772 5890 27792
rect 5582 27770 5588 27772
rect 5644 27770 5668 27772
rect 5724 27770 5748 27772
rect 5804 27770 5828 27772
rect 5884 27770 5890 27772
rect 5644 27718 5646 27770
rect 5826 27718 5828 27770
rect 5582 27716 5588 27718
rect 5644 27716 5668 27718
rect 5724 27716 5748 27718
rect 5804 27716 5828 27718
rect 5884 27716 5890 27718
rect 5582 27696 5890 27716
rect 6196 27606 6224 29294
rect 7102 29200 7158 30000
rect 8390 29200 8446 30000
rect 9678 29200 9734 30000
rect 10966 29200 11022 30000
rect 12254 29322 12310 30000
rect 13542 29322 13598 30000
rect 12254 29294 12388 29322
rect 12254 29200 12310 29294
rect 12360 27606 12388 29294
rect 13542 29294 13768 29322
rect 13542 29200 13598 29294
rect 2044 27600 2096 27606
rect 2044 27542 2096 27548
rect 3332 27600 3384 27606
rect 3332 27542 3384 27548
rect 6184 27600 6236 27606
rect 6184 27542 6236 27548
rect 12348 27600 12400 27606
rect 13740 27588 13768 29294
rect 14830 29200 14886 30000
rect 16118 29200 16174 30000
rect 17406 29200 17462 30000
rect 18694 29200 18750 30000
rect 19982 29200 20038 30000
rect 21270 29200 21326 30000
rect 22558 29200 22614 30000
rect 23846 29200 23902 30000
rect 25134 29200 25190 30000
rect 26422 29322 26478 30000
rect 27710 29322 27766 30000
rect 26422 29294 26556 29322
rect 26422 29200 26478 29294
rect 14844 27962 14872 29200
rect 14752 27934 14872 27962
rect 14752 27606 14780 27934
rect 14846 27772 15154 27792
rect 14846 27770 14852 27772
rect 14908 27770 14932 27772
rect 14988 27770 15012 27772
rect 15068 27770 15092 27772
rect 15148 27770 15154 27772
rect 14908 27718 14910 27770
rect 15090 27718 15092 27770
rect 14846 27716 14852 27718
rect 14908 27716 14932 27718
rect 14988 27716 15012 27718
rect 15068 27716 15092 27718
rect 15148 27716 15154 27718
rect 14846 27696 15154 27716
rect 16132 27606 16160 29200
rect 18708 27606 18736 29200
rect 19996 27606 20024 29200
rect 21284 27606 21312 29200
rect 13820 27600 13872 27606
rect 13740 27560 13820 27588
rect 12348 27542 12400 27548
rect 13820 27542 13872 27548
rect 14740 27600 14792 27606
rect 14740 27542 14792 27548
rect 16120 27600 16172 27606
rect 16120 27542 16172 27548
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 19984 27600 20036 27606
rect 19984 27542 20036 27548
rect 21272 27600 21324 27606
rect 21272 27542 21324 27548
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 1400 27464 1452 27470
rect 13728 27464 13780 27470
rect 1452 27412 1532 27418
rect 1400 27406 1532 27412
rect 13728 27406 13780 27412
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 16304 27464 16356 27470
rect 16304 27406 16356 27412
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 1412 27390 1532 27406
rect 1398 27296 1454 27305
rect 1398 27231 1454 27240
rect 1412 26994 1440 27231
rect 1504 27130 1532 27390
rect 4436 27396 4488 27402
rect 4436 27338 4488 27344
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1492 27124 1544 27130
rect 1492 27066 1544 27072
rect 1400 26988 1452 26994
rect 1400 26930 1452 26936
rect 1400 23520 1452 23526
rect 1400 23462 1452 23468
rect 1412 23225 1440 23462
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1412 21865 1440 21966
rect 1398 21856 1454 21865
rect 1398 21791 1454 21800
rect 1400 17808 1452 17814
rect 1398 17776 1400 17785
rect 1452 17776 1454 17785
rect 1398 17711 1454 17720
rect 1492 16448 1544 16454
rect 1398 16416 1454 16425
rect 1492 16390 1544 16396
rect 1398 16351 1454 16360
rect 1412 16114 1440 16351
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1504 8498 1532 16390
rect 1596 12102 1624 27270
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 1688 25945 1716 26318
rect 1768 26308 1820 26314
rect 1768 26250 1820 26256
rect 1674 25936 1730 25945
rect 1674 25871 1730 25880
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1596 9625 1624 9930
rect 1582 9616 1638 9625
rect 1582 9551 1638 9560
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 8265 1624 8298
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1412 4185 1440 4558
rect 1398 4176 1454 4185
rect 1398 4111 1454 4120
rect 1492 2848 1544 2854
rect 1490 2816 1492 2825
rect 1544 2816 1546 2825
rect 1490 2751 1546 2760
rect 1688 2446 1716 18022
rect 1780 12209 1808 26250
rect 4448 22098 4476 27338
rect 10214 27228 10522 27248
rect 10214 27226 10220 27228
rect 10276 27226 10300 27228
rect 10356 27226 10380 27228
rect 10436 27226 10460 27228
rect 10516 27226 10522 27228
rect 10276 27174 10278 27226
rect 10458 27174 10460 27226
rect 10214 27172 10220 27174
rect 10276 27172 10300 27174
rect 10356 27172 10380 27174
rect 10436 27172 10460 27174
rect 10516 27172 10522 27174
rect 10214 27152 10522 27172
rect 5582 26684 5890 26704
rect 5582 26682 5588 26684
rect 5644 26682 5668 26684
rect 5724 26682 5748 26684
rect 5804 26682 5828 26684
rect 5884 26682 5890 26684
rect 5644 26630 5646 26682
rect 5826 26630 5828 26682
rect 5582 26628 5588 26630
rect 5644 26628 5668 26630
rect 5724 26628 5748 26630
rect 5804 26628 5828 26630
rect 5884 26628 5890 26630
rect 5582 26608 5890 26628
rect 10214 26140 10522 26160
rect 10214 26138 10220 26140
rect 10276 26138 10300 26140
rect 10356 26138 10380 26140
rect 10436 26138 10460 26140
rect 10516 26138 10522 26140
rect 10276 26086 10278 26138
rect 10458 26086 10460 26138
rect 10214 26084 10220 26086
rect 10276 26084 10300 26086
rect 10356 26084 10380 26086
rect 10436 26084 10460 26086
rect 10516 26084 10522 26086
rect 10214 26064 10522 26084
rect 5582 25596 5890 25616
rect 5582 25594 5588 25596
rect 5644 25594 5668 25596
rect 5724 25594 5748 25596
rect 5804 25594 5828 25596
rect 5884 25594 5890 25596
rect 5644 25542 5646 25594
rect 5826 25542 5828 25594
rect 5582 25540 5588 25542
rect 5644 25540 5668 25542
rect 5724 25540 5748 25542
rect 5804 25540 5828 25542
rect 5884 25540 5890 25542
rect 5582 25520 5890 25540
rect 10214 25052 10522 25072
rect 10214 25050 10220 25052
rect 10276 25050 10300 25052
rect 10356 25050 10380 25052
rect 10436 25050 10460 25052
rect 10516 25050 10522 25052
rect 10276 24998 10278 25050
rect 10458 24998 10460 25050
rect 10214 24996 10220 24998
rect 10276 24996 10300 24998
rect 10356 24996 10380 24998
rect 10436 24996 10460 24998
rect 10516 24996 10522 24998
rect 10214 24976 10522 24996
rect 5582 24508 5890 24528
rect 5582 24506 5588 24508
rect 5644 24506 5668 24508
rect 5724 24506 5748 24508
rect 5804 24506 5828 24508
rect 5884 24506 5890 24508
rect 5644 24454 5646 24506
rect 5826 24454 5828 24506
rect 5582 24452 5588 24454
rect 5644 24452 5668 24454
rect 5724 24452 5748 24454
rect 5804 24452 5828 24454
rect 5884 24452 5890 24454
rect 5582 24432 5890 24452
rect 13740 24410 13768 27406
rect 14660 27130 14688 27406
rect 16316 27130 16344 27406
rect 17960 27328 18012 27334
rect 17960 27270 18012 27276
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 16304 27124 16356 27130
rect 16304 27066 16356 27072
rect 17972 27062 18000 27270
rect 14740 27056 14792 27062
rect 14740 26998 14792 27004
rect 15384 27056 15436 27062
rect 15384 26998 15436 27004
rect 17960 27056 18012 27062
rect 17960 26998 18012 27004
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 10214 23964 10522 23984
rect 10214 23962 10220 23964
rect 10276 23962 10300 23964
rect 10356 23962 10380 23964
rect 10436 23962 10460 23964
rect 10516 23962 10522 23964
rect 10276 23910 10278 23962
rect 10458 23910 10460 23962
rect 10214 23908 10220 23910
rect 10276 23908 10300 23910
rect 10356 23908 10380 23910
rect 10436 23908 10460 23910
rect 10516 23908 10522 23910
rect 10214 23888 10522 23908
rect 5582 23420 5890 23440
rect 5582 23418 5588 23420
rect 5644 23418 5668 23420
rect 5724 23418 5748 23420
rect 5804 23418 5828 23420
rect 5884 23418 5890 23420
rect 5644 23366 5646 23418
rect 5826 23366 5828 23418
rect 5582 23364 5588 23366
rect 5644 23364 5668 23366
rect 5724 23364 5748 23366
rect 5804 23364 5828 23366
rect 5884 23364 5890 23366
rect 5582 23344 5890 23364
rect 10214 22876 10522 22896
rect 10214 22874 10220 22876
rect 10276 22874 10300 22876
rect 10356 22874 10380 22876
rect 10436 22874 10460 22876
rect 10516 22874 10522 22876
rect 10276 22822 10278 22874
rect 10458 22822 10460 22874
rect 10214 22820 10220 22822
rect 10276 22820 10300 22822
rect 10356 22820 10380 22822
rect 10436 22820 10460 22822
rect 10516 22820 10522 22822
rect 10214 22800 10522 22820
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 5582 22332 5890 22352
rect 5582 22330 5588 22332
rect 5644 22330 5668 22332
rect 5724 22330 5748 22332
rect 5804 22330 5828 22332
rect 5884 22330 5890 22332
rect 5644 22278 5646 22330
rect 5826 22278 5828 22330
rect 5582 22276 5588 22278
rect 5644 22276 5668 22278
rect 5724 22276 5748 22278
rect 5804 22276 5828 22278
rect 5884 22276 5890 22278
rect 5582 22256 5890 22276
rect 4436 22092 4488 22098
rect 4436 22034 4488 22040
rect 11992 21962 12020 22374
rect 11980 21956 12032 21962
rect 11980 21898 12032 21904
rect 10214 21788 10522 21808
rect 10214 21786 10220 21788
rect 10276 21786 10300 21788
rect 10356 21786 10380 21788
rect 10436 21786 10460 21788
rect 10516 21786 10522 21788
rect 10276 21734 10278 21786
rect 10458 21734 10460 21786
rect 10214 21732 10220 21734
rect 10276 21732 10300 21734
rect 10356 21732 10380 21734
rect 10436 21732 10460 21734
rect 10516 21732 10522 21734
rect 10214 21712 10522 21732
rect 11520 21480 11572 21486
rect 11520 21422 11572 21428
rect 5582 21244 5890 21264
rect 5582 21242 5588 21244
rect 5644 21242 5668 21244
rect 5724 21242 5748 21244
rect 5804 21242 5828 21244
rect 5884 21242 5890 21244
rect 5644 21190 5646 21242
rect 5826 21190 5828 21242
rect 5582 21188 5588 21190
rect 5644 21188 5668 21190
rect 5724 21188 5748 21190
rect 5804 21188 5828 21190
rect 5884 21188 5890 21190
rect 5582 21168 5890 21188
rect 10214 20700 10522 20720
rect 10214 20698 10220 20700
rect 10276 20698 10300 20700
rect 10356 20698 10380 20700
rect 10436 20698 10460 20700
rect 10516 20698 10522 20700
rect 10276 20646 10278 20698
rect 10458 20646 10460 20698
rect 10214 20644 10220 20646
rect 10276 20644 10300 20646
rect 10356 20644 10380 20646
rect 10436 20644 10460 20646
rect 10516 20644 10522 20646
rect 10214 20624 10522 20644
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 5582 20156 5890 20176
rect 5582 20154 5588 20156
rect 5644 20154 5668 20156
rect 5724 20154 5748 20156
rect 5804 20154 5828 20156
rect 5884 20154 5890 20156
rect 5644 20102 5646 20154
rect 5826 20102 5828 20154
rect 5582 20100 5588 20102
rect 5644 20100 5668 20102
rect 5724 20100 5748 20102
rect 5804 20100 5828 20102
rect 5884 20100 5890 20102
rect 5582 20080 5890 20100
rect 8404 19854 8432 20198
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8864 19718 8892 20334
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 5582 19068 5890 19088
rect 5582 19066 5588 19068
rect 5644 19066 5668 19068
rect 5724 19066 5748 19068
rect 5804 19066 5828 19068
rect 5884 19066 5890 19068
rect 5644 19014 5646 19066
rect 5826 19014 5828 19066
rect 5582 19012 5588 19014
rect 5644 19012 5668 19014
rect 5724 19012 5748 19014
rect 5804 19012 5828 19014
rect 5884 19012 5890 19014
rect 5582 18992 5890 19012
rect 8312 18766 8340 19178
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6656 18222 6684 18634
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6932 18358 6960 18566
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 5184 15570 5212 18158
rect 5582 17980 5890 18000
rect 5582 17978 5588 17980
rect 5644 17978 5668 17980
rect 5724 17978 5748 17980
rect 5804 17978 5828 17980
rect 5884 17978 5890 17980
rect 5644 17926 5646 17978
rect 5826 17926 5828 17978
rect 5582 17924 5588 17926
rect 5644 17924 5668 17926
rect 5724 17924 5748 17926
rect 5804 17924 5828 17926
rect 5884 17924 5890 17926
rect 5582 17904 5890 17924
rect 7116 17882 7144 18702
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7208 17678 7236 17818
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7208 17202 7236 17614
rect 7392 17338 7420 18362
rect 8312 17678 8340 18702
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8404 17746 8432 18022
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 5582 16892 5890 16912
rect 5582 16890 5588 16892
rect 5644 16890 5668 16892
rect 5724 16890 5748 16892
rect 5804 16890 5828 16892
rect 5884 16890 5890 16892
rect 5644 16838 5646 16890
rect 5826 16838 5828 16890
rect 5582 16836 5588 16838
rect 5644 16836 5668 16838
rect 5724 16836 5748 16838
rect 5804 16836 5828 16838
rect 5884 16836 5890 16838
rect 5582 16816 5890 16836
rect 6012 16590 6040 16934
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5460 15502 5488 15846
rect 5582 15804 5890 15824
rect 5582 15802 5588 15804
rect 5644 15802 5668 15804
rect 5724 15802 5748 15804
rect 5804 15802 5828 15804
rect 5884 15802 5890 15804
rect 5644 15750 5646 15802
rect 5826 15750 5828 15802
rect 5582 15748 5588 15750
rect 5644 15748 5668 15750
rect 5724 15748 5748 15750
rect 5804 15748 5828 15750
rect 5884 15748 5890 15750
rect 5582 15728 5890 15748
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4080 15065 4108 15098
rect 5920 15094 5948 16050
rect 5908 15088 5960 15094
rect 4066 15056 4122 15065
rect 5908 15030 5960 15036
rect 4066 14991 4122 15000
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5582 14716 5890 14736
rect 5582 14714 5588 14716
rect 5644 14714 5668 14716
rect 5724 14714 5748 14716
rect 5804 14714 5828 14716
rect 5884 14714 5890 14716
rect 5644 14662 5646 14714
rect 5826 14662 5828 14714
rect 5582 14660 5588 14662
rect 5644 14660 5668 14662
rect 5724 14660 5748 14662
rect 5804 14660 5828 14662
rect 5884 14660 5890 14662
rect 5582 14640 5890 14660
rect 5920 14278 5948 14894
rect 6748 14890 6776 16934
rect 7116 16454 7144 17070
rect 7392 16658 7420 17274
rect 7668 17134 7696 17478
rect 8404 17134 8432 17478
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8404 16794 8432 17070
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 14958 6868 15302
rect 7116 15026 7144 16390
rect 7852 16114 7880 16390
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7208 15094 7236 15302
rect 7196 15088 7248 15094
rect 7196 15030 7248 15036
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6550 14376 6606 14385
rect 6550 14311 6606 14320
rect 6564 14278 6592 14311
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 5582 13628 5890 13648
rect 5582 13626 5588 13628
rect 5644 13626 5668 13628
rect 5724 13626 5748 13628
rect 5804 13626 5828 13628
rect 5884 13626 5890 13628
rect 5644 13574 5646 13626
rect 5826 13574 5828 13626
rect 5582 13572 5588 13574
rect 5644 13572 5668 13574
rect 5724 13572 5748 13574
rect 5804 13572 5828 13574
rect 5884 13572 5890 13574
rect 5582 13552 5890 13572
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5184 12306 5212 13330
rect 5920 13326 5948 14010
rect 6564 13870 6592 14214
rect 6748 13954 6776 14826
rect 6840 14006 6868 14894
rect 7576 14890 7604 16050
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7760 15502 7788 15846
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 8220 14958 8248 16526
rect 8496 15450 8524 19314
rect 8864 19310 8892 19654
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8864 17882 8892 19246
rect 8956 18698 8984 19790
rect 9692 19514 9720 20402
rect 11532 20398 11560 21422
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9876 19378 9904 19654
rect 10214 19612 10522 19632
rect 10214 19610 10220 19612
rect 10276 19610 10300 19612
rect 10356 19610 10380 19612
rect 10436 19610 10460 19612
rect 10516 19610 10522 19612
rect 10276 19558 10278 19610
rect 10458 19558 10460 19610
rect 10214 19556 10220 19558
rect 10276 19556 10300 19558
rect 10356 19556 10380 19558
rect 10436 19556 10460 19558
rect 10516 19556 10522 19558
rect 10214 19536 10522 19556
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 9048 18970 9076 19314
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 8944 18692 8996 18698
rect 8944 18634 8996 18640
rect 9048 18222 9076 18770
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9416 18222 9444 18634
rect 9508 18290 9536 19110
rect 9876 18766 9904 19314
rect 10324 19304 10376 19310
rect 10322 19272 10324 19281
rect 10376 19272 10378 19281
rect 10322 19207 10378 19216
rect 10336 18834 10364 19207
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9048 17898 9076 18158
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8956 17870 9076 17898
rect 8956 17814 8984 17870
rect 8944 17808 8996 17814
rect 8944 17750 8996 17756
rect 9232 17678 9260 18022
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8956 16794 8984 17138
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 8576 16720 8628 16726
rect 9784 16697 9812 16934
rect 8576 16662 8628 16668
rect 9770 16688 9826 16697
rect 8588 15570 8616 16662
rect 9770 16623 9826 16632
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 16250 9168 16526
rect 9784 16454 9812 16623
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8496 15422 8616 15450
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 6656 13926 6776 13954
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 6564 12918 6592 13806
rect 6656 13734 6684 13926
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 6000 12912 6052 12918
rect 6000 12854 6052 12860
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 5828 12782 5856 12854
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5276 12238 5304 12582
rect 5582 12540 5890 12560
rect 5582 12538 5588 12540
rect 5644 12538 5668 12540
rect 5724 12538 5748 12540
rect 5804 12538 5828 12540
rect 5884 12538 5890 12540
rect 5644 12486 5646 12538
rect 5826 12486 5828 12538
rect 5582 12484 5588 12486
rect 5644 12484 5668 12486
rect 5724 12484 5748 12486
rect 5804 12484 5828 12486
rect 5884 12484 5890 12486
rect 5582 12464 5890 12484
rect 5264 12232 5316 12238
rect 1766 12200 1822 12209
rect 5264 12174 5316 12180
rect 1766 12135 1822 12144
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1780 8945 1808 12038
rect 6012 11898 6040 12854
rect 6656 12850 6684 13670
rect 6748 13394 6776 13738
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7208 13530 7236 13670
rect 7576 13530 7604 14350
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8036 14006 8064 14214
rect 8220 14006 8248 14894
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6748 12986 6776 13330
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 7852 12850 7880 13670
rect 8220 13394 8248 13942
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6564 12374 6592 12718
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6656 12306 6684 12786
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6656 11762 6684 12038
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 7300 11694 7328 12038
rect 7760 11762 7788 12038
rect 7944 11898 7972 12786
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7288 11688 7340 11694
rect 8220 11642 8248 12174
rect 8588 11898 8616 15422
rect 9232 14958 9260 15982
rect 9588 15972 9640 15978
rect 9588 15914 9640 15920
rect 9600 15570 9628 15914
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9232 14482 9260 14894
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8956 13841 8984 14010
rect 8942 13832 8998 13841
rect 8942 13767 8998 13776
rect 8956 13326 8984 13767
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 8852 12436 8904 12442
rect 9140 12434 9168 13194
rect 9232 12986 9260 13262
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9324 12714 9352 14282
rect 9416 14074 9444 14962
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9784 13734 9812 14418
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9692 12730 9720 13398
rect 9784 13326 9812 13670
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9876 12782 9904 18702
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9968 18086 9996 18566
rect 10214 18524 10522 18544
rect 10214 18522 10220 18524
rect 10276 18522 10300 18524
rect 10356 18522 10380 18524
rect 10436 18522 10460 18524
rect 10516 18522 10522 18524
rect 10276 18470 10278 18522
rect 10458 18470 10460 18522
rect 10214 18468 10220 18470
rect 10276 18468 10300 18470
rect 10356 18468 10380 18470
rect 10436 18468 10460 18470
rect 10516 18468 10522 18470
rect 10214 18448 10522 18468
rect 10782 18320 10838 18329
rect 10782 18255 10838 18264
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9968 17542 9996 18022
rect 10796 17542 10824 18255
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 9968 16250 9996 17478
rect 10214 17436 10522 17456
rect 10214 17434 10220 17436
rect 10276 17434 10300 17436
rect 10356 17434 10380 17436
rect 10436 17434 10460 17436
rect 10516 17434 10522 17436
rect 10276 17382 10278 17434
rect 10458 17382 10460 17434
rect 10214 17380 10220 17382
rect 10276 17380 10300 17382
rect 10356 17380 10380 17382
rect 10436 17380 10460 17382
rect 10516 17380 10522 17382
rect 10214 17360 10522 17380
rect 10214 16348 10522 16368
rect 10214 16346 10220 16348
rect 10276 16346 10300 16348
rect 10356 16346 10380 16348
rect 10436 16346 10460 16348
rect 10516 16346 10522 16348
rect 10276 16294 10278 16346
rect 10458 16294 10460 16346
rect 10214 16292 10220 16294
rect 10276 16292 10300 16294
rect 10356 16292 10380 16294
rect 10436 16292 10460 16294
rect 10516 16292 10522 16294
rect 10214 16272 10522 16292
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 9968 14770 9996 15982
rect 10704 15910 10732 16118
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 10060 14890 10088 15370
rect 10152 15026 10180 15846
rect 10214 15260 10522 15280
rect 10214 15258 10220 15260
rect 10276 15258 10300 15260
rect 10356 15258 10380 15260
rect 10436 15258 10460 15260
rect 10516 15258 10522 15260
rect 10276 15206 10278 15258
rect 10458 15206 10460 15258
rect 10214 15204 10220 15206
rect 10276 15204 10300 15206
rect 10356 15204 10380 15206
rect 10436 15204 10460 15206
rect 10516 15204 10522 15206
rect 10214 15184 10522 15204
rect 10704 15162 10732 15846
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 10140 14816 10192 14822
rect 9968 14742 10088 14770
rect 10140 14758 10192 14764
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9968 12850 9996 14350
rect 10060 14006 10088 14742
rect 10152 14414 10180 14758
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10214 14172 10522 14192
rect 10214 14170 10220 14172
rect 10276 14170 10300 14172
rect 10356 14170 10380 14172
rect 10436 14170 10460 14172
rect 10516 14170 10522 14172
rect 10276 14118 10278 14170
rect 10458 14118 10460 14170
rect 10214 14116 10220 14118
rect 10276 14116 10300 14118
rect 10356 14116 10380 14118
rect 10436 14116 10460 14118
rect 10516 14116 10522 14118
rect 10214 14096 10522 14116
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10214 13084 10522 13104
rect 10214 13082 10220 13084
rect 10276 13082 10300 13084
rect 10356 13082 10380 13084
rect 10436 13082 10460 13084
rect 10516 13082 10522 13084
rect 10276 13030 10278 13082
rect 10458 13030 10460 13082
rect 10214 13028 10220 13030
rect 10276 13028 10300 13030
rect 10356 13028 10380 13030
rect 10436 13028 10460 13030
rect 10516 13028 10522 13030
rect 10214 13008 10522 13028
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9864 12776 9916 12782
rect 9600 12714 9812 12730
rect 9864 12718 9916 12724
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9588 12708 9812 12714
rect 9640 12702 9812 12708
rect 9588 12650 9640 12656
rect 9140 12406 9260 12434
rect 8852 12378 8904 12384
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 7288 11630 7340 11636
rect 5582 11452 5890 11472
rect 5582 11450 5588 11452
rect 5644 11450 5668 11452
rect 5724 11450 5748 11452
rect 5804 11450 5828 11452
rect 5884 11450 5890 11452
rect 5644 11398 5646 11450
rect 5826 11398 5828 11450
rect 5582 11396 5588 11398
rect 5644 11396 5668 11398
rect 5724 11396 5748 11398
rect 5804 11396 5828 11398
rect 5884 11396 5890 11398
rect 5582 11376 5890 11396
rect 7300 11354 7328 11630
rect 8036 11614 8248 11642
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7392 11150 7420 11494
rect 8036 11150 8064 11614
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11150 8248 11494
rect 8588 11354 8616 11834
rect 8864 11762 8892 12378
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8312 10742 8340 11154
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 5582 10364 5890 10384
rect 5582 10362 5588 10364
rect 5644 10362 5668 10364
rect 5724 10362 5748 10364
rect 5804 10362 5828 10364
rect 5884 10362 5890 10364
rect 5644 10310 5646 10362
rect 5826 10310 5828 10362
rect 5582 10308 5588 10310
rect 5644 10308 5668 10310
rect 5724 10308 5748 10310
rect 5804 10308 5828 10310
rect 5884 10308 5890 10310
rect 5582 10288 5890 10308
rect 8312 10130 8340 10678
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8588 9722 8616 10610
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8772 9586 8800 11018
rect 8864 10810 8892 11698
rect 9140 11694 9168 12242
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9232 11626 9260 12406
rect 9324 12238 9352 12650
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9416 12442 9444 12582
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 5582 9276 5890 9296
rect 5582 9274 5588 9276
rect 5644 9274 5668 9276
rect 5724 9274 5748 9276
rect 5804 9274 5828 9276
rect 5884 9274 5890 9276
rect 5644 9222 5646 9274
rect 5826 9222 5828 9274
rect 5582 9220 5588 9222
rect 5644 9220 5668 9222
rect 5724 9220 5748 9222
rect 5804 9220 5828 9222
rect 5884 9220 5890 9222
rect 5582 9200 5890 9220
rect 8956 9042 8984 10066
rect 9232 10062 9260 11562
rect 9324 10130 9352 11630
rect 9508 11286 9536 11698
rect 9496 11280 9548 11286
rect 9692 11257 9720 12038
rect 9496 11222 9548 11228
rect 9678 11248 9734 11257
rect 9678 11183 9734 11192
rect 9784 11200 9812 12702
rect 9968 12170 9996 12786
rect 10612 12782 10640 13942
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 10214 11996 10522 12016
rect 10214 11994 10220 11996
rect 10276 11994 10300 11996
rect 10356 11994 10380 11996
rect 10436 11994 10460 11996
rect 10516 11994 10522 11996
rect 10276 11942 10278 11994
rect 10458 11942 10460 11994
rect 10214 11940 10220 11942
rect 10276 11940 10300 11942
rect 10356 11940 10380 11942
rect 10436 11940 10460 11942
rect 10516 11940 10522 11942
rect 10214 11920 10522 11940
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9692 10266 9720 11183
rect 9784 11172 9904 11200
rect 9876 11082 9904 11172
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9876 10606 9904 11018
rect 10152 10810 10180 11290
rect 10214 10908 10522 10928
rect 10214 10906 10220 10908
rect 10276 10906 10300 10908
rect 10356 10906 10380 10908
rect 10436 10906 10460 10908
rect 10516 10906 10522 10908
rect 10276 10854 10278 10906
rect 10458 10854 10460 10906
rect 10214 10852 10220 10854
rect 10276 10852 10300 10854
rect 10356 10852 10380 10854
rect 10436 10852 10460 10854
rect 10516 10852 10522 10854
rect 10214 10832 10522 10852
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9600 9722 9628 9930
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9784 9586 9812 10406
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8392 8968 8444 8974
rect 1766 8936 1822 8945
rect 8392 8910 8444 8916
rect 1766 8871 1822 8880
rect 8404 8634 8432 8910
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 5582 8188 5890 8208
rect 5582 8186 5588 8188
rect 5644 8186 5668 8188
rect 5724 8186 5748 8188
rect 5804 8186 5828 8188
rect 5884 8186 5890 8188
rect 5644 8134 5646 8186
rect 5826 8134 5828 8186
rect 5582 8132 5588 8134
rect 5644 8132 5668 8134
rect 5724 8132 5748 8134
rect 5804 8132 5828 8134
rect 5884 8132 5890 8134
rect 5582 8112 5890 8132
rect 5582 7100 5890 7120
rect 5582 7098 5588 7100
rect 5644 7098 5668 7100
rect 5724 7098 5748 7100
rect 5804 7098 5828 7100
rect 5884 7098 5890 7100
rect 5644 7046 5646 7098
rect 5826 7046 5828 7098
rect 5582 7044 5588 7046
rect 5644 7044 5668 7046
rect 5724 7044 5748 7046
rect 5804 7044 5828 7046
rect 5884 7044 5890 7046
rect 5582 7024 5890 7044
rect 5582 6012 5890 6032
rect 5582 6010 5588 6012
rect 5644 6010 5668 6012
rect 5724 6010 5748 6012
rect 5804 6010 5828 6012
rect 5884 6010 5890 6012
rect 5644 5958 5646 6010
rect 5826 5958 5828 6010
rect 5582 5956 5588 5958
rect 5644 5956 5668 5958
rect 5724 5956 5748 5958
rect 5804 5956 5828 5958
rect 5884 5956 5890 5958
rect 5582 5936 5890 5956
rect 5582 4924 5890 4944
rect 5582 4922 5588 4924
rect 5644 4922 5668 4924
rect 5724 4922 5748 4924
rect 5804 4922 5828 4924
rect 5884 4922 5890 4924
rect 5644 4870 5646 4922
rect 5826 4870 5828 4922
rect 5582 4868 5588 4870
rect 5644 4868 5668 4870
rect 5724 4868 5748 4870
rect 5804 4868 5828 4870
rect 5884 4868 5890 4870
rect 5582 4848 5890 4868
rect 5582 3836 5890 3856
rect 5582 3834 5588 3836
rect 5644 3834 5668 3836
rect 5724 3834 5748 3836
rect 5804 3834 5828 3836
rect 5884 3834 5890 3836
rect 5644 3782 5646 3834
rect 5826 3782 5828 3834
rect 5582 3780 5588 3782
rect 5644 3780 5668 3782
rect 5724 3780 5748 3782
rect 5804 3780 5828 3782
rect 5884 3780 5890 3782
rect 5582 3760 5890 3780
rect 5582 2748 5890 2768
rect 5582 2746 5588 2748
rect 5644 2746 5668 2748
rect 5724 2746 5748 2748
rect 5804 2746 5828 2748
rect 5884 2746 5890 2748
rect 5644 2694 5646 2746
rect 5826 2694 5828 2746
rect 5582 2692 5588 2694
rect 5644 2692 5668 2694
rect 5724 2692 5748 2694
rect 5804 2692 5828 2694
rect 5884 2692 5890 2694
rect 5582 2672 5890 2692
rect 9232 2650 9260 9318
rect 9876 8430 9904 10542
rect 10060 9722 10088 10610
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10214 9820 10522 9840
rect 10214 9818 10220 9820
rect 10276 9818 10300 9820
rect 10356 9818 10380 9820
rect 10436 9818 10460 9820
rect 10516 9818 10522 9820
rect 10276 9766 10278 9818
rect 10458 9766 10460 9818
rect 10214 9764 10220 9766
rect 10276 9764 10300 9766
rect 10356 9764 10380 9766
rect 10436 9764 10460 9766
rect 10516 9764 10522 9766
rect 10214 9744 10522 9764
rect 10704 9722 10732 9862
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10796 9450 10824 17478
rect 11072 17241 11100 18022
rect 11348 17610 11376 19314
rect 11532 18834 11560 20334
rect 11808 20058 11836 20402
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11992 19446 12020 21898
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12360 21146 12388 21490
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12256 20868 12308 20874
rect 12256 20810 12308 20816
rect 12268 20058 12296 20810
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12072 19848 12124 19854
rect 12070 19816 12072 19825
rect 12124 19816 12126 19825
rect 12070 19751 12126 19760
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11900 18970 11928 19314
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11520 18692 11572 18698
rect 11520 18634 11572 18640
rect 11532 18426 11560 18634
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11702 18320 11758 18329
rect 11520 18284 11572 18290
rect 11992 18290 12020 19110
rect 11702 18255 11704 18264
rect 11520 18226 11572 18232
rect 11756 18255 11758 18264
rect 11980 18284 12032 18290
rect 11704 18226 11756 18232
rect 11980 18226 12032 18232
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11058 17232 11114 17241
rect 11348 17202 11376 17546
rect 11532 17338 11560 18226
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11900 17542 11928 18022
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11058 17167 11060 17176
rect 11112 17167 11114 17176
rect 11336 17196 11388 17202
rect 11060 17138 11112 17144
rect 11336 17138 11388 17144
rect 11150 16416 11206 16425
rect 11150 16351 11206 16360
rect 11164 16250 11192 16351
rect 11152 16244 11204 16250
rect 11204 16204 11284 16232
rect 11152 16186 11204 16192
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11072 15706 11100 16050
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11150 13968 11206 13977
rect 11150 13903 11206 13912
rect 11164 13802 11192 13903
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12986 10916 13194
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10980 12850 11008 13126
rect 11072 12918 11100 13126
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11072 12345 11100 12718
rect 11164 12442 11192 13262
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 11058 12336 11114 12345
rect 11058 12271 11114 12280
rect 11072 12238 11100 12271
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10888 11150 10916 11834
rect 11164 11694 11192 12378
rect 11256 11898 11284 16204
rect 11348 15502 11376 17138
rect 11888 17060 11940 17066
rect 11808 17020 11888 17048
rect 11426 16960 11482 16969
rect 11426 16895 11482 16904
rect 11440 16794 11468 16895
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11440 15502 11468 16730
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11716 15638 11744 16662
rect 11808 16454 11836 17020
rect 11888 17002 11940 17008
rect 11992 16998 12020 17818
rect 12084 17202 12112 19654
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12176 18086 12204 18226
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11796 16448 11848 16454
rect 11900 16425 11928 16458
rect 11796 16390 11848 16396
rect 11886 16416 11942 16425
rect 11886 16351 11942 16360
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11808 15706 11836 16050
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11702 15192 11758 15201
rect 11702 15127 11758 15136
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11624 14278 11652 14554
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11624 14074 11652 14214
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11716 13938 11744 15127
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11808 14822 11836 14894
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11624 12986 11652 13194
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11808 12850 11836 14758
rect 11992 13814 12020 16934
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 12084 14482 12112 14962
rect 12176 14550 12204 17682
rect 12268 17678 12296 19994
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12256 17672 12308 17678
rect 12360 17660 12388 18158
rect 12440 17672 12492 17678
rect 12360 17632 12440 17660
rect 12256 17614 12308 17620
rect 12440 17614 12492 17620
rect 12268 15910 12296 17614
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12360 16590 12388 17478
rect 12452 17134 12480 17614
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12256 15632 12308 15638
rect 12256 15574 12308 15580
rect 12268 15502 12296 15574
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12360 15484 12388 16526
rect 12452 16522 12480 17070
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12452 15706 12480 16458
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12544 15586 12572 22374
rect 12716 21956 12768 21962
rect 12716 21898 12768 21904
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12636 20942 12664 21830
rect 12728 21690 12756 21898
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12636 19922 12664 20198
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12716 19848 12768 19854
rect 12714 19816 12716 19825
rect 12768 19816 12770 19825
rect 12714 19751 12770 19760
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12636 18290 12664 19110
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12636 17338 12664 17546
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12728 16726 12756 17138
rect 12820 16794 12848 24074
rect 13832 23322 13860 24142
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 13360 23044 13412 23050
rect 13360 22986 13412 22992
rect 13372 22030 13400 22986
rect 13832 22710 13860 23258
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13176 21072 13228 21078
rect 12898 21040 12954 21049
rect 13176 21014 13228 21020
rect 12898 20975 12954 20984
rect 12912 20942 12940 20975
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12912 19718 12940 20878
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13096 19922 13124 20538
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 18272 12940 19110
rect 13084 18692 13136 18698
rect 13084 18634 13136 18640
rect 13096 18426 13124 18634
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 12992 18284 13044 18290
rect 12912 18244 12992 18272
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12820 15638 12848 16594
rect 12808 15632 12860 15638
rect 12544 15558 12664 15586
rect 12808 15574 12860 15580
rect 12532 15496 12584 15502
rect 12360 15456 12532 15484
rect 12268 15162 12296 15438
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12268 14770 12296 15098
rect 12360 14958 12388 15456
rect 12532 15438 12584 15444
rect 12636 15178 12664 15558
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12544 15150 12664 15178
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12268 14742 12480 14770
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12254 13968 12310 13977
rect 12254 13903 12310 13912
rect 11900 13786 12020 13814
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11900 12322 11928 13786
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11992 12434 12020 12718
rect 11992 12406 12112 12434
rect 11900 12294 12020 12322
rect 12084 12306 12112 12406
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11520 12096 11572 12102
rect 11518 12064 11520 12073
rect 11572 12064 11574 12073
rect 11518 11999 11574 12008
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10888 10742 10916 11086
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 11164 10130 11192 11630
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11256 11014 11284 11494
rect 11900 11150 11928 12174
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11440 10062 11468 10406
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11716 9722 11744 10610
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 11256 9042 11284 9590
rect 11808 9586 11836 9930
rect 11992 9722 12020 12294
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12084 11898 12112 12242
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12176 11354 12204 12038
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 11980 9716 12032 9722
rect 11900 9676 11980 9704
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10214 8732 10522 8752
rect 10214 8730 10220 8732
rect 10276 8730 10300 8732
rect 10356 8730 10380 8732
rect 10436 8730 10460 8732
rect 10516 8730 10522 8732
rect 10276 8678 10278 8730
rect 10458 8678 10460 8730
rect 10214 8676 10220 8678
rect 10276 8676 10300 8678
rect 10356 8676 10380 8678
rect 10436 8676 10460 8678
rect 10516 8676 10522 8678
rect 10214 8656 10522 8676
rect 10612 8498 10640 8774
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 9864 8424 9916 8430
rect 10796 8401 10824 8434
rect 11256 8430 11284 8978
rect 11900 8974 11928 9676
rect 11980 9658 12032 9664
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11244 8424 11296 8430
rect 9864 8366 9916 8372
rect 10782 8392 10838 8401
rect 9876 7478 9904 8366
rect 11244 8366 11296 8372
rect 10782 8327 10838 8336
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10060 7546 10088 7822
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 10152 7410 10180 8230
rect 11532 8022 11560 8434
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11532 7818 11560 7958
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 10214 7644 10522 7664
rect 10214 7642 10220 7644
rect 10276 7642 10300 7644
rect 10356 7642 10380 7644
rect 10436 7642 10460 7644
rect 10516 7642 10522 7644
rect 10276 7590 10278 7642
rect 10458 7590 10460 7642
rect 10214 7588 10220 7590
rect 10276 7588 10300 7590
rect 10356 7588 10380 7590
rect 10436 7588 10460 7590
rect 10516 7588 10522 7590
rect 10214 7568 10522 7588
rect 11624 7546 11652 8910
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 8498 11928 8774
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11992 8022 12020 8910
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 12268 7886 12296 13903
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12360 12170 12388 13806
rect 12452 12986 12480 14742
rect 12544 14074 12572 15150
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12360 11150 12388 12106
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12452 10130 12480 11154
rect 12544 10538 12572 11698
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 9654 12480 10066
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12636 9110 12664 15030
rect 12728 15026 12756 15302
rect 12912 15201 12940 18244
rect 12992 18226 13044 18232
rect 13188 17954 13216 21014
rect 13372 20942 13400 21966
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13556 20534 13584 21898
rect 14016 21690 14044 26930
rect 14752 25362 14780 26998
rect 14846 26684 15154 26704
rect 14846 26682 14852 26684
rect 14908 26682 14932 26684
rect 14988 26682 15012 26684
rect 15068 26682 15092 26684
rect 15148 26682 15154 26684
rect 14908 26630 14910 26682
rect 15090 26630 15092 26682
rect 14846 26628 14852 26630
rect 14908 26628 14932 26630
rect 14988 26628 15012 26630
rect 15068 26628 15092 26630
rect 15148 26628 15154 26630
rect 14846 26608 15154 26628
rect 15292 25696 15344 25702
rect 15292 25638 15344 25644
rect 14846 25596 15154 25616
rect 14846 25594 14852 25596
rect 14908 25594 14932 25596
rect 14988 25594 15012 25596
rect 15068 25594 15092 25596
rect 15148 25594 15154 25596
rect 14908 25542 14910 25594
rect 15090 25542 15092 25594
rect 14846 25540 14852 25542
rect 14908 25540 14932 25542
rect 14988 25540 15012 25542
rect 15068 25540 15092 25542
rect 15148 25540 15154 25542
rect 14846 25520 15154 25540
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14752 24206 14780 25298
rect 15304 25226 15332 25638
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 14846 24508 15154 24528
rect 14846 24506 14852 24508
rect 14908 24506 14932 24508
rect 14988 24506 15012 24508
rect 15068 24506 15092 24508
rect 15148 24506 15154 24508
rect 14908 24454 14910 24506
rect 15090 24454 15092 24506
rect 14846 24452 14852 24454
rect 14908 24452 14932 24454
rect 14988 24452 15012 24454
rect 15068 24452 15092 24454
rect 15148 24452 15154 24454
rect 14846 24432 15154 24452
rect 15212 24342 15240 24550
rect 15200 24336 15252 24342
rect 15200 24278 15252 24284
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14832 24132 14884 24138
rect 14832 24074 14884 24080
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14464 23588 14516 23594
rect 14464 23530 14516 23536
rect 14476 23186 14504 23530
rect 14464 23180 14516 23186
rect 14464 23122 14516 23128
rect 14568 23118 14596 24006
rect 14844 23730 14872 24074
rect 14648 23724 14700 23730
rect 14648 23666 14700 23672
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14660 23322 14688 23666
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 14648 23316 14700 23322
rect 14648 23258 14700 23264
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14752 22710 14780 23462
rect 14846 23420 15154 23440
rect 14846 23418 14852 23420
rect 14908 23418 14932 23420
rect 14988 23418 15012 23420
rect 15068 23418 15092 23420
rect 15148 23418 15154 23420
rect 14908 23366 14910 23418
rect 15090 23366 15092 23418
rect 14846 23364 14852 23366
rect 14908 23364 14932 23366
rect 14988 23364 15012 23366
rect 15068 23364 15092 23366
rect 15148 23364 15154 23366
rect 14846 23344 15154 23364
rect 14740 22704 14792 22710
rect 14740 22646 14792 22652
rect 14846 22332 15154 22352
rect 14846 22330 14852 22332
rect 14908 22330 14932 22332
rect 14988 22330 15012 22332
rect 15068 22330 15092 22332
rect 15148 22330 15154 22332
rect 14908 22278 14910 22330
rect 15090 22278 15092 22330
rect 14846 22276 14852 22278
rect 14908 22276 14932 22278
rect 14988 22276 15012 22278
rect 15068 22276 15092 22278
rect 15148 22276 15154 22278
rect 14846 22256 15154 22276
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 13832 21078 13860 21558
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13556 18850 13584 20470
rect 13832 20466 13860 21014
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13648 18970 13676 19314
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13556 18822 13676 18850
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 13188 17926 13308 17954
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13096 17202 13124 17274
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12990 16824 13046 16833
rect 12990 16759 13046 16768
rect 13004 16658 13032 16759
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 13096 16590 13124 17138
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13096 16114 13124 16526
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13004 15638 13032 15846
rect 12992 15632 13044 15638
rect 12992 15574 13044 15580
rect 13084 15496 13136 15502
rect 12990 15464 13046 15473
rect 13084 15438 13136 15444
rect 12990 15399 13046 15408
rect 12898 15192 12954 15201
rect 12898 15127 12954 15136
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12912 14346 12940 14758
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 13004 14226 13032 15399
rect 13096 15026 13124 15438
rect 13188 15337 13216 15846
rect 13174 15328 13230 15337
rect 13280 15314 13308 17926
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13372 16794 13400 17478
rect 13464 17202 13492 17478
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13452 15496 13504 15502
rect 13450 15464 13452 15473
rect 13504 15464 13506 15473
rect 13450 15399 13506 15408
rect 13556 15366 13584 18090
rect 13648 16726 13676 18822
rect 13740 18290 13768 19654
rect 13832 19514 13860 19654
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 14016 18902 14044 21490
rect 14200 20942 14228 22034
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14188 20936 14240 20942
rect 14186 20904 14188 20913
rect 14240 20904 14242 20913
rect 14186 20839 14242 20848
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14108 20534 14136 20742
rect 14096 20528 14148 20534
rect 14096 20470 14148 20476
rect 14292 19990 14320 21966
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 14384 21554 14412 21830
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14846 21244 15154 21264
rect 14846 21242 14852 21244
rect 14908 21242 14932 21244
rect 14988 21242 15012 21244
rect 15068 21242 15092 21244
rect 15148 21242 15154 21244
rect 14908 21190 14910 21242
rect 15090 21190 15092 21242
rect 14846 21188 14852 21190
rect 14908 21188 14932 21190
rect 14988 21188 15012 21190
rect 15068 21188 15092 21190
rect 15148 21188 15154 21190
rect 14846 21168 15154 21188
rect 14738 21040 14794 21049
rect 14738 20975 14794 20984
rect 14752 20942 14780 20975
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 15200 20868 15252 20874
rect 15200 20810 15252 20816
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 15212 20262 15240 20810
rect 15304 20602 15332 20810
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 14846 20156 15154 20176
rect 14846 20154 14852 20156
rect 14908 20154 14932 20156
rect 14988 20154 15012 20156
rect 15068 20154 15092 20156
rect 15148 20154 15154 20156
rect 14908 20102 14910 20154
rect 15090 20102 15092 20154
rect 14846 20100 14852 20102
rect 14908 20100 14932 20102
rect 14988 20100 15012 20102
rect 15068 20100 15092 20102
rect 15148 20100 15154 20102
rect 14846 20080 15154 20100
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14924 19984 14976 19990
rect 14924 19926 14976 19932
rect 15108 19984 15160 19990
rect 15108 19926 15160 19932
rect 14936 19854 14964 19926
rect 15120 19854 15148 19926
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14924 19848 14976 19854
rect 15108 19848 15160 19854
rect 14924 19790 14976 19796
rect 15028 19808 15108 19836
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 13832 18358 13860 18838
rect 14200 18698 14228 19314
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13740 17202 13768 17614
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 13740 16250 13768 17138
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 16250 13860 16390
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13648 15706 13676 15982
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13452 15360 13504 15366
rect 13280 15286 13400 15314
rect 13452 15302 13504 15308
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13174 15263 13230 15272
rect 13372 15144 13400 15286
rect 13464 15178 13492 15302
rect 13464 15150 13584 15178
rect 13740 15162 13768 15438
rect 13280 15116 13400 15144
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13082 14920 13138 14929
rect 13082 14855 13084 14864
rect 13136 14855 13138 14864
rect 13084 14826 13136 14832
rect 12912 14198 13032 14226
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12986 12756 13126
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12912 12866 12940 14198
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13004 13938 13032 14010
rect 13096 13938 13124 14214
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12912 12838 13124 12866
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12716 12096 12768 12102
rect 12714 12064 12716 12073
rect 12768 12064 12770 12073
rect 12714 11999 12770 12008
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12728 10674 12756 11290
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10198 12756 10406
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12716 9648 12768 9654
rect 12714 9616 12716 9625
rect 12768 9616 12770 9625
rect 12714 9551 12770 9560
rect 12728 9450 12756 9551
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 7954 12572 8774
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 12268 7410 12296 7822
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 10214 6556 10522 6576
rect 10214 6554 10220 6556
rect 10276 6554 10300 6556
rect 10356 6554 10380 6556
rect 10436 6554 10460 6556
rect 10516 6554 10522 6556
rect 10276 6502 10278 6554
rect 10458 6502 10460 6554
rect 10214 6500 10220 6502
rect 10276 6500 10300 6502
rect 10356 6500 10380 6502
rect 10436 6500 10460 6502
rect 10516 6500 10522 6502
rect 10214 6480 10522 6500
rect 12268 6458 12296 6666
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12452 6322 12480 7142
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 10214 5468 10522 5488
rect 10214 5466 10220 5468
rect 10276 5466 10300 5468
rect 10356 5466 10380 5468
rect 10436 5466 10460 5468
rect 10516 5466 10522 5468
rect 10276 5414 10278 5466
rect 10458 5414 10460 5466
rect 10214 5412 10220 5414
rect 10276 5412 10300 5414
rect 10356 5412 10380 5414
rect 10436 5412 10460 5414
rect 10516 5412 10522 5414
rect 10214 5392 10522 5412
rect 10214 4380 10522 4400
rect 10214 4378 10220 4380
rect 10276 4378 10300 4380
rect 10356 4378 10380 4380
rect 10436 4378 10460 4380
rect 10516 4378 10522 4380
rect 10276 4326 10278 4378
rect 10458 4326 10460 4378
rect 10214 4324 10220 4326
rect 10276 4324 10300 4326
rect 10356 4324 10380 4326
rect 10436 4324 10460 4326
rect 10516 4324 10522 4326
rect 10214 4304 10522 4324
rect 10214 3292 10522 3312
rect 10214 3290 10220 3292
rect 10276 3290 10300 3292
rect 10356 3290 10380 3292
rect 10436 3290 10460 3292
rect 10516 3290 10522 3292
rect 10276 3238 10278 3290
rect 10458 3238 10460 3290
rect 10214 3236 10220 3238
rect 10276 3236 10300 3238
rect 10356 3236 10380 3238
rect 10436 3236 10460 3238
rect 10516 3236 10522 3238
rect 10214 3216 10522 3236
rect 12360 3058 12388 5510
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12820 2774 12848 12582
rect 12912 12238 12940 12718
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 11694 12940 12038
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 13004 11150 13032 12242
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12992 10736 13044 10742
rect 12992 10678 13044 10684
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12912 9110 12940 9454
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12912 8566 12940 9046
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12912 8090 12940 8502
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12912 6866 12940 8026
rect 13004 7886 13032 10678
rect 13096 10266 13124 12838
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 13280 11234 13308 15116
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13452 15020 13504 15026
rect 13556 15008 13584 15150
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13636 15020 13688 15026
rect 13556 14980 13636 15008
rect 13452 14962 13504 14968
rect 13636 14962 13688 14968
rect 13740 15008 13768 15098
rect 13820 15020 13872 15026
rect 13740 14980 13820 15008
rect 13372 14414 13400 14962
rect 13464 14618 13492 14962
rect 13648 14822 13676 14962
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13372 14074 13400 14350
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13464 14074 13492 14282
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13372 11558 13400 13874
rect 13648 13870 13676 14758
rect 13740 13938 13768 14980
rect 13820 14962 13872 14968
rect 13820 14544 13872 14550
rect 13818 14512 13820 14521
rect 13872 14512 13874 14521
rect 13818 14447 13874 14456
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13924 13734 13952 17070
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 14016 15570 14044 16934
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 14004 14952 14056 14958
rect 14108 14929 14136 17682
rect 14292 17610 14320 18634
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14384 18086 14412 18566
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14280 17604 14332 17610
rect 14280 17546 14332 17552
rect 14292 17202 14320 17546
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 14200 15994 14228 16662
rect 14292 16114 14320 16934
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14200 15966 14320 15994
rect 14384 15978 14412 18022
rect 14476 16998 14504 19382
rect 14568 18970 14596 19722
rect 14752 19242 14780 19790
rect 14936 19514 14964 19790
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 14924 19372 14976 19378
rect 15028 19360 15056 19808
rect 15108 19790 15160 19796
rect 14976 19332 15056 19360
rect 14924 19314 14976 19320
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14752 18698 14780 19178
rect 14846 19068 15154 19088
rect 14846 19066 14852 19068
rect 14908 19066 14932 19068
rect 14988 19066 15012 19068
rect 15068 19066 15092 19068
rect 15148 19066 15154 19068
rect 14908 19014 14910 19066
rect 15090 19014 15092 19066
rect 14846 19012 14852 19014
rect 14908 19012 14932 19014
rect 14988 19012 15012 19014
rect 15068 19012 15092 19014
rect 15148 19012 15154 19014
rect 14846 18992 15154 19012
rect 15212 18834 15240 20198
rect 15396 19514 15424 26998
rect 17500 26920 17552 26926
rect 17500 26862 17552 26868
rect 17512 26382 17540 26862
rect 18064 26586 18092 27406
rect 20260 27328 20312 27334
rect 20260 27270 20312 27276
rect 19478 27228 19786 27248
rect 19478 27226 19484 27228
rect 19540 27226 19564 27228
rect 19620 27226 19644 27228
rect 19700 27226 19724 27228
rect 19780 27226 19786 27228
rect 19540 27174 19542 27226
rect 19722 27174 19724 27226
rect 19478 27172 19484 27174
rect 19540 27172 19564 27174
rect 19620 27172 19644 27174
rect 19700 27172 19724 27174
rect 19780 27172 19786 27174
rect 19478 27152 19786 27172
rect 19524 26852 19576 26858
rect 19524 26794 19576 26800
rect 19064 26784 19116 26790
rect 19340 26784 19392 26790
rect 19116 26732 19196 26738
rect 19064 26726 19196 26732
rect 19340 26726 19392 26732
rect 19076 26710 19196 26726
rect 18052 26580 18104 26586
rect 18052 26522 18104 26528
rect 18236 26580 18288 26586
rect 18236 26522 18288 26528
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 16672 26308 16724 26314
rect 16672 26250 16724 26256
rect 16684 26042 16712 26250
rect 17592 26240 17644 26246
rect 17592 26182 17644 26188
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 17316 26036 17368 26042
rect 17316 25978 17368 25984
rect 17328 25906 17356 25978
rect 15476 25900 15528 25906
rect 15476 25842 15528 25848
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17316 25900 17368 25906
rect 17316 25842 17368 25848
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17604 25888 17632 26182
rect 18248 26042 18276 26522
rect 18328 26308 18380 26314
rect 18328 26250 18380 26256
rect 18420 26308 18472 26314
rect 18420 26250 18472 26256
rect 18236 26036 18288 26042
rect 18236 25978 18288 25984
rect 18340 25922 18368 26250
rect 17684 25900 17736 25906
rect 17604 25860 17684 25888
rect 15488 24954 15516 25842
rect 17144 25498 17172 25842
rect 17224 25696 17276 25702
rect 17224 25638 17276 25644
rect 17236 25498 17264 25638
rect 17132 25492 17184 25498
rect 17132 25434 17184 25440
rect 17224 25492 17276 25498
rect 17224 25434 17276 25440
rect 16580 25424 16632 25430
rect 16580 25366 16632 25372
rect 16856 25424 16908 25430
rect 17328 25401 17356 25842
rect 16856 25366 16908 25372
rect 17314 25392 17370 25401
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 15476 24948 15528 24954
rect 15476 24890 15528 24896
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15488 24410 15516 24754
rect 16224 24750 16252 25094
rect 16302 24984 16358 24993
rect 16302 24919 16358 24928
rect 16316 24886 16344 24919
rect 16304 24880 16356 24886
rect 16304 24822 16356 24828
rect 16592 24818 16620 25366
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 16684 25158 16712 25230
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 15752 24744 15804 24750
rect 15752 24686 15804 24692
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 16212 24744 16264 24750
rect 16212 24686 16264 24692
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15660 24200 15712 24206
rect 15764 24177 15792 24686
rect 15660 24142 15712 24148
rect 15750 24168 15806 24177
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15488 23662 15516 24006
rect 15568 23724 15620 23730
rect 15672 23712 15700 24142
rect 15856 24138 15884 24686
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 16212 24268 16264 24274
rect 16212 24210 16264 24216
rect 15750 24103 15806 24112
rect 15844 24132 15896 24138
rect 15844 24074 15896 24080
rect 15752 23724 15804 23730
rect 15672 23684 15752 23712
rect 15568 23666 15620 23672
rect 15752 23666 15804 23672
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 15580 23322 15608 23666
rect 15568 23316 15620 23322
rect 15568 23258 15620 23264
rect 15764 23118 15792 23666
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15948 23118 15976 23462
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 16224 22778 16252 24210
rect 16500 23798 16528 24618
rect 16684 24410 16712 25094
rect 16868 24750 16896 25366
rect 17314 25327 17370 25336
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17420 24750 17448 25230
rect 17512 25158 17540 25842
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 16672 24404 16724 24410
rect 16672 24346 16724 24352
rect 17052 24206 17080 24550
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 17604 24138 17632 25860
rect 17684 25842 17736 25848
rect 18248 25894 18368 25922
rect 17776 24812 17828 24818
rect 17776 24754 17828 24760
rect 17788 24138 17816 24754
rect 18248 24342 18276 25894
rect 18328 25832 18380 25838
rect 18328 25774 18380 25780
rect 18340 25430 18368 25774
rect 18328 25424 18380 25430
rect 18328 25366 18380 25372
rect 18340 24750 18368 25366
rect 18432 24886 18460 26250
rect 18512 26036 18564 26042
rect 18512 25978 18564 25984
rect 18524 25362 18552 25978
rect 19168 25974 19196 26710
rect 19352 26382 19380 26726
rect 19536 26382 19564 26794
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19524 26376 19576 26382
rect 19524 26318 19576 26324
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 19156 25968 19208 25974
rect 19156 25910 19208 25916
rect 18696 25900 18748 25906
rect 18696 25842 18748 25848
rect 19064 25900 19116 25906
rect 19064 25842 19116 25848
rect 18708 25770 18736 25842
rect 18696 25764 18748 25770
rect 18696 25706 18748 25712
rect 18972 25764 19024 25770
rect 18972 25706 19024 25712
rect 18604 25696 18656 25702
rect 18984 25650 19012 25706
rect 18656 25644 19012 25650
rect 18604 25638 19012 25644
rect 18616 25622 19012 25638
rect 18512 25356 18564 25362
rect 18512 25298 18564 25304
rect 18420 24880 18472 24886
rect 18420 24822 18472 24828
rect 18328 24744 18380 24750
rect 18328 24686 18380 24692
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18432 24410 18460 24686
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18616 24410 18644 24550
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18604 24404 18656 24410
rect 18604 24346 18656 24352
rect 18236 24336 18288 24342
rect 18236 24278 18288 24284
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 16488 23792 16540 23798
rect 16488 23734 16540 23740
rect 16684 23730 16712 24074
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16684 23254 16712 23666
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16672 23248 16724 23254
rect 16672 23190 16724 23196
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16224 22030 16252 22714
rect 16396 22092 16448 22098
rect 16396 22034 16448 22040
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 15672 21622 15700 21830
rect 15660 21616 15712 21622
rect 15660 21558 15712 21564
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14568 17678 14596 18226
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14568 17270 14596 17614
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14568 16726 14596 17206
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14660 16969 14688 17138
rect 14646 16960 14702 16969
rect 14646 16895 14702 16904
rect 14556 16720 14608 16726
rect 14608 16668 14688 16674
rect 14556 16662 14688 16668
rect 14568 16646 14688 16662
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14004 14894 14056 14900
rect 14094 14920 14150 14929
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 14016 13410 14044 14894
rect 14094 14855 14150 14864
rect 14200 14482 14228 14962
rect 14292 14906 14320 15966
rect 14372 15972 14424 15978
rect 14372 15914 14424 15920
rect 14476 15502 14504 16050
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14384 15162 14412 15438
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 14370 15056 14426 15065
rect 14370 14991 14372 15000
rect 14424 14991 14426 15000
rect 14372 14962 14424 14968
rect 14292 14878 14412 14906
rect 14384 14822 14412 14878
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 14006 14136 14350
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 13924 13382 14044 13410
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13464 11626 13492 13194
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13464 11354 13492 11562
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13096 10062 13124 10202
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13188 9654 13216 11222
rect 13280 11206 13492 11234
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13280 10538 13308 11018
rect 13372 10606 13400 11086
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13280 10198 13308 10474
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13280 9654 13308 10134
rect 13464 9926 13492 11206
rect 13556 10742 13584 12106
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 11082 13768 11630
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13924 11014 13952 13382
rect 14004 13320 14056 13326
rect 14108 13274 14136 13738
rect 14056 13268 14136 13274
rect 14004 13262 14136 13268
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14016 13246 14136 13262
rect 14108 12850 14136 13246
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13464 9654 13492 9862
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8634 13124 8842
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13188 8362 13216 8978
rect 13464 8974 13492 9590
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13556 8974 13584 9318
rect 13832 9042 13860 9998
rect 13924 9994 13952 10950
rect 14016 10130 14044 12786
rect 14108 12646 14136 12786
rect 14200 12714 14228 13262
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14188 12436 14240 12442
rect 14292 12434 14320 14758
rect 14462 14512 14518 14521
rect 14462 14447 14464 14456
rect 14516 14447 14518 14456
rect 14464 14418 14516 14424
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14384 13394 14412 13806
rect 14476 13462 14504 13942
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14476 12850 14504 13398
rect 14568 12986 14596 16526
rect 14660 16114 14688 16646
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14648 15972 14700 15978
rect 14648 15914 14700 15920
rect 14660 14346 14688 15914
rect 14752 15162 14780 18226
rect 14846 17980 15154 18000
rect 14846 17978 14852 17980
rect 14908 17978 14932 17980
rect 14988 17978 15012 17980
rect 15068 17978 15092 17980
rect 15148 17978 15154 17980
rect 14908 17926 14910 17978
rect 15090 17926 15092 17978
rect 14846 17924 14852 17926
rect 14908 17924 14932 17926
rect 14988 17924 15012 17926
rect 15068 17924 15092 17926
rect 15148 17924 15154 17926
rect 14846 17904 15154 17924
rect 15212 17882 15240 18566
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14844 17338 14872 17682
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15120 17338 15148 17614
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 14846 16892 15154 16912
rect 14846 16890 14852 16892
rect 14908 16890 14932 16892
rect 14988 16890 15012 16892
rect 15068 16890 15092 16892
rect 15148 16890 15154 16892
rect 14908 16838 14910 16890
rect 15090 16838 15092 16890
rect 14846 16836 14852 16838
rect 14908 16836 14932 16838
rect 14988 16836 15012 16838
rect 15068 16836 15092 16838
rect 15148 16836 15154 16838
rect 14846 16816 15154 16836
rect 15304 16794 15332 19450
rect 15580 18426 15608 21286
rect 15764 21146 15792 21966
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 16408 20942 16436 22034
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16500 21350 16528 21830
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 15948 20602 15976 20878
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 16408 20466 16436 20878
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 16500 20398 16528 21286
rect 16868 20806 16896 23462
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17236 21078 17264 21354
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 16856 20800 16908 20806
rect 16856 20742 16908 20748
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 16212 20324 16264 20330
rect 16212 20266 16264 20272
rect 15842 19816 15898 19825
rect 15660 19780 15712 19786
rect 15842 19751 15844 19760
rect 15660 19722 15712 19728
rect 15896 19751 15898 19760
rect 15844 19722 15896 19728
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15396 18154 15424 18362
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15672 17882 15700 19722
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15764 18970 15792 19246
rect 16132 18970 16160 19314
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15764 18290 15792 18906
rect 16224 18834 16252 20266
rect 16304 19236 16356 19242
rect 16304 19178 16356 19184
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15566 17776 15622 17785
rect 15566 17711 15568 17720
rect 15620 17711 15622 17720
rect 15568 17682 15620 17688
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 15028 16182 15056 16458
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 14846 15804 15154 15824
rect 14846 15802 14852 15804
rect 14908 15802 14932 15804
rect 14988 15802 15012 15804
rect 15068 15802 15092 15804
rect 15148 15802 15154 15804
rect 14908 15750 14910 15802
rect 15090 15750 15092 15802
rect 14846 15748 14852 15750
rect 14908 15748 14932 15750
rect 14988 15748 15012 15750
rect 15068 15748 15092 15750
rect 15148 15748 15154 15750
rect 14846 15728 15154 15748
rect 15212 15570 15240 16390
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15304 15502 15332 15846
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14738 15056 14794 15065
rect 15212 15026 15240 15370
rect 14738 14991 14794 15000
rect 15200 15020 15252 15026
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14646 13832 14702 13841
rect 14646 13767 14702 13776
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14660 12850 14688 13767
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14752 12434 14780 14991
rect 15200 14962 15252 14968
rect 14846 14716 15154 14736
rect 14846 14714 14852 14716
rect 14908 14714 14932 14716
rect 14988 14714 15012 14716
rect 15068 14714 15092 14716
rect 15148 14714 15154 14716
rect 14908 14662 14910 14714
rect 15090 14662 15092 14714
rect 14846 14660 14852 14662
rect 14908 14660 14932 14662
rect 14988 14660 15012 14662
rect 15068 14660 15092 14662
rect 15148 14660 15154 14662
rect 14846 14640 15154 14660
rect 15212 14414 15240 14962
rect 15396 14958 15424 15438
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 14550 15332 14758
rect 15396 14550 15424 14894
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15290 14376 15346 14385
rect 15290 14311 15346 14320
rect 15304 14278 15332 14311
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15304 13734 15332 14214
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 14846 13628 15154 13648
rect 14846 13626 14852 13628
rect 14908 13626 14932 13628
rect 14988 13626 15012 13628
rect 15068 13626 15092 13628
rect 15148 13626 15154 13628
rect 14908 13574 14910 13626
rect 15090 13574 15092 13626
rect 14846 13572 14852 13574
rect 14908 13572 14932 13574
rect 14988 13572 15012 13574
rect 15068 13572 15092 13574
rect 15148 13572 15154 13574
rect 14846 13552 15154 13572
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14844 12918 14872 13126
rect 15488 12986 15516 17138
rect 15764 16454 15792 17206
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15764 16114 15792 16390
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15672 15162 15700 15370
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 15672 12764 15700 15098
rect 15856 13530 15884 17614
rect 15948 17542 15976 18634
rect 16132 18426 16160 18702
rect 16316 18698 16344 19178
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 16028 18352 16080 18358
rect 16028 18294 16080 18300
rect 16040 17542 16068 18294
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 16040 16114 16068 17478
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15948 14414 15976 15506
rect 16132 14482 16160 18362
rect 16408 17814 16436 18566
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16224 17202 16252 17614
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16794 16252 16934
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16224 15706 16252 16730
rect 16304 16720 16356 16726
rect 16304 16662 16356 16668
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15948 14006 15976 14350
rect 15936 14000 15988 14006
rect 15936 13942 15988 13948
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15948 13394 15976 13942
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15752 12776 15804 12782
rect 15672 12736 15752 12764
rect 15752 12718 15804 12724
rect 15108 12708 15160 12714
rect 15160 12668 15240 12696
rect 15108 12650 15160 12656
rect 14846 12540 15154 12560
rect 14846 12538 14852 12540
rect 14908 12538 14932 12540
rect 14988 12538 15012 12540
rect 15068 12538 15092 12540
rect 15148 12538 15154 12540
rect 14908 12486 14910 12538
rect 15090 12486 15092 12538
rect 14846 12484 14852 12486
rect 14908 12484 14932 12486
rect 14988 12484 15012 12486
rect 15068 12484 15092 12486
rect 15148 12484 15154 12486
rect 14846 12464 15154 12484
rect 15212 12434 15240 12668
rect 15948 12646 15976 13330
rect 16224 13258 16252 13942
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16040 12782 16068 13126
rect 16224 12850 16252 13194
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 14292 12406 14412 12434
rect 14188 12378 14240 12384
rect 14200 11762 14228 12378
rect 14278 12336 14334 12345
rect 14278 12271 14334 12280
rect 14292 12238 14320 12271
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14292 11150 14320 11494
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14200 10266 14228 11086
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14292 10062 14320 10610
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13280 7410 13308 8230
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 13372 6662 13400 8366
rect 13464 8090 13492 8910
rect 13634 8664 13690 8673
rect 14200 8634 14228 9998
rect 14292 9722 14320 9998
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14384 9058 14412 12406
rect 14660 12406 14780 12434
rect 15120 12406 15240 12434
rect 14660 12170 14688 12406
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14568 11354 14596 11698
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14292 9030 14412 9058
rect 13634 8599 13636 8608
rect 13688 8599 13690 8608
rect 14188 8628 14240 8634
rect 13636 8570 13688 8576
rect 14188 8570 14240 8576
rect 13648 8378 13676 8570
rect 14292 8498 14320 9030
rect 14476 8974 14504 11290
rect 14660 11098 14688 12106
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11218 14780 12038
rect 15120 11540 15148 12406
rect 16040 12238 16068 12718
rect 16224 12646 16252 12786
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16118 12200 16174 12209
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15120 11512 15240 11540
rect 14846 11452 15154 11472
rect 14846 11450 14852 11452
rect 14908 11450 14932 11452
rect 14988 11450 15012 11452
rect 15068 11450 15092 11452
rect 15148 11450 15154 11452
rect 14908 11398 14910 11450
rect 15090 11398 15092 11450
rect 14846 11396 14852 11398
rect 14908 11396 14932 11398
rect 14988 11396 15012 11398
rect 15068 11396 15092 11398
rect 15148 11396 15154 11398
rect 14846 11376 15154 11396
rect 15212 11336 15240 11512
rect 15120 11308 15240 11336
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14660 11070 14780 11098
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14660 9926 14688 10950
rect 14752 10674 14780 11070
rect 15120 11014 15148 11308
rect 15672 11150 15700 11834
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14846 10364 15154 10384
rect 14846 10362 14852 10364
rect 14908 10362 14932 10364
rect 14988 10362 15012 10364
rect 15068 10362 15092 10364
rect 15148 10362 15154 10364
rect 14908 10310 14910 10362
rect 15090 10310 15092 10362
rect 14846 10308 14852 10310
rect 14908 10308 14932 10310
rect 14988 10308 15012 10310
rect 15068 10308 15092 10310
rect 15148 10308 15154 10310
rect 14846 10288 15154 10308
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 15212 9518 15240 11018
rect 15304 10266 15332 11086
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15396 10062 15424 10406
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 14846 9276 15154 9296
rect 14846 9274 14852 9276
rect 14908 9274 14932 9276
rect 14988 9274 15012 9276
rect 15068 9274 15092 9276
rect 15148 9274 15154 9276
rect 14908 9222 14910 9274
rect 15090 9222 15092 9274
rect 14846 9220 14852 9222
rect 14908 9220 14932 9222
rect 14988 9220 15012 9222
rect 15068 9220 15092 9222
rect 15148 9220 15154 9222
rect 14846 9200 15154 9220
rect 15212 9178 15240 9454
rect 15488 9450 15516 10678
rect 15764 10606 15792 11086
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 10266 15608 10474
rect 15764 10266 15792 10542
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15568 9648 15620 9654
rect 15566 9616 15568 9625
rect 15752 9648 15804 9654
rect 15620 9616 15752 9636
rect 15622 9608 15752 9616
rect 15752 9590 15804 9596
rect 15566 9551 15622 9560
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 14384 8634 14412 8842
rect 14568 8634 14596 9114
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14936 8498 14964 8774
rect 15488 8566 15516 9386
rect 15856 8974 15884 12174
rect 16118 12135 16174 12144
rect 16132 11762 16160 12135
rect 16316 11801 16344 16662
rect 16408 15434 16436 17614
rect 16500 17610 16528 20334
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16592 15586 16620 18770
rect 16684 18630 16712 20198
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16854 18456 16910 18465
rect 16854 18391 16856 18400
rect 16908 18391 16910 18400
rect 16856 18362 16908 18368
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16684 17338 16712 18226
rect 16960 18222 16988 20402
rect 17144 20058 17172 20742
rect 17236 20398 17264 21014
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 17052 18970 17080 19722
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 17144 18306 17172 19994
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17236 18766 17264 19382
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17328 18426 17356 19314
rect 17420 18426 17448 22034
rect 17604 22030 17632 24074
rect 17788 22642 17816 24074
rect 18432 23730 18460 24074
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18156 23322 18184 23666
rect 18524 23322 18552 24142
rect 18984 24138 19012 25622
rect 19076 25430 19104 25842
rect 19168 25838 19196 25910
rect 19156 25832 19208 25838
rect 19156 25774 19208 25780
rect 19064 25424 19116 25430
rect 19064 25366 19116 25372
rect 19064 25152 19116 25158
rect 19064 25094 19116 25100
rect 19076 24954 19104 25094
rect 19168 24954 19196 25774
rect 19248 25152 19300 25158
rect 19248 25094 19300 25100
rect 19064 24948 19116 24954
rect 19064 24890 19116 24896
rect 19156 24948 19208 24954
rect 19156 24890 19208 24896
rect 19076 24614 19104 24890
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 19260 24206 19288 25094
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 18972 24132 19024 24138
rect 18972 24074 19024 24080
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 18512 23316 18564 23322
rect 18512 23258 18564 23264
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17776 22092 17828 22098
rect 17776 22034 17828 22040
rect 18052 22092 18104 22098
rect 18052 22034 18104 22040
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 17592 21344 17644 21350
rect 17592 21286 17644 21292
rect 17604 20942 17632 21286
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17512 19854 17540 20878
rect 17788 20058 17816 22034
rect 18064 21554 18092 22034
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 17972 20602 18000 21490
rect 18328 20868 18380 20874
rect 18328 20810 18380 20816
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 18340 20466 18368 20810
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17512 19514 17540 19790
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17512 18834 17540 19450
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17144 18278 17356 18306
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16776 16590 16804 18022
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16868 15638 16896 17546
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16960 15638 16988 15846
rect 16856 15632 16908 15638
rect 16592 15558 16712 15586
rect 16856 15574 16908 15580
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16396 15428 16448 15434
rect 16396 15370 16448 15376
rect 16592 14890 16620 15438
rect 16684 15162 16712 15558
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16776 15026 16804 15302
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 16592 14482 16620 14826
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16776 13938 16804 14962
rect 16868 14414 16896 15370
rect 17052 15026 17080 17546
rect 17144 17270 17172 18022
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17236 16726 17264 17546
rect 17328 17218 17356 18278
rect 17420 17338 17448 18362
rect 17512 17882 17540 18770
rect 17604 18766 17632 19110
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17696 18426 17724 19110
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17590 18320 17646 18329
rect 17590 18255 17592 18264
rect 17644 18255 17646 18264
rect 17592 18226 17644 18232
rect 17880 18222 17908 19314
rect 18340 19310 18368 20402
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18432 19961 18460 20198
rect 18418 19952 18474 19961
rect 18418 19887 18474 19896
rect 18432 19854 18460 19887
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18524 18222 18552 23122
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18616 22778 18644 22918
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 18708 20806 18736 21490
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 20534 18736 20742
rect 18696 20528 18748 20534
rect 18696 20470 18748 20476
rect 18800 20346 18828 23258
rect 18984 23118 19012 24074
rect 19352 23798 19380 26318
rect 19892 26308 19944 26314
rect 19892 26250 19944 26256
rect 19478 26140 19786 26160
rect 19478 26138 19484 26140
rect 19540 26138 19564 26140
rect 19620 26138 19644 26140
rect 19700 26138 19724 26140
rect 19780 26138 19786 26140
rect 19540 26086 19542 26138
rect 19722 26086 19724 26138
rect 19478 26084 19484 26086
rect 19540 26084 19564 26086
rect 19620 26084 19644 26086
rect 19700 26084 19724 26086
rect 19780 26084 19786 26086
rect 19478 26064 19786 26084
rect 19524 25696 19576 25702
rect 19524 25638 19576 25644
rect 19536 25294 19564 25638
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19478 25052 19786 25072
rect 19478 25050 19484 25052
rect 19540 25050 19564 25052
rect 19620 25050 19644 25052
rect 19700 25050 19724 25052
rect 19780 25050 19786 25052
rect 19540 24998 19542 25050
rect 19722 24998 19724 25050
rect 19478 24996 19484 24998
rect 19540 24996 19564 24998
rect 19620 24996 19644 24998
rect 19700 24996 19724 24998
rect 19780 24996 19786 24998
rect 19478 24976 19786 24996
rect 19708 24812 19760 24818
rect 19708 24754 19760 24760
rect 19720 24274 19748 24754
rect 19904 24682 19932 26250
rect 19996 25838 20024 26318
rect 20272 26314 20300 27270
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20456 26586 20484 26930
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20260 26308 20312 26314
rect 20260 26250 20312 26256
rect 20260 26036 20312 26042
rect 20260 25978 20312 25984
rect 20272 25838 20300 25978
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 20260 25832 20312 25838
rect 20260 25774 20312 25780
rect 20168 25220 20220 25226
rect 20168 25162 20220 25168
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 19892 24676 19944 24682
rect 19892 24618 19944 24624
rect 19708 24268 19760 24274
rect 19708 24210 19760 24216
rect 19478 23964 19786 23984
rect 19478 23962 19484 23964
rect 19540 23962 19564 23964
rect 19620 23962 19644 23964
rect 19700 23962 19724 23964
rect 19780 23962 19786 23964
rect 19540 23910 19542 23962
rect 19722 23910 19724 23962
rect 19478 23908 19484 23910
rect 19540 23908 19564 23910
rect 19620 23908 19644 23910
rect 19700 23908 19724 23910
rect 19780 23908 19786 23910
rect 19478 23888 19786 23908
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19904 23610 19932 24618
rect 19996 23730 20024 24890
rect 20180 24886 20208 25162
rect 20168 24880 20220 24886
rect 20168 24822 20220 24828
rect 20272 24410 20300 25774
rect 20640 25770 20668 27406
rect 20996 27396 21048 27402
rect 20996 27338 21048 27344
rect 21008 26382 21036 27338
rect 20996 26376 21048 26382
rect 20996 26318 21048 26324
rect 20720 25968 20772 25974
rect 20720 25910 20772 25916
rect 20536 25764 20588 25770
rect 20536 25706 20588 25712
rect 20628 25764 20680 25770
rect 20628 25706 20680 25712
rect 20352 25220 20404 25226
rect 20352 25162 20404 25168
rect 20364 24750 20392 25162
rect 20548 24818 20576 25706
rect 20640 24818 20668 25706
rect 20732 25362 20760 25910
rect 21008 25906 21036 26318
rect 21100 26246 21128 27474
rect 23860 27130 23888 29200
rect 24110 27772 24418 27792
rect 24110 27770 24116 27772
rect 24172 27770 24196 27772
rect 24252 27770 24276 27772
rect 24332 27770 24356 27772
rect 24412 27770 24418 27772
rect 24172 27718 24174 27770
rect 24354 27718 24356 27770
rect 24110 27716 24116 27718
rect 24172 27716 24196 27718
rect 24252 27716 24276 27718
rect 24332 27716 24356 27718
rect 24412 27716 24418 27718
rect 24110 27696 24418 27716
rect 25148 27606 25176 29200
rect 26528 27606 26556 29294
rect 27710 29294 28120 29322
rect 27710 29200 27766 29294
rect 27526 28656 27582 28665
rect 27526 28591 27582 28600
rect 25136 27600 25188 27606
rect 25136 27542 25188 27548
rect 26516 27600 26568 27606
rect 26516 27542 26568 27548
rect 25872 27396 25924 27402
rect 25872 27338 25924 27344
rect 23848 27124 23900 27130
rect 23848 27066 23900 27072
rect 21732 26988 21784 26994
rect 21732 26930 21784 26936
rect 25504 26988 25556 26994
rect 25504 26930 25556 26936
rect 21744 26518 21772 26930
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 21732 26512 21784 26518
rect 21732 26454 21784 26460
rect 22204 26382 22232 26726
rect 22192 26376 22244 26382
rect 22192 26318 22244 26324
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 21916 26240 21968 26246
rect 21916 26182 21968 26188
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 20720 25356 20772 25362
rect 20720 25298 20772 25304
rect 20904 25288 20956 25294
rect 21008 25276 21036 25842
rect 21100 25838 21128 26182
rect 21928 26042 21956 26182
rect 21456 26036 21508 26042
rect 21456 25978 21508 25984
rect 21916 26036 21968 26042
rect 21916 25978 21968 25984
rect 21088 25832 21140 25838
rect 21088 25774 21140 25780
rect 21086 25392 21142 25401
rect 21086 25327 21142 25336
rect 21100 25294 21128 25327
rect 21468 25294 21496 25978
rect 22204 25974 22232 26318
rect 22192 25968 22244 25974
rect 22192 25910 22244 25916
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22112 25770 22140 25842
rect 22100 25764 22152 25770
rect 22100 25706 22152 25712
rect 22008 25424 22060 25430
rect 22008 25366 22060 25372
rect 20956 25248 21036 25276
rect 21088 25288 21140 25294
rect 20904 25230 20956 25236
rect 21088 25230 21140 25236
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 20916 24954 20944 25230
rect 20904 24948 20956 24954
rect 20904 24890 20956 24896
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20352 24744 20404 24750
rect 20352 24686 20404 24692
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20260 24404 20312 24410
rect 20260 24346 20312 24352
rect 20456 24342 20484 24550
rect 21100 24410 21128 25230
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 21284 24954 21312 25094
rect 21272 24948 21324 24954
rect 21272 24890 21324 24896
rect 22020 24614 22048 25366
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 21088 24404 21140 24410
rect 21088 24346 21140 24352
rect 20444 24336 20496 24342
rect 20444 24278 20496 24284
rect 20260 24200 20312 24206
rect 20260 24142 20312 24148
rect 20352 24200 20404 24206
rect 20904 24200 20956 24206
rect 20352 24142 20404 24148
rect 20718 24168 20774 24177
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19904 23582 20208 23610
rect 20272 23594 20300 24142
rect 20364 23866 20392 24142
rect 20718 24103 20774 24112
rect 20824 24160 20904 24188
rect 20352 23860 20404 23866
rect 20352 23802 20404 23808
rect 20364 23594 20392 23802
rect 20732 23798 20760 24103
rect 20444 23792 20496 23798
rect 20444 23734 20496 23740
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19984 23248 20036 23254
rect 19984 23190 20036 23196
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 19892 22976 19944 22982
rect 19892 22918 19944 22924
rect 19478 22876 19786 22896
rect 19478 22874 19484 22876
rect 19540 22874 19564 22876
rect 19620 22874 19644 22876
rect 19700 22874 19724 22876
rect 19780 22874 19786 22876
rect 19540 22822 19542 22874
rect 19722 22822 19724 22874
rect 19478 22820 19484 22822
rect 19540 22820 19564 22822
rect 19620 22820 19644 22822
rect 19700 22820 19724 22822
rect 19780 22820 19786 22822
rect 19478 22800 19786 22820
rect 19904 22778 19932 22918
rect 19892 22772 19944 22778
rect 19892 22714 19944 22720
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19064 22160 19116 22166
rect 19064 22102 19116 22108
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18892 21486 18920 21966
rect 19076 21554 19104 22102
rect 19352 21894 19380 22510
rect 19892 22500 19944 22506
rect 19892 22442 19944 22448
rect 19904 21978 19932 22442
rect 19996 22166 20024 23190
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19904 21950 20024 21978
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 19478 21788 19786 21808
rect 19478 21786 19484 21788
rect 19540 21786 19564 21788
rect 19620 21786 19644 21788
rect 19700 21786 19724 21788
rect 19780 21786 19786 21788
rect 19540 21734 19542 21786
rect 19722 21734 19724 21786
rect 19478 21732 19484 21734
rect 19540 21732 19564 21734
rect 19620 21732 19644 21734
rect 19700 21732 19724 21734
rect 19780 21732 19786 21734
rect 19478 21712 19786 21732
rect 19904 21690 19932 21830
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18878 20496 18934 20505
rect 18878 20431 18934 20440
rect 19064 20460 19116 20466
rect 18708 20318 18828 20346
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18616 19378 18644 19790
rect 18708 19718 18736 20318
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18800 19378 18828 20198
rect 18892 19961 18920 20431
rect 19064 20402 19116 20408
rect 18878 19952 18934 19961
rect 18878 19887 18934 19896
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18892 19122 18920 19887
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18984 19242 19012 19790
rect 18972 19236 19024 19242
rect 18972 19178 19024 19184
rect 18892 19094 19012 19122
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17328 17190 17448 17218
rect 17224 16720 17276 16726
rect 17130 16688 17186 16697
rect 17224 16662 17276 16668
rect 17130 16623 17186 16632
rect 17144 16153 17172 16623
rect 17130 16144 17186 16153
rect 17130 16079 17132 16088
rect 17184 16079 17186 16088
rect 17132 16050 17184 16056
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17328 15502 17356 15846
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17420 15434 17448 17190
rect 17512 16658 17540 17818
rect 17776 17128 17828 17134
rect 17880 17116 17908 18158
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 17958 17232 18014 17241
rect 17958 17167 17960 17176
rect 18012 17167 18014 17176
rect 17960 17138 18012 17144
rect 17828 17088 17908 17116
rect 17776 17070 17828 17076
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17880 16266 17908 17088
rect 17958 16416 18014 16425
rect 17958 16351 18014 16360
rect 17696 16250 17908 16266
rect 17696 16244 17920 16250
rect 17696 16238 17868 16244
rect 17696 16182 17724 16238
rect 17868 16186 17920 16192
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 17236 15008 17264 15370
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17316 15020 17368 15026
rect 17236 14980 17316 15008
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16592 13462 16620 13738
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16592 12986 16620 13398
rect 16776 13394 16804 13874
rect 17052 13870 17080 14962
rect 17236 14618 17264 14980
rect 17316 14962 17368 14968
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17144 13734 17172 14214
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 13530 17172 13670
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 17144 13326 17172 13466
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16408 11898 16436 12378
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16592 11830 16620 12174
rect 16684 11898 16712 12786
rect 16960 12434 16988 12854
rect 16868 12406 16988 12434
rect 16868 12238 16896 12406
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16580 11824 16632 11830
rect 16302 11792 16358 11801
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16212 11756 16264 11762
rect 16580 11766 16632 11772
rect 16302 11727 16358 11736
rect 16212 11698 16264 11704
rect 16224 11626 16252 11698
rect 16212 11620 16264 11626
rect 16212 11562 16264 11568
rect 16224 11286 16252 11562
rect 16212 11280 16264 11286
rect 16210 11248 16212 11257
rect 16264 11248 16266 11257
rect 16210 11183 16266 11192
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 13648 8350 13860 8378
rect 13832 8090 13860 8350
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 14292 7818 14320 8434
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14476 7410 14504 8298
rect 14568 8090 14596 8434
rect 15382 8392 15438 8401
rect 15382 8327 15438 8336
rect 14846 8188 15154 8208
rect 14846 8186 14852 8188
rect 14908 8186 14932 8188
rect 14988 8186 15012 8188
rect 15068 8186 15092 8188
rect 15148 8186 15154 8188
rect 14908 8134 14910 8186
rect 15090 8134 15092 8186
rect 14846 8132 14852 8134
rect 14908 8132 14932 8134
rect 14988 8132 15012 8134
rect 15068 8132 15092 8134
rect 15148 8132 15154 8134
rect 14846 8112 15154 8132
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13450 6896 13506 6905
rect 13450 6831 13506 6840
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13464 5710 13492 6831
rect 13556 6798 13584 7142
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13740 5778 13768 6802
rect 14200 6186 14228 7346
rect 14476 6662 14504 7346
rect 14568 7342 14596 8026
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14844 7478 14872 7686
rect 15120 7546 15148 7822
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 15396 7410 15424 8327
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 15488 7274 15516 8502
rect 15856 8430 15884 8910
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15476 7268 15528 7274
rect 15476 7210 15528 7216
rect 14846 7100 15154 7120
rect 14846 7098 14852 7100
rect 14908 7098 14932 7100
rect 14988 7098 15012 7100
rect 15068 7098 15092 7100
rect 15148 7098 15154 7100
rect 14908 7046 14910 7098
rect 15090 7046 15092 7098
rect 14846 7044 14852 7046
rect 14908 7044 14932 7046
rect 14988 7044 15012 7046
rect 15068 7044 15092 7046
rect 15148 7044 15154 7046
rect 14846 7024 15154 7044
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15856 6186 15884 6598
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 14846 6012 15154 6032
rect 14846 6010 14852 6012
rect 14908 6010 14932 6012
rect 14988 6010 15012 6012
rect 15068 6010 15092 6012
rect 15148 6010 15154 6012
rect 14908 5958 14910 6010
rect 15090 5958 15092 6010
rect 14846 5956 14852 5958
rect 14908 5956 14932 5958
rect 14988 5956 15012 5958
rect 15068 5956 15092 5958
rect 15148 5956 15154 5958
rect 14846 5936 15154 5956
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 15672 5642 15700 6054
rect 15660 5636 15712 5642
rect 15660 5578 15712 5584
rect 14846 4924 15154 4944
rect 14846 4922 14852 4924
rect 14908 4922 14932 4924
rect 14988 4922 15012 4924
rect 15068 4922 15092 4924
rect 15148 4922 15154 4924
rect 14908 4870 14910 4922
rect 15090 4870 15092 4922
rect 14846 4868 14852 4870
rect 14908 4868 14932 4870
rect 14988 4868 15012 4870
rect 15068 4868 15092 4870
rect 15148 4868 15154 4870
rect 14846 4848 15154 4868
rect 14846 3836 15154 3856
rect 14846 3834 14852 3836
rect 14908 3834 14932 3836
rect 14988 3834 15012 3836
rect 15068 3834 15092 3836
rect 15148 3834 15154 3836
rect 14908 3782 14910 3834
rect 15090 3782 15092 3834
rect 14846 3780 14852 3782
rect 14908 3780 14932 3782
rect 14988 3780 15012 3782
rect 15068 3780 15092 3782
rect 15148 3780 15154 3782
rect 14846 3760 15154 3780
rect 12636 2746 12848 2774
rect 14846 2748 15154 2768
rect 14846 2746 14852 2748
rect 14908 2746 14932 2748
rect 14988 2746 15012 2748
rect 15068 2746 15092 2748
rect 15148 2746 15154 2748
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 1492 2304 1544 2310
rect 1492 2246 1544 2252
rect 1504 1465 1532 2246
rect 1490 1456 1546 1465
rect 1490 1391 1546 1400
rect 2608 800 2636 2382
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 800 5212 2246
rect 6472 800 6500 2382
rect 7760 800 7788 2382
rect 10152 1306 10180 2382
rect 12636 2378 12664 2746
rect 14908 2694 14910 2746
rect 15090 2694 15092 2746
rect 14846 2692 14852 2694
rect 14908 2692 14932 2694
rect 14988 2692 15012 2694
rect 15068 2692 15092 2694
rect 15148 2692 15154 2694
rect 14846 2672 15154 2692
rect 15856 2650 15884 6122
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15948 2582 15976 10950
rect 16316 10810 16344 11727
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16224 9586 16252 10066
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16040 6390 16068 8366
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16224 7546 16252 7754
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16132 6322 16160 6598
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16592 3194 16620 11766
rect 17132 11688 17184 11694
rect 17130 11656 17132 11665
rect 17184 11656 17186 11665
rect 17130 11591 17186 11600
rect 17144 11286 17172 11591
rect 17236 11354 17264 14554
rect 17604 14414 17632 15302
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17512 14006 17540 14282
rect 17500 14000 17552 14006
rect 17696 13977 17724 15982
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17788 14958 17816 15642
rect 17880 15570 17908 15914
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17880 15162 17908 15506
rect 17972 15473 18000 16351
rect 17958 15464 18014 15473
rect 17958 15399 17960 15408
rect 18012 15399 18014 15408
rect 17960 15370 18012 15376
rect 17972 15339 18000 15370
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17500 13942 17552 13948
rect 17682 13968 17738 13977
rect 17682 13903 17738 13912
rect 17788 12850 17816 14894
rect 18248 13852 18276 18022
rect 18524 17882 18552 18158
rect 18892 18086 18920 18226
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18602 17640 18658 17649
rect 18602 17575 18658 17584
rect 18616 17542 18644 17575
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 16425 18644 17478
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18602 16416 18658 16425
rect 18602 16351 18658 16360
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18616 15026 18644 15302
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18340 14006 18368 14894
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18432 14074 18460 14486
rect 18524 14414 18552 14758
rect 18708 14414 18736 16934
rect 18788 16516 18840 16522
rect 18788 16458 18840 16464
rect 18800 16250 18828 16458
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18892 16153 18920 16934
rect 18878 16144 18934 16153
rect 18878 16079 18934 16088
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18800 14618 18828 15438
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18512 14408 18564 14414
rect 18696 14408 18748 14414
rect 18512 14350 18564 14356
rect 18616 14376 18696 14396
rect 18748 14376 18750 14385
rect 18616 14368 18694 14376
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18248 13824 18368 13852
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17788 12238 17816 12786
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17880 12102 17908 12922
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17972 12170 18000 12718
rect 18064 12646 18092 13126
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18064 12306 18092 12582
rect 18156 12442 18184 12650
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17788 11694 17816 12038
rect 17880 11762 17908 12038
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17420 11082 17448 11630
rect 17880 11218 17908 11698
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17972 11082 18000 12106
rect 18248 11830 18276 12582
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18248 11150 18276 11766
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16868 10062 16896 10746
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17328 10062 17356 10406
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 8673 16712 9318
rect 17052 9178 17080 9522
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16670 8664 16726 8673
rect 16868 8634 16896 8910
rect 17328 8634 17356 9114
rect 16670 8599 16726 8608
rect 16856 8628 16908 8634
rect 16684 8430 16712 8599
rect 16856 8570 16908 8576
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16776 7410 16804 8298
rect 17040 7812 17092 7818
rect 17040 7754 17092 7760
rect 17052 7546 17080 7754
rect 17144 7546 17172 8434
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 16868 5846 16896 6598
rect 17052 6322 17080 6598
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 17420 3194 17448 11018
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17696 10266 17724 10610
rect 18340 10538 18368 13824
rect 18432 13394 18460 13874
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18524 13258 18552 14350
rect 18616 13530 18644 14368
rect 18694 14311 18750 14320
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18524 12442 18552 13194
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18616 11354 18644 13466
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18604 11076 18656 11082
rect 18604 11018 18656 11024
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17972 9994 18000 10406
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 18064 9926 18092 10406
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 8906 17540 9318
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17880 8838 17908 9386
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17776 7880 17828 7886
rect 17880 7868 17908 8774
rect 17828 7840 17908 7868
rect 17776 7822 17828 7828
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17696 7546 17724 7686
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17880 7478 17908 7840
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17604 6866 17632 7346
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17604 6458 17632 6802
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17512 5710 17540 6258
rect 17696 5914 17724 6734
rect 17880 6390 17908 7414
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17972 5574 18000 9590
rect 18142 8936 18198 8945
rect 18142 8871 18198 8880
rect 18156 8838 18184 8871
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17972 5370 18000 5510
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 15936 2576 15988 2582
rect 15936 2518 15988 2524
rect 17328 2514 17356 2994
rect 18064 2650 18092 8434
rect 18156 8430 18184 8774
rect 18248 8566 18276 10066
rect 18340 8906 18368 10474
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18432 9586 18460 9930
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18524 8634 18552 11018
rect 18616 10742 18644 11018
rect 18604 10736 18656 10742
rect 18604 10678 18656 10684
rect 18616 9586 18644 10678
rect 18800 10130 18828 11494
rect 18892 10452 18920 16079
rect 18984 14396 19012 19094
rect 19076 18154 19104 20402
rect 19168 20262 19196 21490
rect 19524 21480 19576 21486
rect 19524 21422 19576 21428
rect 19536 21078 19564 21422
rect 19892 21412 19944 21418
rect 19892 21354 19944 21360
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 19536 20942 19564 21014
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19478 20700 19786 20720
rect 19478 20698 19484 20700
rect 19540 20698 19564 20700
rect 19620 20698 19644 20700
rect 19700 20698 19724 20700
rect 19780 20698 19786 20700
rect 19540 20646 19542 20698
rect 19722 20646 19724 20698
rect 19478 20644 19484 20646
rect 19540 20644 19564 20646
rect 19620 20644 19644 20646
rect 19700 20644 19724 20646
rect 19780 20644 19786 20646
rect 19478 20624 19786 20644
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19248 20324 19300 20330
rect 19248 20266 19300 20272
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19260 19922 19288 20266
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 19168 19378 19196 19654
rect 19260 19514 19288 19858
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19352 19446 19380 20470
rect 19904 19854 19932 21354
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19996 19700 20024 21950
rect 20088 21554 20116 23462
rect 20180 22642 20208 23582
rect 20260 23588 20312 23594
rect 20260 23530 20312 23536
rect 20352 23588 20404 23594
rect 20352 23530 20404 23536
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 20272 22094 20300 23530
rect 20456 23118 20484 23734
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20548 23322 20576 23666
rect 20824 23594 20852 24160
rect 20904 24142 20956 24148
rect 21100 24052 21128 24346
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 20916 24024 21128 24052
rect 20812 23588 20864 23594
rect 20812 23530 20864 23536
rect 20536 23316 20588 23322
rect 20588 23276 20668 23304
rect 20536 23258 20588 23264
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20180 22066 20300 22094
rect 20180 21622 20208 22066
rect 20456 22030 20484 23054
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20444 22024 20496 22030
rect 20444 21966 20496 21972
rect 20168 21616 20220 21622
rect 20168 21558 20220 21564
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 20076 21072 20128 21078
rect 20076 21014 20128 21020
rect 20088 20806 20116 21014
rect 20272 21010 20300 21558
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20364 21146 20392 21490
rect 20456 21486 20484 21966
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20260 21004 20312 21010
rect 20260 20946 20312 20952
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 19904 19672 20024 19700
rect 19478 19612 19786 19632
rect 19478 19610 19484 19612
rect 19540 19610 19564 19612
rect 19620 19610 19644 19612
rect 19700 19610 19724 19612
rect 19780 19610 19786 19612
rect 19540 19558 19542 19610
rect 19722 19558 19724 19610
rect 19478 19556 19484 19558
rect 19540 19556 19564 19558
rect 19620 19556 19644 19558
rect 19700 19556 19724 19558
rect 19780 19556 19786 19558
rect 19478 19536 19786 19556
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 19168 14550 19196 19314
rect 19536 18970 19564 19314
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19260 18358 19288 18634
rect 19248 18352 19300 18358
rect 19248 18294 19300 18300
rect 19260 17898 19288 18294
rect 19352 18086 19380 18906
rect 19478 18524 19786 18544
rect 19478 18522 19484 18524
rect 19540 18522 19564 18524
rect 19620 18522 19644 18524
rect 19700 18522 19724 18524
rect 19780 18522 19786 18524
rect 19540 18470 19542 18522
rect 19722 18470 19724 18522
rect 19478 18468 19484 18470
rect 19540 18468 19564 18470
rect 19620 18468 19644 18470
rect 19700 18468 19724 18470
rect 19780 18468 19786 18470
rect 19478 18448 19786 18468
rect 19904 18290 19932 19672
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19996 18902 20024 19246
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19996 18465 20024 18702
rect 19982 18456 20038 18465
rect 19982 18391 20038 18400
rect 19892 18284 19944 18290
rect 19944 18244 20024 18272
rect 19892 18226 19944 18232
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19260 17870 19380 17898
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19260 16658 19288 17546
rect 19352 17202 19380 17870
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19478 17436 19786 17456
rect 19478 17434 19484 17436
rect 19540 17434 19564 17436
rect 19620 17434 19644 17436
rect 19700 17434 19724 17436
rect 19780 17434 19786 17436
rect 19540 17382 19542 17434
rect 19722 17382 19724 17434
rect 19478 17380 19484 17382
rect 19540 17380 19564 17382
rect 19620 17380 19644 17382
rect 19700 17380 19724 17382
rect 19780 17380 19786 17382
rect 19478 17360 19786 17380
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 15994 19288 16594
rect 19352 16590 19380 17138
rect 19720 16658 19748 17138
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19812 16590 19840 17206
rect 19904 17134 19932 17614
rect 19996 17270 20024 18244
rect 20088 17524 20116 20742
rect 20364 20466 20392 20742
rect 20168 20460 20220 20466
rect 20352 20460 20404 20466
rect 20220 20420 20300 20448
rect 20168 20402 20220 20408
rect 20168 20052 20220 20058
rect 20272 20040 20300 20420
rect 20352 20402 20404 20408
rect 20352 20052 20404 20058
rect 20272 20012 20352 20040
rect 20168 19994 20220 20000
rect 20352 19994 20404 20000
rect 20180 19446 20208 19994
rect 20168 19440 20220 19446
rect 20220 19400 20300 19428
rect 20168 19382 20220 19388
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 20180 18290 20208 18770
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20180 17678 20208 18226
rect 20272 18222 20300 19400
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 20088 17496 20208 17524
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 19892 17128 19944 17134
rect 19944 17088 20024 17116
rect 19892 17070 19944 17076
rect 19892 16652 19944 16658
rect 19892 16594 19944 16600
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19352 16114 19380 16526
rect 19478 16348 19786 16368
rect 19478 16346 19484 16348
rect 19540 16346 19564 16348
rect 19620 16346 19644 16348
rect 19700 16346 19724 16348
rect 19780 16346 19786 16348
rect 19540 16294 19542 16346
rect 19722 16294 19724 16346
rect 19478 16292 19484 16294
rect 19540 16292 19564 16294
rect 19620 16292 19644 16294
rect 19700 16292 19724 16294
rect 19780 16292 19786 16294
rect 19478 16272 19786 16292
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19260 15966 19380 15994
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 19352 14482 19380 15966
rect 19904 15586 19932 16594
rect 19996 16046 20024 17088
rect 20088 16250 20116 17138
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19904 15570 20116 15586
rect 19892 15564 20116 15570
rect 19944 15558 20116 15564
rect 19892 15506 19944 15512
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19892 15428 19944 15434
rect 19892 15370 19944 15376
rect 19478 15260 19786 15280
rect 19478 15258 19484 15260
rect 19540 15258 19564 15260
rect 19620 15258 19644 15260
rect 19700 15258 19724 15260
rect 19780 15258 19786 15260
rect 19540 15206 19542 15258
rect 19722 15206 19724 15258
rect 19478 15204 19484 15206
rect 19540 15204 19564 15206
rect 19620 15204 19644 15206
rect 19700 15204 19724 15206
rect 19780 15204 19786 15206
rect 19478 15184 19786 15204
rect 19904 15162 19932 15370
rect 19892 15156 19944 15162
rect 19892 15098 19944 15104
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19720 14822 19748 14894
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 18984 14368 19196 14396
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18984 11626 19012 12718
rect 19076 11762 19104 12786
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 18972 10464 19024 10470
rect 18892 10424 18972 10452
rect 18972 10406 19024 10412
rect 19076 10266 19104 10610
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18616 9110 18644 9522
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 18340 8022 18368 8230
rect 18328 8016 18380 8022
rect 18328 7958 18380 7964
rect 18432 7868 18460 8298
rect 18340 7840 18460 7868
rect 18340 7342 18368 7840
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18800 7410 18828 7686
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18340 6934 18368 7278
rect 18328 6928 18380 6934
rect 18328 6870 18380 6876
rect 18340 6390 18368 6870
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5778 18184 6054
rect 18340 5778 18368 6326
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 19076 4554 19104 8434
rect 19168 6866 19196 14368
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 14006 19288 14214
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19352 13326 19380 14282
rect 19478 14172 19786 14192
rect 19478 14170 19484 14172
rect 19540 14170 19564 14172
rect 19620 14170 19644 14172
rect 19700 14170 19724 14172
rect 19780 14170 19786 14172
rect 19540 14118 19542 14170
rect 19722 14118 19724 14170
rect 19478 14116 19484 14118
rect 19540 14116 19564 14118
rect 19620 14116 19644 14118
rect 19700 14116 19724 14118
rect 19780 14116 19786 14118
rect 19478 14096 19786 14116
rect 19904 13462 19932 15098
rect 19996 15094 20024 15438
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 19996 13394 20024 15030
rect 20088 14958 20116 15558
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19340 13320 19392 13326
rect 19812 13297 19840 13330
rect 19892 13320 19944 13326
rect 19340 13262 19392 13268
rect 19798 13288 19854 13297
rect 19892 13262 19944 13268
rect 19798 13223 19854 13232
rect 19478 13084 19786 13104
rect 19478 13082 19484 13084
rect 19540 13082 19564 13084
rect 19620 13082 19644 13084
rect 19700 13082 19724 13084
rect 19780 13082 19786 13084
rect 19540 13030 19542 13082
rect 19722 13030 19724 13082
rect 19478 13028 19484 13030
rect 19540 13028 19564 13030
rect 19620 13028 19644 13030
rect 19700 13028 19724 13030
rect 19780 13028 19786 13030
rect 19478 13008 19786 13028
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11898 19288 12038
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19260 11286 19288 11834
rect 19352 11506 19380 12786
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19444 12442 19472 12718
rect 19904 12442 19932 13262
rect 19996 12986 20024 13330
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 19892 12232 19944 12238
rect 19996 12220 20024 12922
rect 20088 12918 20116 13398
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19944 12192 20024 12220
rect 19892 12174 19944 12180
rect 19478 11996 19786 12016
rect 19478 11994 19484 11996
rect 19540 11994 19564 11996
rect 19620 11994 19644 11996
rect 19700 11994 19724 11996
rect 19780 11994 19786 11996
rect 19540 11942 19542 11994
rect 19722 11942 19724 11994
rect 19478 11940 19484 11942
rect 19540 11940 19564 11942
rect 19620 11940 19644 11942
rect 19700 11940 19724 11942
rect 19780 11940 19786 11942
rect 19478 11920 19786 11940
rect 19798 11792 19854 11801
rect 19798 11727 19800 11736
rect 19852 11727 19854 11736
rect 19800 11698 19852 11704
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19536 11506 19564 11562
rect 19352 11478 19564 11506
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19352 9586 19380 11478
rect 19478 10908 19786 10928
rect 19478 10906 19484 10908
rect 19540 10906 19564 10908
rect 19620 10906 19644 10908
rect 19700 10906 19724 10908
rect 19780 10906 19786 10908
rect 19540 10854 19542 10906
rect 19722 10854 19724 10906
rect 19478 10852 19484 10854
rect 19540 10852 19564 10854
rect 19620 10852 19644 10854
rect 19700 10852 19724 10854
rect 19780 10852 19786 10854
rect 19478 10832 19786 10852
rect 19904 10606 19932 12174
rect 20088 11286 20116 12582
rect 20180 12102 20208 17496
rect 20260 17264 20312 17270
rect 20260 17206 20312 17212
rect 20272 16658 20300 17206
rect 20364 16776 20392 19994
rect 20456 18766 20484 20810
rect 20548 20534 20576 22986
rect 20640 21418 20668 23276
rect 20824 22642 20852 23530
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20732 21418 20760 21898
rect 20824 21622 20852 22578
rect 20812 21616 20864 21622
rect 20812 21558 20864 21564
rect 20916 21536 20944 24024
rect 21284 23118 21312 24142
rect 21732 23656 21784 23662
rect 21732 23598 21784 23604
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21744 21894 21772 23598
rect 21836 23186 21864 24550
rect 22008 24200 22060 24206
rect 22008 24142 22060 24148
rect 22020 23798 22048 24142
rect 22008 23792 22060 23798
rect 22008 23734 22060 23740
rect 22112 23662 22140 25706
rect 22204 24818 22232 25910
rect 23400 25838 23428 26862
rect 24676 26852 24728 26858
rect 24676 26794 24728 26800
rect 24110 26684 24418 26704
rect 24110 26682 24116 26684
rect 24172 26682 24196 26684
rect 24252 26682 24276 26684
rect 24332 26682 24356 26684
rect 24412 26682 24418 26684
rect 24172 26630 24174 26682
rect 24354 26630 24356 26682
rect 24110 26628 24116 26630
rect 24172 26628 24196 26630
rect 24252 26628 24276 26630
rect 24332 26628 24356 26630
rect 24412 26628 24418 26630
rect 24110 26608 24418 26628
rect 23756 25900 23808 25906
rect 23756 25842 23808 25848
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 22376 25356 22428 25362
rect 22376 25298 22428 25304
rect 22388 24954 22416 25298
rect 23400 25294 23428 25774
rect 23768 25498 23796 25842
rect 24110 25596 24418 25616
rect 24110 25594 24116 25596
rect 24172 25594 24196 25596
rect 24252 25594 24276 25596
rect 24332 25594 24356 25596
rect 24412 25594 24418 25596
rect 24172 25542 24174 25594
rect 24354 25542 24356 25594
rect 24110 25540 24116 25542
rect 24172 25540 24196 25542
rect 24252 25540 24276 25542
rect 24332 25540 24356 25542
rect 24412 25540 24418 25542
rect 24110 25520 24418 25540
rect 23756 25492 23808 25498
rect 23756 25434 23808 25440
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 22376 24948 22428 24954
rect 22376 24890 22428 24896
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22388 24614 22416 24754
rect 22468 24676 22520 24682
rect 22468 24618 22520 24624
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 22204 23730 22232 24142
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21928 23050 21956 23462
rect 22112 23118 22140 23598
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22388 23066 22416 24006
rect 22480 23322 22508 24618
rect 22664 24206 22692 25230
rect 23020 24880 23072 24886
rect 23020 24822 23072 24828
rect 23032 24682 23060 24822
rect 23020 24676 23072 24682
rect 23020 24618 23072 24624
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22664 23322 22692 24142
rect 23296 24132 23348 24138
rect 23296 24074 23348 24080
rect 23308 23866 23336 24074
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23860 23730 23888 24550
rect 24110 24508 24418 24528
rect 24110 24506 24116 24508
rect 24172 24506 24196 24508
rect 24252 24506 24276 24508
rect 24332 24506 24356 24508
rect 24412 24506 24418 24508
rect 24172 24454 24174 24506
rect 24354 24454 24356 24506
rect 24110 24452 24116 24454
rect 24172 24452 24196 24454
rect 24252 24452 24276 24454
rect 24332 24452 24356 24454
rect 24412 24452 24418 24454
rect 24110 24432 24418 24452
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24504 23798 24532 24006
rect 24492 23792 24544 23798
rect 24492 23734 24544 23740
rect 23848 23724 23900 23730
rect 23848 23666 23900 23672
rect 23756 23656 23808 23662
rect 23492 23616 23756 23644
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22468 23112 22520 23118
rect 22388 23060 22468 23066
rect 22388 23054 22520 23060
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 22388 23038 22508 23054
rect 21824 22636 21876 22642
rect 21928 22624 21956 22986
rect 21876 22596 21956 22624
rect 21824 22578 21876 22584
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 20916 21508 21036 21536
rect 20628 21412 20680 21418
rect 20628 21354 20680 21360
rect 20720 21412 20772 21418
rect 20720 21354 20772 21360
rect 21008 21078 21036 21508
rect 21192 21350 21220 21626
rect 21928 21554 21956 22596
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 20996 21072 21048 21078
rect 20996 21014 21048 21020
rect 21824 21072 21876 21078
rect 21824 21014 21876 21020
rect 21008 20942 21036 21014
rect 21364 21004 21416 21010
rect 21364 20946 21416 20952
rect 20628 20936 20680 20942
rect 20628 20878 20680 20884
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 20640 20602 20668 20878
rect 20628 20596 20680 20602
rect 20680 20556 20760 20584
rect 20628 20538 20680 20544
rect 20536 20528 20588 20534
rect 20536 20470 20588 20476
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 19258 20668 19654
rect 20732 19378 20760 20556
rect 20824 19514 20852 20878
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 21100 20058 21128 20334
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20720 19372 20772 19378
rect 21376 19360 21404 20946
rect 21836 20942 21864 21014
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21928 20330 21956 21490
rect 22112 21146 22140 21490
rect 22192 21344 22244 21350
rect 22192 21286 22244 21292
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 22204 20942 22232 21286
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 21916 20324 21968 20330
rect 21916 20266 21968 20272
rect 22388 19854 22416 23038
rect 22664 22710 22692 23258
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 22928 23044 22980 23050
rect 22928 22986 22980 22992
rect 22652 22704 22704 22710
rect 22652 22646 22704 22652
rect 22940 22574 22968 22986
rect 23400 22642 23428 23190
rect 23492 23186 23520 23616
rect 23756 23598 23808 23604
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 23480 23180 23532 23186
rect 23480 23122 23532 23128
rect 23952 23118 23980 23598
rect 24110 23420 24418 23440
rect 24110 23418 24116 23420
rect 24172 23418 24196 23420
rect 24252 23418 24276 23420
rect 24332 23418 24356 23420
rect 24412 23418 24418 23420
rect 24172 23366 24174 23418
rect 24354 23366 24356 23418
rect 24110 23364 24116 23366
rect 24172 23364 24196 23366
rect 24252 23364 24276 23366
rect 24332 23364 24356 23366
rect 24412 23364 24418 23366
rect 24110 23344 24418 23364
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23940 23112 23992 23118
rect 23940 23054 23992 23060
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 22928 22568 22980 22574
rect 22928 22510 22980 22516
rect 23492 22234 23520 22918
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 23480 22228 23532 22234
rect 23480 22170 23532 22176
rect 23584 22030 23612 22442
rect 23676 22094 23704 22918
rect 23768 22778 23796 23054
rect 24492 23044 24544 23050
rect 24492 22986 24544 22992
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 23952 22522 23980 22646
rect 24216 22636 24268 22642
rect 23860 22506 23980 22522
rect 23848 22500 23980 22506
rect 23900 22494 23980 22500
rect 24044 22596 24216 22624
rect 23848 22442 23900 22448
rect 23676 22066 23796 22094
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23492 21690 23520 21830
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 22926 21448 22982 21457
rect 22926 21383 22982 21392
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 21468 19689 21496 19790
rect 21454 19680 21510 19689
rect 21454 19615 21510 19624
rect 21456 19372 21508 19378
rect 21376 19332 21456 19360
rect 20720 19314 20772 19320
rect 21456 19314 21508 19320
rect 20640 19230 20760 19258
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 20536 18964 20588 18970
rect 20640 18952 20668 19110
rect 20588 18924 20668 18952
rect 20536 18906 20588 18912
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20456 18290 20484 18702
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20640 17218 20668 18924
rect 20732 18766 20760 19230
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20732 18086 20760 18702
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 21192 18086 21220 18158
rect 21376 18154 21404 18566
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 20720 18080 20772 18086
rect 21180 18080 21232 18086
rect 20772 18040 20852 18068
rect 20720 18022 20772 18028
rect 20824 17678 20852 18040
rect 21180 18022 21232 18028
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20732 17338 20760 17614
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20640 17202 20760 17218
rect 20640 17196 20772 17202
rect 20640 17190 20720 17196
rect 20720 17138 20772 17144
rect 20732 16998 20760 17138
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20444 16788 20496 16794
rect 20364 16748 20444 16776
rect 20444 16730 20496 16736
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20260 15428 20312 15434
rect 20260 15370 20312 15376
rect 20272 14890 20300 15370
rect 20456 15026 20484 15846
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20260 14884 20312 14890
rect 20260 14826 20312 14832
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20272 14074 20300 14350
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20272 12646 20300 13466
rect 20364 13190 20392 14962
rect 20548 14890 20576 15302
rect 20732 15178 20760 16390
rect 20916 16114 20944 16662
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20824 15434 20852 16050
rect 21008 15502 21036 17478
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 21100 16182 21128 16934
rect 21192 16522 21220 18022
rect 21376 17134 21404 18090
rect 21560 17542 21588 19790
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22192 19712 22244 19718
rect 22296 19689 22324 19722
rect 22192 19654 22244 19660
rect 22282 19680 22338 19689
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 21548 17536 21600 17542
rect 21548 17478 21600 17484
rect 21652 17354 21680 18362
rect 21560 17326 21680 17354
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21468 16250 21496 16390
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21088 16176 21140 16182
rect 21088 16118 21140 16124
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20640 15150 20760 15178
rect 20640 15094 20668 15150
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20536 14884 20588 14890
rect 20536 14826 20588 14832
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20456 13938 20484 14350
rect 20824 13938 20852 15370
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20916 14278 20944 14758
rect 20996 14408 21048 14414
rect 20994 14376 20996 14385
rect 21048 14376 21050 14385
rect 20994 14311 21050 14320
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 14113 20944 14214
rect 20902 14104 20958 14113
rect 20902 14039 20958 14048
rect 21100 14006 21128 16118
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21284 15570 21312 16050
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21376 15094 21404 15302
rect 21364 15088 21416 15094
rect 21364 15030 21416 15036
rect 21362 14104 21418 14113
rect 21362 14039 21418 14048
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20364 12918 20392 13126
rect 20456 12986 20484 13194
rect 20548 13025 20576 13874
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20534 13016 20590 13025
rect 20444 12980 20496 12986
rect 20534 12951 20590 12960
rect 20444 12922 20496 12928
rect 20352 12912 20404 12918
rect 20352 12854 20404 12860
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19892 10600 19944 10606
rect 19892 10542 19944 10548
rect 19444 10198 19472 10542
rect 19996 10266 20024 11086
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19982 10160 20038 10169
rect 19982 10095 20038 10104
rect 19996 10062 20024 10095
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19478 9820 19786 9840
rect 19478 9818 19484 9820
rect 19540 9818 19564 9820
rect 19620 9818 19644 9820
rect 19700 9818 19724 9820
rect 19780 9818 19786 9820
rect 19540 9766 19542 9818
rect 19722 9766 19724 9818
rect 19478 9764 19484 9766
rect 19540 9764 19564 9766
rect 19620 9764 19644 9766
rect 19700 9764 19724 9766
rect 19780 9764 19786 9766
rect 19478 9744 19786 9764
rect 19904 9586 19932 9862
rect 20088 9654 20116 11222
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20180 10130 20208 11154
rect 20272 11014 20300 12378
rect 20548 11694 20576 12951
rect 20640 12850 20668 13670
rect 21100 13530 21128 13806
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12850 21128 13126
rect 21376 12986 21404 14039
rect 21560 13938 21588 17326
rect 21836 16726 21864 19314
rect 22204 19281 22232 19654
rect 22282 19615 22338 19624
rect 22296 19378 22324 19615
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22190 19272 22246 19281
rect 22190 19207 22246 19216
rect 22296 18970 22324 19314
rect 22572 18970 22600 20878
rect 22652 19236 22704 19242
rect 22652 19178 22704 19184
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22468 18896 22520 18902
rect 22468 18838 22520 18844
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22112 18290 22140 18770
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22008 18216 22060 18222
rect 22008 18158 22060 18164
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21928 17746 21956 17818
rect 21916 17740 21968 17746
rect 21916 17682 21968 17688
rect 21928 17202 21956 17682
rect 22020 17678 22048 18158
rect 22112 17678 22140 18226
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 21916 17196 21968 17202
rect 21916 17138 21968 17144
rect 22388 17066 22416 18566
rect 22480 17270 22508 18838
rect 22664 18834 22692 19178
rect 22652 18828 22704 18834
rect 22652 18770 22704 18776
rect 22940 18426 22968 21383
rect 23584 21350 23612 21966
rect 23676 21418 23704 21966
rect 23664 21412 23716 21418
rect 23664 21354 23716 21360
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 23124 20466 23152 20946
rect 23676 20942 23704 21354
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23204 20868 23256 20874
rect 23204 20810 23256 20816
rect 23296 20868 23348 20874
rect 23296 20810 23348 20816
rect 23112 20460 23164 20466
rect 23112 20402 23164 20408
rect 23216 20398 23244 20810
rect 23204 20392 23256 20398
rect 23204 20334 23256 20340
rect 23308 20058 23336 20810
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23492 19854 23520 20402
rect 23676 19990 23704 20538
rect 23664 19984 23716 19990
rect 23664 19926 23716 19932
rect 23676 19854 23704 19926
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23294 18456 23350 18465
rect 22928 18420 22980 18426
rect 23294 18391 23350 18400
rect 22928 18362 22980 18368
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 22940 18154 22968 18226
rect 23308 18154 23336 18391
rect 22928 18148 22980 18154
rect 22928 18090 22980 18096
rect 23296 18148 23348 18154
rect 23296 18090 23348 18096
rect 22468 17264 22520 17270
rect 22468 17206 22520 17212
rect 21916 17060 21968 17066
rect 21916 17002 21968 17008
rect 22376 17060 22428 17066
rect 22376 17002 22428 17008
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21652 15706 21680 16526
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 21744 15162 21772 15506
rect 21928 15484 21956 17002
rect 22008 16720 22060 16726
rect 22008 16662 22060 16668
rect 22020 16182 22048 16662
rect 22008 16176 22060 16182
rect 22008 16118 22060 16124
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 22296 15502 22324 15846
rect 22284 15496 22336 15502
rect 21928 15456 22048 15484
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21652 14074 21680 14214
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21468 13433 21496 13670
rect 21652 13530 21680 13874
rect 21744 13734 21772 14962
rect 21916 14544 21968 14550
rect 21916 14486 21968 14492
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21928 13530 21956 14486
rect 22020 14414 22048 15456
rect 22284 15438 22336 15444
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22112 14414 22140 15030
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22112 14278 22140 14350
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21454 13424 21510 13433
rect 21454 13359 21510 13368
rect 21836 13190 21864 13466
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21836 12850 21864 13126
rect 21928 12968 21956 13466
rect 21928 12940 22048 12968
rect 22020 12850 22048 12940
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 20626 12744 20682 12753
rect 20626 12679 20628 12688
rect 20680 12679 20682 12688
rect 20628 12650 20680 12656
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20640 11898 20668 12174
rect 20732 12170 20760 12582
rect 22112 12481 22140 14214
rect 22296 13938 22324 15438
rect 22560 15428 22612 15434
rect 22560 15370 22612 15376
rect 22572 15162 22600 15370
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22560 14952 22612 14958
rect 22560 14894 22612 14900
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22296 13530 22324 13670
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22388 13190 22416 13670
rect 22480 13190 22508 14350
rect 22572 14278 22600 14894
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22572 14074 22600 14214
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22480 13002 22508 13126
rect 22558 13016 22614 13025
rect 22480 12974 22558 13002
rect 22558 12951 22560 12960
rect 22612 12951 22614 12960
rect 22560 12922 22612 12928
rect 22098 12472 22154 12481
rect 22098 12407 22154 12416
rect 22112 12238 22140 12407
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22468 12232 22520 12238
rect 22572 12220 22600 12922
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22520 12192 22600 12220
rect 22468 12174 22520 12180
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 21008 11762 21036 12038
rect 21744 11762 21772 12174
rect 22008 12164 22060 12170
rect 22008 12106 22060 12112
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 22020 11626 22048 12106
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22572 11762 22600 12038
rect 22376 11756 22428 11762
rect 22560 11756 22612 11762
rect 22428 11716 22508 11744
rect 22376 11698 22428 11704
rect 22282 11656 22338 11665
rect 22008 11620 22060 11626
rect 22282 11591 22338 11600
rect 22008 11562 22060 11568
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20824 11082 20852 11494
rect 22020 11354 22048 11562
rect 22296 11354 22324 11591
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20640 10266 20668 10610
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 20180 9518 20208 10066
rect 20732 10062 20760 11018
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 21284 10198 21312 10406
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 21192 9586 21220 9862
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 19720 9042 19748 9454
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19352 8498 19380 8978
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19478 8732 19786 8752
rect 19478 8730 19484 8732
rect 19540 8730 19564 8732
rect 19620 8730 19644 8732
rect 19700 8730 19724 8732
rect 19780 8730 19786 8732
rect 19540 8678 19542 8730
rect 19722 8678 19724 8730
rect 19478 8676 19484 8678
rect 19540 8676 19564 8678
rect 19620 8676 19644 8678
rect 19700 8676 19724 8678
rect 19780 8676 19786 8678
rect 19478 8656 19786 8676
rect 19996 8566 20024 8774
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19352 7886 19380 8230
rect 19812 8090 19840 8434
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 20364 7954 20392 8910
rect 20824 8906 20852 9046
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21008 8498 21036 8774
rect 21100 8634 21128 8774
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 19478 7644 19786 7664
rect 19478 7642 19484 7644
rect 19540 7642 19564 7644
rect 19620 7642 19644 7644
rect 19700 7642 19724 7644
rect 19780 7642 19786 7644
rect 19540 7590 19542 7642
rect 19722 7590 19724 7642
rect 19478 7588 19484 7590
rect 19540 7588 19564 7590
rect 19620 7588 19644 7590
rect 19700 7588 19724 7590
rect 19780 7588 19786 7590
rect 19478 7568 19786 7588
rect 19904 7206 19932 7754
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19260 5234 19288 6598
rect 19352 5914 19380 6734
rect 19478 6556 19786 6576
rect 19478 6554 19484 6556
rect 19540 6554 19564 6556
rect 19620 6554 19644 6556
rect 19700 6554 19724 6556
rect 19780 6554 19786 6556
rect 19540 6502 19542 6554
rect 19722 6502 19724 6554
rect 19478 6500 19484 6502
rect 19540 6500 19564 6502
rect 19620 6500 19644 6502
rect 19700 6500 19724 6502
rect 19780 6500 19786 6502
rect 19478 6480 19786 6500
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19720 5710 19748 6054
rect 19812 5846 19840 6258
rect 19800 5840 19852 5846
rect 19800 5782 19852 5788
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 19904 5642 19932 7142
rect 19996 6866 20024 7890
rect 20364 7478 20392 7890
rect 20456 7886 20484 8230
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 19996 6254 20024 6802
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 20364 5778 20392 7414
rect 21284 6798 21312 10134
rect 22112 9586 22140 10406
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21376 8022 21404 8910
rect 22112 8906 22140 9522
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 21836 8634 21864 8842
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21364 8016 21416 8022
rect 21364 7958 21416 7964
rect 21376 7478 21404 7958
rect 22112 7954 22140 8842
rect 22204 8498 22232 9862
rect 22296 9586 22324 11018
rect 22388 10742 22416 11494
rect 22480 11218 22508 11716
rect 22560 11698 22612 11704
rect 22664 11626 22692 12718
rect 22756 12646 22784 13262
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22940 12434 22968 18090
rect 23676 17746 23704 19314
rect 23768 19258 23796 22066
rect 23848 22024 23900 22030
rect 24044 21978 24072 22596
rect 24216 22578 24268 22584
rect 24110 22332 24418 22352
rect 24110 22330 24116 22332
rect 24172 22330 24196 22332
rect 24252 22330 24276 22332
rect 24332 22330 24356 22332
rect 24412 22330 24418 22332
rect 24172 22278 24174 22330
rect 24354 22278 24356 22330
rect 24110 22276 24116 22278
rect 24172 22276 24196 22278
rect 24252 22276 24276 22278
rect 24332 22276 24356 22278
rect 24412 22276 24418 22278
rect 24110 22256 24418 22276
rect 24306 22128 24362 22137
rect 24306 22063 24308 22072
rect 24360 22063 24362 22072
rect 24308 22034 24360 22040
rect 23900 21972 24072 21978
rect 23848 21966 24072 21972
rect 23860 21950 24072 21966
rect 24306 21992 24362 22001
rect 24306 21927 24308 21936
rect 24360 21927 24362 21936
rect 24308 21898 24360 21904
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23848 21412 23900 21418
rect 23848 21354 23900 21360
rect 23860 21146 23888 21354
rect 23952 21350 23980 21490
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 24110 21244 24418 21264
rect 24110 21242 24116 21244
rect 24172 21242 24196 21244
rect 24252 21242 24276 21244
rect 24332 21242 24356 21244
rect 24412 21242 24418 21244
rect 24172 21190 24174 21242
rect 24354 21190 24356 21242
rect 24110 21188 24116 21190
rect 24172 21188 24196 21190
rect 24252 21188 24276 21190
rect 24332 21188 24356 21190
rect 24412 21188 24418 21190
rect 24110 21168 24418 21188
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 24400 21072 24452 21078
rect 24504 21060 24532 22986
rect 24596 22778 24624 23598
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24584 22500 24636 22506
rect 24584 22442 24636 22448
rect 24596 22166 24624 22442
rect 24584 22160 24636 22166
rect 24584 22102 24636 22108
rect 24688 21894 24716 26794
rect 25516 26353 25544 26930
rect 25134 26344 25190 26353
rect 25134 26279 25136 26288
rect 25188 26279 25190 26288
rect 25502 26344 25558 26353
rect 25502 26279 25558 26288
rect 25136 26250 25188 26256
rect 25688 25968 25740 25974
rect 25688 25910 25740 25916
rect 25412 25900 25464 25906
rect 25412 25842 25464 25848
rect 25596 25900 25648 25906
rect 25596 25842 25648 25848
rect 24768 25696 24820 25702
rect 24768 25638 24820 25644
rect 24780 25362 24808 25638
rect 24768 25356 24820 25362
rect 24768 25298 24820 25304
rect 24780 24818 24808 25298
rect 24860 25288 24912 25294
rect 24912 25248 24992 25276
rect 24860 25230 24912 25236
rect 24768 24812 24820 24818
rect 24768 24754 24820 24760
rect 24780 24138 24808 24754
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24768 24132 24820 24138
rect 24768 24074 24820 24080
rect 24780 23798 24808 24074
rect 24872 23798 24900 24142
rect 24768 23792 24820 23798
rect 24768 23734 24820 23740
rect 24860 23792 24912 23798
rect 24860 23734 24912 23740
rect 24964 22982 24992 25248
rect 25424 25226 25452 25842
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 25608 24954 25636 25842
rect 25700 25498 25728 25910
rect 25780 25900 25832 25906
rect 25780 25842 25832 25848
rect 25688 25492 25740 25498
rect 25688 25434 25740 25440
rect 25596 24948 25648 24954
rect 25596 24890 25648 24896
rect 25700 24818 25728 25434
rect 25792 25362 25820 25842
rect 25780 25356 25832 25362
rect 25780 25298 25832 25304
rect 25780 25220 25832 25226
rect 25780 25162 25832 25168
rect 25688 24812 25740 24818
rect 25688 24754 25740 24760
rect 25136 24676 25188 24682
rect 25136 24618 25188 24624
rect 25148 24138 25176 24618
rect 25700 24410 25728 24754
rect 25792 24410 25820 25162
rect 25688 24404 25740 24410
rect 25688 24346 25740 24352
rect 25780 24404 25832 24410
rect 25780 24346 25832 24352
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25412 24268 25464 24274
rect 25412 24210 25464 24216
rect 25136 24132 25188 24138
rect 25136 24074 25188 24080
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 25056 23254 25084 23666
rect 25148 23594 25176 24074
rect 25240 23866 25268 24210
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25228 23656 25280 23662
rect 25228 23598 25280 23604
rect 25136 23588 25188 23594
rect 25136 23530 25188 23536
rect 25240 23322 25268 23598
rect 25424 23338 25452 24210
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 25504 23724 25556 23730
rect 25504 23666 25556 23672
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 25332 23310 25452 23338
rect 25516 23322 25544 23666
rect 25504 23316 25556 23322
rect 25044 23248 25096 23254
rect 25044 23190 25096 23196
rect 24952 22976 25004 22982
rect 24952 22918 25004 22924
rect 25044 22772 25096 22778
rect 25044 22714 25096 22720
rect 24768 22500 24820 22506
rect 24768 22442 24820 22448
rect 24780 22234 24808 22442
rect 24768 22228 24820 22234
rect 24768 22170 24820 22176
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24780 21690 24808 22170
rect 24952 22092 25004 22098
rect 24952 22034 25004 22040
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24780 21554 24808 21626
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24872 21434 24900 21966
rect 24964 21457 24992 22034
rect 25056 22001 25084 22714
rect 25240 22574 25268 23258
rect 25332 22710 25360 23310
rect 25504 23258 25556 23264
rect 25792 23186 25820 24006
rect 25780 23180 25832 23186
rect 25780 23122 25832 23128
rect 25504 23112 25556 23118
rect 25884 23066 25912 27338
rect 27344 27328 27396 27334
rect 27344 27270 27396 27276
rect 26148 27056 26200 27062
rect 26148 26998 26200 27004
rect 25964 25696 26016 25702
rect 25964 25638 26016 25644
rect 25976 25226 26004 25638
rect 26160 25294 26188 26998
rect 26700 26920 26752 26926
rect 26700 26862 26752 26868
rect 26712 26314 26740 26862
rect 26700 26308 26752 26314
rect 26700 26250 26752 26256
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 25964 25220 26016 25226
rect 25964 25162 26016 25168
rect 25964 23860 26016 23866
rect 25964 23802 26016 23808
rect 25976 23118 26004 23802
rect 26148 23792 26200 23798
rect 26148 23734 26200 23740
rect 26160 23118 26188 23734
rect 25504 23054 25556 23060
rect 25320 22704 25372 22710
rect 25320 22646 25372 22652
rect 25228 22568 25280 22574
rect 25228 22510 25280 22516
rect 25042 21992 25098 22001
rect 25098 21950 25176 21978
rect 25042 21927 25098 21936
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 24452 21032 24532 21060
rect 24400 21014 24452 21020
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23860 20466 23888 20878
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23860 20058 23888 20402
rect 24032 20256 24084 20262
rect 24032 20198 24084 20204
rect 23848 20052 23900 20058
rect 23848 19994 23900 20000
rect 24044 19854 24072 20198
rect 24110 20156 24418 20176
rect 24110 20154 24116 20156
rect 24172 20154 24196 20156
rect 24252 20154 24276 20156
rect 24332 20154 24356 20156
rect 24412 20154 24418 20156
rect 24172 20102 24174 20154
rect 24354 20102 24356 20154
rect 24110 20100 24116 20102
rect 24172 20100 24196 20102
rect 24252 20100 24276 20102
rect 24332 20100 24356 20102
rect 24412 20100 24418 20102
rect 24110 20080 24418 20100
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 23940 19712 23992 19718
rect 23940 19654 23992 19660
rect 23952 19514 23980 19654
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 23938 19408 23994 19417
rect 23938 19343 23940 19352
rect 23992 19343 23994 19352
rect 23940 19314 23992 19320
rect 23768 19230 23888 19258
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 23768 18766 23796 19110
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23860 17882 23888 19230
rect 23952 18465 23980 19314
rect 24044 18970 24072 19790
rect 24504 19446 24532 21032
rect 24596 21406 24900 21434
rect 24950 21448 25006 21457
rect 24596 20330 24624 21406
rect 24950 21383 25006 21392
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24688 21146 24716 21286
rect 24676 21140 24728 21146
rect 24676 21082 24728 21088
rect 24688 21010 24716 21082
rect 24860 21072 24912 21078
rect 25056 21060 25084 21490
rect 24912 21032 25084 21060
rect 24860 21014 24912 21020
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24584 20324 24636 20330
rect 24584 20266 24636 20272
rect 24492 19440 24544 19446
rect 24492 19382 24544 19388
rect 24596 19334 24624 20266
rect 24688 19854 24716 20946
rect 24768 20936 24820 20942
rect 24952 20936 25004 20942
rect 24768 20878 24820 20884
rect 24872 20884 24952 20890
rect 24872 20878 25004 20884
rect 24780 20398 24808 20878
rect 24872 20862 24992 20878
rect 24768 20392 24820 20398
rect 24768 20334 24820 20340
rect 24780 19922 24808 20334
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24872 19854 24900 20862
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24492 19304 24544 19310
rect 24596 19306 24716 19334
rect 24492 19246 24544 19252
rect 24110 19068 24418 19088
rect 24110 19066 24116 19068
rect 24172 19066 24196 19068
rect 24252 19066 24276 19068
rect 24332 19066 24356 19068
rect 24412 19066 24418 19068
rect 24172 19014 24174 19066
rect 24354 19014 24356 19066
rect 24110 19012 24116 19014
rect 24172 19012 24196 19014
rect 24252 19012 24276 19014
rect 24332 19012 24356 19014
rect 24412 19012 24418 19014
rect 24110 18992 24418 19012
rect 24504 18970 24532 19246
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24032 18964 24084 18970
rect 24032 18906 24084 18912
rect 24492 18964 24544 18970
rect 24492 18906 24544 18912
rect 23938 18456 23994 18465
rect 23938 18391 23994 18400
rect 24044 18290 24072 18906
rect 24596 18426 24624 19110
rect 24688 18902 24716 19306
rect 24872 19009 24900 19790
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 24858 19000 24914 19009
rect 24858 18935 24914 18944
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 25056 18766 25084 19450
rect 25148 19446 25176 21950
rect 25332 21026 25360 22646
rect 25516 22438 25544 23054
rect 25792 23038 25912 23066
rect 25964 23112 26016 23118
rect 25964 23054 26016 23060
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 25412 22432 25464 22438
rect 25412 22374 25464 22380
rect 25504 22432 25556 22438
rect 25504 22374 25556 22380
rect 25424 21622 25452 22374
rect 25502 22128 25558 22137
rect 25608 22114 25636 22578
rect 25558 22086 25636 22114
rect 25502 22063 25558 22072
rect 25516 21962 25544 22063
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25516 21622 25544 21898
rect 25412 21616 25464 21622
rect 25412 21558 25464 21564
rect 25504 21616 25556 21622
rect 25504 21558 25556 21564
rect 25240 20998 25360 21026
rect 25240 20806 25268 20998
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25228 20800 25280 20806
rect 25228 20742 25280 20748
rect 25332 20466 25360 20878
rect 25320 20460 25372 20466
rect 25320 20402 25372 20408
rect 25424 19854 25452 21558
rect 25688 21004 25740 21010
rect 25688 20946 25740 20952
rect 25700 20534 25728 20946
rect 25504 20528 25556 20534
rect 25504 20470 25556 20476
rect 25688 20528 25740 20534
rect 25792 20505 25820 23038
rect 26056 22500 26108 22506
rect 26056 22442 26108 22448
rect 25872 22432 25924 22438
rect 25872 22374 25924 22380
rect 25884 21350 25912 22374
rect 26068 22098 26096 22442
rect 26056 22092 26108 22098
rect 26056 22034 26108 22040
rect 25964 22024 26016 22030
rect 25964 21966 26016 21972
rect 25976 21894 26004 21966
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 26516 21888 26568 21894
rect 26516 21830 26568 21836
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25872 20936 25924 20942
rect 25872 20878 25924 20884
rect 25884 20602 25912 20878
rect 25872 20596 25924 20602
rect 25872 20538 25924 20544
rect 25688 20470 25740 20476
rect 25778 20496 25834 20505
rect 25516 20398 25544 20470
rect 25596 20460 25648 20466
rect 25778 20431 25834 20440
rect 25596 20402 25648 20408
rect 25504 20392 25556 20398
rect 25504 20334 25556 20340
rect 25608 19990 25636 20402
rect 25596 19984 25648 19990
rect 25596 19926 25648 19932
rect 25412 19848 25464 19854
rect 25332 19796 25412 19802
rect 25332 19790 25464 19796
rect 25332 19774 25452 19790
rect 25136 19440 25188 19446
rect 25136 19382 25188 19388
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 25148 18698 25176 19382
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24110 17980 24418 18000
rect 24110 17978 24116 17980
rect 24172 17978 24196 17980
rect 24252 17978 24276 17980
rect 24332 17978 24356 17980
rect 24412 17978 24418 17980
rect 24172 17926 24174 17978
rect 24354 17926 24356 17978
rect 24110 17924 24116 17926
rect 24172 17924 24196 17926
rect 24252 17924 24276 17926
rect 24332 17924 24356 17926
rect 24412 17924 24418 17926
rect 24110 17904 24418 17924
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 24492 17740 24544 17746
rect 24492 17682 24544 17688
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23124 17202 23152 17614
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 23216 14346 23244 17478
rect 24504 17134 24532 17682
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24584 17196 24636 17202
rect 24872 17184 24900 17614
rect 25136 17604 25188 17610
rect 25332 17592 25360 19774
rect 25884 19718 25912 20538
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25504 19712 25556 19718
rect 25504 19654 25556 19660
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 25424 18426 25452 19654
rect 25516 19514 25544 19654
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25976 19394 26004 21830
rect 26148 21548 26200 21554
rect 26148 21490 26200 21496
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 26068 20942 26096 21286
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 26068 20398 26096 20878
rect 26056 20392 26108 20398
rect 26056 20334 26108 20340
rect 25884 19366 26004 19394
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 25516 17882 25544 18770
rect 25884 18766 25912 19366
rect 25964 19304 26016 19310
rect 25964 19246 26016 19252
rect 25976 18970 26004 19246
rect 25964 18964 26016 18970
rect 25964 18906 26016 18912
rect 25872 18760 25924 18766
rect 25872 18702 25924 18708
rect 25884 18290 25912 18702
rect 26068 18290 26096 20334
rect 25872 18284 25924 18290
rect 25872 18226 25924 18232
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 25504 17876 25556 17882
rect 25504 17818 25556 17824
rect 25516 17610 25544 17818
rect 25188 17564 25360 17592
rect 25504 17604 25556 17610
rect 25136 17546 25188 17552
rect 25504 17546 25556 17552
rect 25688 17604 25740 17610
rect 25688 17546 25740 17552
rect 24952 17196 25004 17202
rect 24636 17156 24952 17184
rect 24584 17138 24636 17144
rect 24952 17138 25004 17144
rect 25148 17134 25176 17546
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 23388 16992 23440 16998
rect 24952 16992 25004 16998
rect 23440 16940 23796 16946
rect 23388 16934 23796 16940
rect 24952 16934 25004 16940
rect 23400 16918 23796 16934
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23492 16114 23520 16390
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23584 15706 23612 16050
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23294 14512 23350 14521
rect 23294 14447 23350 14456
rect 23308 14414 23336 14447
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 23020 14340 23072 14346
rect 23020 14282 23072 14288
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 23032 13870 23060 14282
rect 23294 14104 23350 14113
rect 23294 14039 23296 14048
rect 23348 14039 23350 14048
rect 23296 14010 23348 14016
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 23216 13326 23244 13874
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23216 12918 23244 13262
rect 23308 13190 23336 13738
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23204 12912 23256 12918
rect 23204 12854 23256 12860
rect 23112 12640 23164 12646
rect 23112 12582 23164 12588
rect 22940 12406 23060 12434
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 22744 12164 22796 12170
rect 22744 12106 22796 12112
rect 22652 11620 22704 11626
rect 22652 11562 22704 11568
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22652 11144 22704 11150
rect 22756 11132 22784 12106
rect 22940 12102 22968 12174
rect 22928 12096 22980 12102
rect 22928 12038 22980 12044
rect 23032 11762 23060 12406
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 22848 11354 22876 11698
rect 23032 11665 23060 11698
rect 23018 11656 23074 11665
rect 23018 11591 23074 11600
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 23124 11150 23152 12582
rect 23216 12442 23244 12854
rect 23400 12832 23428 14758
rect 23676 14550 23704 14962
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23768 14249 23796 16918
rect 24110 16892 24418 16912
rect 24110 16890 24116 16892
rect 24172 16890 24196 16892
rect 24252 16890 24276 16892
rect 24332 16890 24356 16892
rect 24412 16890 24418 16892
rect 24172 16838 24174 16890
rect 24354 16838 24356 16890
rect 24110 16836 24116 16838
rect 24172 16836 24196 16838
rect 24252 16836 24276 16838
rect 24332 16836 24356 16838
rect 24412 16836 24418 16838
rect 24110 16816 24418 16836
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23860 16114 23888 16730
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23860 14278 23888 16050
rect 24110 15804 24418 15824
rect 24110 15802 24116 15804
rect 24172 15802 24196 15804
rect 24252 15802 24276 15804
rect 24332 15802 24356 15804
rect 24412 15802 24418 15804
rect 24172 15750 24174 15802
rect 24354 15750 24356 15802
rect 24110 15748 24116 15750
rect 24172 15748 24196 15750
rect 24252 15748 24276 15750
rect 24332 15748 24356 15750
rect 24412 15748 24418 15750
rect 24110 15728 24418 15748
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24872 15434 24900 15642
rect 24964 15502 24992 16934
rect 25136 16720 25188 16726
rect 25136 16662 25188 16668
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25056 15706 25084 16526
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 24044 14618 24072 14758
rect 24110 14716 24418 14736
rect 24110 14714 24116 14716
rect 24172 14714 24196 14716
rect 24252 14714 24276 14716
rect 24332 14714 24356 14716
rect 24412 14714 24418 14716
rect 24172 14662 24174 14714
rect 24354 14662 24356 14714
rect 24110 14660 24116 14662
rect 24172 14660 24196 14662
rect 24252 14660 24276 14662
rect 24332 14660 24356 14662
rect 24412 14660 24418 14662
rect 24110 14640 24418 14660
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 23848 14272 23900 14278
rect 23754 14240 23810 14249
rect 24044 14260 24072 14554
rect 24766 14512 24822 14521
rect 24584 14476 24636 14482
rect 24766 14447 24822 14456
rect 24584 14418 24636 14424
rect 24216 14272 24268 14278
rect 24044 14232 24164 14260
rect 23848 14214 23900 14220
rect 23754 14175 23810 14184
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 23584 13462 23612 13806
rect 23676 13530 23704 14010
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23572 13456 23624 13462
rect 23572 13398 23624 13404
rect 23768 12918 23796 14175
rect 24136 14074 24164 14232
rect 24216 14214 24268 14220
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 24044 13530 24072 13942
rect 24228 13938 24256 14214
rect 24596 14006 24624 14418
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24596 13870 24624 13942
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24492 13728 24544 13734
rect 24492 13670 24544 13676
rect 24110 13628 24418 13648
rect 24110 13626 24116 13628
rect 24172 13626 24196 13628
rect 24252 13626 24276 13628
rect 24332 13626 24356 13628
rect 24412 13626 24418 13628
rect 24172 13574 24174 13626
rect 24354 13574 24356 13626
rect 24110 13572 24116 13574
rect 24172 13572 24196 13574
rect 24252 13572 24276 13574
rect 24332 13572 24356 13574
rect 24412 13572 24418 13574
rect 24110 13552 24418 13572
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 24398 13424 24454 13433
rect 24398 13359 24454 13368
rect 24412 13326 24440 13359
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24504 12918 24532 13670
rect 24688 13530 24716 13874
rect 24676 13524 24728 13530
rect 24676 13466 24728 13472
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 24492 12912 24544 12918
rect 24492 12854 24544 12860
rect 23480 12844 23532 12850
rect 23308 12804 23480 12832
rect 23308 12442 23336 12804
rect 23480 12786 23532 12792
rect 23572 12776 23624 12782
rect 23400 12724 23572 12730
rect 23400 12718 23624 12724
rect 23400 12702 23612 12718
rect 23664 12708 23716 12714
rect 23400 12481 23428 12702
rect 23664 12650 23716 12656
rect 23386 12472 23442 12481
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 23296 12436 23348 12442
rect 23386 12407 23442 12416
rect 23296 12378 23348 12384
rect 23216 12306 23244 12378
rect 23204 12300 23256 12306
rect 23204 12242 23256 12248
rect 23204 12164 23256 12170
rect 23204 12106 23256 12112
rect 23216 11626 23244 12106
rect 23204 11620 23256 11626
rect 23204 11562 23256 11568
rect 23204 11280 23256 11286
rect 23308 11234 23336 12378
rect 23400 11694 23428 12407
rect 23676 12170 23704 12650
rect 23768 12238 23796 12854
rect 24110 12540 24418 12560
rect 24110 12538 24116 12540
rect 24172 12538 24196 12540
rect 24252 12538 24276 12540
rect 24332 12538 24356 12540
rect 24412 12538 24418 12540
rect 24172 12486 24174 12538
rect 24354 12486 24356 12538
rect 24110 12484 24116 12486
rect 24172 12484 24196 12486
rect 24252 12484 24276 12486
rect 24332 12484 24356 12486
rect 24412 12484 24418 12486
rect 24110 12464 24418 12484
rect 24780 12434 24808 14447
rect 24872 14346 24900 15370
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 25056 14414 25084 14758
rect 25148 14618 25176 16662
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25240 15910 25268 16526
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25240 14890 25268 15846
rect 25228 14884 25280 14890
rect 25228 14826 25280 14832
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 24860 14340 24912 14346
rect 24860 14282 24912 14288
rect 25044 14272 25096 14278
rect 25044 14214 25096 14220
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24872 12646 24900 13806
rect 25056 13734 25084 14214
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 25056 13394 25084 13670
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 25056 12986 25084 13330
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25148 12866 25176 14554
rect 25332 13258 25360 17138
rect 25700 16998 25728 17546
rect 25884 17542 25912 18226
rect 26160 18170 26188 21490
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26344 21078 26372 21286
rect 26332 21072 26384 21078
rect 26332 21014 26384 21020
rect 26344 20262 26372 21014
rect 26436 20330 26464 21490
rect 26528 20602 26556 21830
rect 26608 20936 26660 20942
rect 26608 20878 26660 20884
rect 26516 20596 26568 20602
rect 26516 20538 26568 20544
rect 26424 20324 26476 20330
rect 26424 20266 26476 20272
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26344 19922 26372 20198
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 26240 19712 26292 19718
rect 26240 19654 26292 19660
rect 26252 19514 26280 19654
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26344 19378 26372 19858
rect 26620 19854 26648 20878
rect 26608 19848 26660 19854
rect 26712 19825 26740 26250
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27264 22234 27292 22578
rect 27252 22228 27304 22234
rect 27252 22170 27304 22176
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 26884 20936 26936 20942
rect 26884 20878 26936 20884
rect 26792 20460 26844 20466
rect 26792 20402 26844 20408
rect 26804 20058 26832 20402
rect 26896 20398 26924 20878
rect 26884 20392 26936 20398
rect 26884 20334 26936 20340
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26608 19790 26660 19796
rect 26698 19816 26754 19825
rect 26424 19780 26476 19786
rect 26698 19751 26754 19760
rect 26424 19722 26476 19728
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 26252 18970 26280 19110
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 26436 18850 26464 19722
rect 26514 19408 26570 19417
rect 26514 19343 26516 19352
rect 26568 19343 26570 19352
rect 26516 19314 26568 19320
rect 26896 19242 26924 20334
rect 27080 19514 27108 21966
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 26884 19236 26936 19242
rect 26884 19178 26936 19184
rect 26068 18142 26188 18170
rect 26252 18822 26464 18850
rect 25964 18080 26016 18086
rect 25964 18022 26016 18028
rect 25976 17678 26004 18022
rect 25964 17672 26016 17678
rect 25964 17614 26016 17620
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 25780 17264 25832 17270
rect 25780 17206 25832 17212
rect 25412 16992 25464 16998
rect 25412 16934 25464 16940
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25424 16794 25452 16934
rect 25412 16788 25464 16794
rect 25412 16730 25464 16736
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 25412 16040 25464 16046
rect 25412 15982 25464 15988
rect 25424 14521 25452 15982
rect 25516 15706 25544 16390
rect 25792 16114 25820 17206
rect 26068 17134 26096 18142
rect 26252 17678 26280 18822
rect 26332 18760 26384 18766
rect 26332 18702 26384 18708
rect 26344 18290 26372 18702
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26332 18284 26384 18290
rect 26332 18226 26384 18232
rect 26436 18086 26464 18566
rect 26424 18080 26476 18086
rect 26424 18022 26476 18028
rect 26436 17678 26464 18022
rect 26896 17678 26924 19178
rect 27068 18896 27120 18902
rect 27068 18838 27120 18844
rect 26240 17672 26292 17678
rect 26240 17614 26292 17620
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26884 17672 26936 17678
rect 26884 17614 26936 17620
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 26160 16590 26188 16934
rect 26240 16720 26292 16726
rect 26240 16662 26292 16668
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26252 16114 26280 16662
rect 26344 16590 26372 17478
rect 26436 17338 26464 17614
rect 26424 17332 26476 17338
rect 26424 17274 26476 17280
rect 26424 17060 26476 17066
rect 26424 17002 26476 17008
rect 26332 16584 26384 16590
rect 26332 16526 26384 16532
rect 26436 16522 26464 17002
rect 26896 16590 26924 17614
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26424 16516 26476 16522
rect 26424 16458 26476 16464
rect 26896 16182 26924 16526
rect 26884 16176 26936 16182
rect 26884 16118 26936 16124
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 25504 15700 25556 15706
rect 25504 15642 25556 15648
rect 25410 14512 25466 14521
rect 25516 14482 25544 15642
rect 26160 15570 26188 16050
rect 26884 16040 26936 16046
rect 26884 15982 26936 15988
rect 26896 15706 26924 15982
rect 26884 15700 26936 15706
rect 26884 15642 26936 15648
rect 26792 15632 26844 15638
rect 26792 15574 26844 15580
rect 26148 15564 26200 15570
rect 26148 15506 26200 15512
rect 26516 15496 26568 15502
rect 26516 15438 26568 15444
rect 25596 15428 25648 15434
rect 25596 15370 25648 15376
rect 26056 15428 26108 15434
rect 26056 15370 26108 15376
rect 25608 14958 25636 15370
rect 26068 15026 26096 15370
rect 26056 15020 26108 15026
rect 26056 14962 26108 14968
rect 25596 14952 25648 14958
rect 25596 14894 25648 14900
rect 25872 14884 25924 14890
rect 25872 14826 25924 14832
rect 25410 14447 25466 14456
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25884 14346 25912 14826
rect 26068 14618 26096 14962
rect 26148 14952 26200 14958
rect 26148 14894 26200 14900
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 25872 14340 25924 14346
rect 25872 14282 25924 14288
rect 25504 14272 25556 14278
rect 25502 14240 25504 14249
rect 25556 14240 25558 14249
rect 25502 14175 25558 14184
rect 25884 14074 25912 14282
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 25688 13796 25740 13802
rect 25688 13738 25740 13744
rect 25700 13297 25728 13738
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 25872 13320 25924 13326
rect 25686 13288 25742 13297
rect 25320 13252 25372 13258
rect 25872 13262 25924 13268
rect 25686 13223 25688 13232
rect 25320 13194 25372 13200
rect 25740 13223 25742 13232
rect 25688 13194 25740 13200
rect 25056 12838 25176 12866
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 23952 12406 24808 12434
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 23664 12164 23716 12170
rect 23664 12106 23716 12112
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23388 11688 23440 11694
rect 23388 11630 23440 11636
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23492 11506 23520 11630
rect 23256 11228 23336 11234
rect 23204 11222 23336 11228
rect 23216 11206 23336 11222
rect 23400 11478 23520 11506
rect 23400 11218 23428 11478
rect 23388 11212 23440 11218
rect 23388 11154 23440 11160
rect 22704 11104 22784 11132
rect 23112 11144 23164 11150
rect 22652 11086 22704 11092
rect 23112 11086 23164 11092
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 22376 10736 22428 10742
rect 22376 10678 22428 10684
rect 23308 10470 23336 11086
rect 23400 10810 23428 11154
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23296 10464 23348 10470
rect 23296 10406 23348 10412
rect 23308 10130 23336 10406
rect 23584 10198 23612 12038
rect 23768 11762 23796 12174
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 23860 11898 23888 12038
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 23662 11656 23718 11665
rect 23662 11591 23718 11600
rect 23572 10192 23624 10198
rect 23572 10134 23624 10140
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 22468 9920 22520 9926
rect 22468 9862 22520 9868
rect 22480 9722 22508 9862
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22296 8566 22324 9522
rect 22376 9512 22428 9518
rect 22376 9454 22428 9460
rect 22388 9110 22416 9454
rect 22376 9104 22428 9110
rect 22376 9046 22428 9052
rect 22388 8838 22416 9046
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 23308 8566 23336 10066
rect 23572 9988 23624 9994
rect 23572 9930 23624 9936
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23492 9450 23520 9862
rect 23480 9444 23532 9450
rect 23480 9386 23532 9392
rect 23492 9042 23520 9386
rect 23584 9178 23612 9930
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 22284 8560 22336 8566
rect 22284 8502 22336 8508
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22744 8424 22796 8430
rect 22744 8366 22796 8372
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22112 7546 22140 7754
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 21364 7472 21416 7478
rect 21364 7414 21416 7420
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22204 7002 22232 7346
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22192 6996 22244 7002
rect 22192 6938 22244 6944
rect 22388 6798 22416 7142
rect 22756 6866 22784 8366
rect 22836 8288 22888 8294
rect 22836 8230 22888 8236
rect 22848 7342 22876 8230
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 22848 6934 22876 7278
rect 22836 6928 22888 6934
rect 22836 6870 22888 6876
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 20824 6458 20852 6598
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 19892 5636 19944 5642
rect 19892 5578 19944 5584
rect 19478 5468 19786 5488
rect 19478 5466 19484 5468
rect 19540 5466 19564 5468
rect 19620 5466 19644 5468
rect 19700 5466 19724 5468
rect 19780 5466 19786 5468
rect 19540 5414 19542 5466
rect 19722 5414 19724 5466
rect 19478 5412 19484 5414
rect 19540 5412 19564 5414
rect 19620 5412 19644 5414
rect 19700 5412 19724 5414
rect 19780 5412 19786 5414
rect 19478 5392 19786 5412
rect 20364 5302 20392 5714
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 20456 5098 20484 6258
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20640 5234 20668 6054
rect 21100 5710 21128 6190
rect 22112 5914 22140 6598
rect 22664 6254 22692 6598
rect 22652 6248 22704 6254
rect 22652 6190 22704 6196
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 20824 5370 20852 5578
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 22112 5302 22140 5850
rect 22204 5370 22232 6054
rect 22664 5914 22692 6190
rect 22652 5908 22704 5914
rect 22652 5850 22704 5856
rect 22756 5710 22784 6802
rect 22848 6254 22876 6870
rect 23676 6798 23704 11591
rect 23860 11354 23888 11834
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23952 10062 23980 12406
rect 24584 12368 24636 12374
rect 24584 12310 24636 12316
rect 24492 12164 24544 12170
rect 24492 12106 24544 12112
rect 24032 11756 24084 11762
rect 24032 11698 24084 11704
rect 24044 11558 24072 11698
rect 24032 11552 24084 11558
rect 24032 11494 24084 11500
rect 24044 11286 24072 11494
rect 24110 11452 24418 11472
rect 24110 11450 24116 11452
rect 24172 11450 24196 11452
rect 24252 11450 24276 11452
rect 24332 11450 24356 11452
rect 24412 11450 24418 11452
rect 24172 11398 24174 11450
rect 24354 11398 24356 11450
rect 24110 11396 24116 11398
rect 24172 11396 24196 11398
rect 24252 11396 24276 11398
rect 24332 11396 24356 11398
rect 24412 11396 24418 11398
rect 24110 11376 24418 11396
rect 24032 11280 24084 11286
rect 24032 11222 24084 11228
rect 24504 11082 24532 12106
rect 24032 11076 24084 11082
rect 24032 11018 24084 11024
rect 24492 11076 24544 11082
rect 24492 11018 24544 11024
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 24044 9994 24072 11018
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24110 10364 24418 10384
rect 24110 10362 24116 10364
rect 24172 10362 24196 10364
rect 24252 10362 24276 10364
rect 24332 10362 24356 10364
rect 24412 10362 24418 10364
rect 24172 10310 24174 10362
rect 24354 10310 24356 10362
rect 24110 10308 24116 10310
rect 24172 10308 24196 10310
rect 24252 10308 24276 10310
rect 24332 10308 24356 10310
rect 24412 10308 24418 10310
rect 24110 10288 24418 10308
rect 24032 9988 24084 9994
rect 24032 9930 24084 9936
rect 23848 9920 23900 9926
rect 23848 9862 23900 9868
rect 23860 8498 23888 9862
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 24044 8634 24072 9522
rect 24110 9276 24418 9296
rect 24110 9274 24116 9276
rect 24172 9274 24196 9276
rect 24252 9274 24276 9276
rect 24332 9274 24356 9276
rect 24412 9274 24418 9276
rect 24172 9222 24174 9274
rect 24354 9222 24356 9274
rect 24110 9220 24116 9222
rect 24172 9220 24196 9222
rect 24252 9220 24276 9222
rect 24332 9220 24356 9222
rect 24412 9220 24418 9222
rect 24110 9200 24418 9220
rect 24032 8628 24084 8634
rect 24032 8570 24084 8576
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 24110 8188 24418 8208
rect 24110 8186 24116 8188
rect 24172 8186 24196 8188
rect 24252 8186 24276 8188
rect 24332 8186 24356 8188
rect 24412 8186 24418 8188
rect 24172 8134 24174 8186
rect 24354 8134 24356 8186
rect 24110 8132 24116 8134
rect 24172 8132 24196 8134
rect 24252 8132 24276 8134
rect 24332 8132 24356 8134
rect 24412 8132 24418 8134
rect 24110 8112 24418 8132
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 24044 7546 24072 7958
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 24110 7100 24418 7120
rect 24110 7098 24116 7100
rect 24172 7098 24196 7100
rect 24252 7098 24276 7100
rect 24332 7098 24356 7100
rect 24412 7098 24418 7100
rect 24172 7046 24174 7098
rect 24354 7046 24356 7098
rect 24110 7044 24116 7046
rect 24172 7044 24196 7046
rect 24252 7044 24276 7046
rect 24332 7044 24356 7046
rect 24412 7044 24418 7046
rect 24110 7024 24418 7044
rect 24504 6882 24532 10746
rect 24596 10674 24624 12310
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24688 11354 24716 12174
rect 24768 12164 24820 12170
rect 24768 12106 24820 12112
rect 24780 11830 24808 12106
rect 24872 11898 24900 12582
rect 25056 12306 25084 12838
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 25240 12442 25268 12718
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 25240 12170 25268 12378
rect 25228 12164 25280 12170
rect 25228 12106 25280 12112
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24768 11824 24820 11830
rect 24964 11778 24992 12038
rect 24768 11766 24820 11772
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 24688 10810 24716 11154
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24688 9382 24716 10066
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 24688 8906 24716 9318
rect 24780 8974 24808 11766
rect 24872 11750 24992 11778
rect 24872 11014 24900 11750
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24860 11008 24912 11014
rect 24860 10950 24912 10956
rect 24872 9994 24900 10950
rect 24964 10810 24992 11494
rect 25240 11150 25268 12106
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 25240 10742 25268 11086
rect 25332 11082 25360 13194
rect 25884 12986 25912 13262
rect 25976 13258 26004 13670
rect 26160 13394 26188 14894
rect 26528 14414 26556 15438
rect 26804 15366 26832 15574
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 26792 15088 26844 15094
rect 26792 15030 26844 15036
rect 26804 14414 26832 15030
rect 26988 14414 27016 15302
rect 27080 14414 27108 18838
rect 27356 18358 27384 27270
rect 27540 26586 27568 28591
rect 28092 27606 28120 29294
rect 28998 29200 29054 30000
rect 28080 27600 28132 27606
rect 28080 27542 28132 27548
rect 27896 27464 27948 27470
rect 27896 27406 27948 27412
rect 27908 27130 27936 27406
rect 27896 27124 27948 27130
rect 27896 27066 27948 27072
rect 28356 26784 28408 26790
rect 28356 26726 28408 26732
rect 27528 26580 27580 26586
rect 27528 26522 27580 26528
rect 28368 26382 28396 26726
rect 28356 26376 28408 26382
rect 28356 26318 28408 26324
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 28276 24585 28304 24754
rect 28262 24576 28318 24585
rect 28262 24511 28318 24520
rect 28264 23724 28316 23730
rect 28264 23666 28316 23672
rect 27988 23588 28040 23594
rect 27988 23530 28040 23536
rect 27802 19000 27858 19009
rect 27802 18935 27804 18944
rect 27856 18935 27858 18944
rect 27804 18906 27856 18912
rect 27344 18352 27396 18358
rect 27344 18294 27396 18300
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27264 14618 27292 14962
rect 27252 14612 27304 14618
rect 27252 14554 27304 14560
rect 26516 14408 26568 14414
rect 26516 14350 26568 14356
rect 26792 14408 26844 14414
rect 26792 14350 26844 14356
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 26344 14006 26372 14214
rect 26804 14074 26832 14350
rect 26792 14068 26844 14074
rect 26792 14010 26844 14016
rect 26332 14000 26384 14006
rect 26332 13942 26384 13948
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26976 13932 27028 13938
rect 26976 13874 27028 13880
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 26160 12782 26188 13330
rect 26148 12776 26200 12782
rect 26148 12718 26200 12724
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25516 11354 25544 11698
rect 25700 11694 25728 12174
rect 26148 12096 26200 12102
rect 26148 12038 26200 12044
rect 25688 11688 25740 11694
rect 25688 11630 25740 11636
rect 25504 11348 25556 11354
rect 25504 11290 25556 11296
rect 26160 11082 26188 12038
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 25332 10742 25360 11018
rect 26252 10810 26280 13874
rect 26988 13530 27016 13874
rect 27080 13870 27108 14350
rect 27896 14340 27948 14346
rect 27896 14282 27948 14288
rect 27908 14006 27936 14282
rect 28000 14113 28028 23530
rect 28276 23225 28304 23666
rect 28262 23216 28318 23225
rect 28262 23151 28318 23160
rect 28356 22160 28408 22166
rect 28356 22102 28408 22108
rect 28368 21865 28396 22102
rect 28354 21856 28410 21865
rect 28354 21791 28410 21800
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 28368 20505 28396 21286
rect 28354 20496 28410 20505
rect 28354 20431 28410 20440
rect 28356 19848 28408 19854
rect 28356 19790 28408 19796
rect 28172 19168 28224 19174
rect 28368 19145 28396 19790
rect 28172 19110 28224 19116
rect 28354 19136 28410 19145
rect 28184 18970 28212 19110
rect 28354 19071 28410 19080
rect 28172 18964 28224 18970
rect 28172 18906 28224 18912
rect 28080 18760 28132 18766
rect 28080 18702 28132 18708
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28092 18290 28120 18702
rect 28080 18284 28132 18290
rect 28080 18226 28132 18232
rect 28092 17882 28120 18226
rect 28172 18080 28224 18086
rect 28172 18022 28224 18028
rect 28080 17876 28132 17882
rect 28080 17818 28132 17824
rect 28184 17785 28212 18022
rect 28170 17776 28226 17785
rect 28170 17711 28226 17720
rect 28170 17640 28226 17649
rect 28170 17575 28226 17584
rect 28184 17338 28212 17575
rect 28172 17332 28224 17338
rect 28172 17274 28224 17280
rect 28276 17270 28304 18702
rect 28448 18284 28500 18290
rect 28448 18226 28500 18232
rect 28264 17264 28316 17270
rect 28264 17206 28316 17212
rect 28276 16794 28304 17206
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 28264 16788 28316 16794
rect 28264 16730 28316 16736
rect 28368 16425 28396 17138
rect 28354 16416 28410 16425
rect 28354 16351 28410 16360
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28368 15570 28396 15846
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 27986 14104 28042 14113
rect 27986 14039 28042 14048
rect 27896 14000 27948 14006
rect 27896 13942 27948 13948
rect 27068 13864 27120 13870
rect 27068 13806 27120 13812
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 27172 12918 27200 13670
rect 27252 13252 27304 13258
rect 27252 13194 27304 13200
rect 27160 12912 27212 12918
rect 27160 12854 27212 12860
rect 27066 12744 27122 12753
rect 27066 12679 27122 12688
rect 27080 12238 27108 12679
rect 27264 12442 27292 13194
rect 27908 12986 27936 13942
rect 28276 13938 28304 15302
rect 28356 14816 28408 14822
rect 28356 14758 28408 14764
rect 28368 14414 28396 14758
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 28264 13932 28316 13938
rect 28264 13874 28316 13880
rect 28276 13705 28304 13874
rect 28262 13696 28318 13705
rect 28262 13631 28318 13640
rect 28460 13530 28488 18226
rect 28448 13524 28500 13530
rect 28448 13466 28500 13472
rect 27896 12980 27948 12986
rect 27896 12922 27948 12928
rect 27252 12436 27304 12442
rect 27252 12378 27304 12384
rect 28354 12336 28410 12345
rect 28354 12271 28356 12280
rect 28408 12271 28410 12280
rect 28356 12242 28408 12248
rect 27068 12232 27120 12238
rect 27068 12174 27120 12180
rect 28356 11144 28408 11150
rect 28356 11086 28408 11092
rect 28368 10985 28396 11086
rect 28354 10976 28410 10985
rect 28354 10911 28410 10920
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 25228 10736 25280 10742
rect 25228 10678 25280 10684
rect 25320 10736 25372 10742
rect 25320 10678 25372 10684
rect 25780 10668 25832 10674
rect 25780 10610 25832 10616
rect 25792 10266 25820 10610
rect 26252 10470 26280 10746
rect 26792 10668 26844 10674
rect 26792 10610 26844 10616
rect 26240 10464 26292 10470
rect 26240 10406 26292 10412
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 26804 10198 26832 10610
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 26792 10192 26844 10198
rect 26792 10134 26844 10140
rect 27356 10062 27384 10406
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24872 9042 24900 9930
rect 25148 9042 25176 9998
rect 25332 9178 25360 9998
rect 25504 9920 25556 9926
rect 25504 9862 25556 9868
rect 26516 9920 26568 9926
rect 26516 9862 26568 9868
rect 28080 9920 28132 9926
rect 28080 9862 28132 9868
rect 25516 9654 25544 9862
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 26528 9450 26556 9862
rect 26516 9444 26568 9450
rect 26516 9386 26568 9392
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 26528 9110 26556 9386
rect 26516 9104 26568 9110
rect 26516 9046 26568 9052
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 25136 9036 25188 9042
rect 25136 8978 25188 8984
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24676 8900 24728 8906
rect 24676 8842 24728 8848
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24596 8022 24624 8366
rect 24584 8016 24636 8022
rect 24584 7958 24636 7964
rect 24688 7886 24716 8842
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24504 6854 24624 6882
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 24492 6792 24544 6798
rect 24492 6734 24544 6740
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23676 6322 23704 6598
rect 24504 6458 24532 6734
rect 24596 6730 24624 6854
rect 24584 6724 24636 6730
rect 24584 6666 24636 6672
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24688 6390 24716 7822
rect 24964 7546 24992 8434
rect 25148 8430 25176 8978
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 25412 7744 25464 7750
rect 25412 7686 25464 7692
rect 25424 7546 25452 7686
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24872 6866 24900 7346
rect 25608 7342 25636 8910
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 25792 7546 25820 8774
rect 26516 8356 26568 8362
rect 26516 8298 26568 8304
rect 26528 7886 26556 8298
rect 26516 7880 26568 7886
rect 26516 7822 26568 7828
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 25596 7336 25648 7342
rect 25596 7278 25648 7284
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24872 6458 24900 6802
rect 24860 6452 24912 6458
rect 24860 6394 24912 6400
rect 24676 6384 24728 6390
rect 24676 6326 24728 6332
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22100 5296 22152 5302
rect 22100 5238 22152 5244
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 22296 5166 22324 5646
rect 23216 5370 23244 6258
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 23308 5710 23336 6054
rect 23768 5778 23796 6258
rect 24110 6012 24418 6032
rect 24110 6010 24116 6012
rect 24172 6010 24196 6012
rect 24252 6010 24276 6012
rect 24332 6010 24356 6012
rect 24412 6010 24418 6012
rect 24172 5958 24174 6010
rect 24354 5958 24356 6010
rect 24110 5956 24116 5958
rect 24172 5956 24196 5958
rect 24252 5956 24276 5958
rect 24332 5956 24356 5958
rect 24412 5956 24418 5958
rect 24110 5936 24418 5956
rect 23756 5772 23808 5778
rect 23756 5714 23808 5720
rect 28092 5710 28120 9862
rect 28262 9616 28318 9625
rect 28262 9551 28264 9560
rect 28316 9551 28318 9560
rect 28264 9522 28316 9528
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28172 8288 28224 8294
rect 28368 8265 28396 8434
rect 28172 8230 28224 8236
rect 28354 8256 28410 8265
rect 28184 8090 28212 8230
rect 28354 8191 28410 8200
rect 28172 8084 28224 8090
rect 28172 8026 28224 8032
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 28184 6730 28212 7142
rect 28368 6905 28396 7346
rect 28354 6896 28410 6905
rect 28354 6831 28410 6840
rect 28172 6724 28224 6730
rect 28172 6666 28224 6672
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 28264 5568 28316 5574
rect 28262 5536 28264 5545
rect 28316 5536 28318 5545
rect 28262 5471 28318 5480
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 20444 5092 20496 5098
rect 20444 5034 20496 5040
rect 24110 4924 24418 4944
rect 24110 4922 24116 4924
rect 24172 4922 24196 4924
rect 24252 4922 24276 4924
rect 24332 4922 24356 4924
rect 24412 4922 24418 4924
rect 24172 4870 24174 4922
rect 24354 4870 24356 4922
rect 24110 4868 24116 4870
rect 24172 4868 24196 4870
rect 24252 4868 24276 4870
rect 24332 4868 24356 4870
rect 24412 4868 24418 4870
rect 24110 4848 24418 4868
rect 28356 4616 28408 4622
rect 28356 4558 28408 4564
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 19478 4380 19786 4400
rect 19478 4378 19484 4380
rect 19540 4378 19564 4380
rect 19620 4378 19644 4380
rect 19700 4378 19724 4380
rect 19780 4378 19786 4380
rect 19540 4326 19542 4378
rect 19722 4326 19724 4378
rect 19478 4324 19484 4326
rect 19540 4324 19564 4326
rect 19620 4324 19644 4326
rect 19700 4324 19724 4326
rect 19780 4324 19786 4326
rect 19478 4304 19786 4324
rect 28368 4185 28396 4558
rect 28354 4176 28410 4185
rect 28354 4111 28410 4120
rect 24110 3836 24418 3856
rect 24110 3834 24116 3836
rect 24172 3834 24196 3836
rect 24252 3834 24276 3836
rect 24332 3834 24356 3836
rect 24412 3834 24418 3836
rect 24172 3782 24174 3834
rect 24354 3782 24356 3834
rect 24110 3780 24116 3782
rect 24172 3780 24196 3782
rect 24252 3780 24276 3782
rect 24332 3780 24356 3782
rect 24412 3780 24418 3782
rect 24110 3760 24418 3780
rect 19478 3292 19786 3312
rect 19478 3290 19484 3292
rect 19540 3290 19564 3292
rect 19620 3290 19644 3292
rect 19700 3290 19724 3292
rect 19780 3290 19786 3292
rect 19540 3238 19542 3290
rect 19722 3238 19724 3290
rect 19478 3236 19484 3238
rect 19540 3236 19564 3238
rect 19620 3236 19644 3238
rect 19700 3236 19724 3238
rect 19780 3236 19786 3238
rect 19478 3216 19786 3236
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24110 2748 24418 2768
rect 24110 2746 24116 2748
rect 24172 2746 24196 2748
rect 24252 2746 24276 2748
rect 24332 2746 24356 2748
rect 24412 2746 24418 2748
rect 24172 2694 24174 2746
rect 24354 2694 24356 2746
rect 24110 2692 24116 2694
rect 24172 2692 24196 2694
rect 24252 2692 24276 2694
rect 24332 2692 24356 2694
rect 24412 2692 24418 2694
rect 24110 2672 24418 2692
rect 24596 2650 24624 2994
rect 28356 2848 28408 2854
rect 28354 2816 28356 2825
rect 28408 2816 28410 2825
rect 28354 2751 28410 2760
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 27528 2440 27580 2446
rect 27528 2382 27580 2388
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 10214 2204 10522 2224
rect 10214 2202 10220 2204
rect 10276 2202 10300 2204
rect 10356 2202 10380 2204
rect 10436 2202 10460 2204
rect 10516 2202 10522 2204
rect 10276 2150 10278 2202
rect 10458 2150 10460 2202
rect 10214 2148 10220 2150
rect 10276 2148 10300 2150
rect 10356 2148 10380 2150
rect 10436 2148 10460 2150
rect 10516 2148 10522 2150
rect 10214 2128 10522 2148
rect 10152 1278 10364 1306
rect 10336 800 10364 1278
rect 15488 800 15516 2382
rect 18064 800 18092 2382
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 19478 2204 19786 2224
rect 19478 2202 19484 2204
rect 19540 2202 19564 2204
rect 19620 2202 19644 2204
rect 19700 2202 19724 2204
rect 19780 2202 19786 2204
rect 19540 2150 19542 2202
rect 19722 2150 19724 2202
rect 19478 2148 19484 2150
rect 19540 2148 19564 2150
rect 19620 2148 19644 2150
rect 19700 2148 19724 2150
rect 19780 2148 19786 2150
rect 19478 2128 19786 2148
rect 20640 800 20668 2246
rect 24504 800 24532 2382
rect 25792 800 25820 2382
rect 27080 800 27108 2382
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 27540 105 27568 2382
rect 27526 96 27582 105
rect 27526 31 27582 40
rect 28354 0 28410 800
<< via2 >>
rect 1398 28600 1454 28656
rect 5588 27770 5644 27772
rect 5668 27770 5724 27772
rect 5748 27770 5804 27772
rect 5828 27770 5884 27772
rect 5588 27718 5634 27770
rect 5634 27718 5644 27770
rect 5668 27718 5698 27770
rect 5698 27718 5710 27770
rect 5710 27718 5724 27770
rect 5748 27718 5762 27770
rect 5762 27718 5774 27770
rect 5774 27718 5804 27770
rect 5828 27718 5838 27770
rect 5838 27718 5884 27770
rect 5588 27716 5644 27718
rect 5668 27716 5724 27718
rect 5748 27716 5804 27718
rect 5828 27716 5884 27718
rect 14852 27770 14908 27772
rect 14932 27770 14988 27772
rect 15012 27770 15068 27772
rect 15092 27770 15148 27772
rect 14852 27718 14898 27770
rect 14898 27718 14908 27770
rect 14932 27718 14962 27770
rect 14962 27718 14974 27770
rect 14974 27718 14988 27770
rect 15012 27718 15026 27770
rect 15026 27718 15038 27770
rect 15038 27718 15068 27770
rect 15092 27718 15102 27770
rect 15102 27718 15148 27770
rect 14852 27716 14908 27718
rect 14932 27716 14988 27718
rect 15012 27716 15068 27718
rect 15092 27716 15148 27718
rect 1398 27240 1454 27296
rect 1398 23160 1454 23216
rect 1398 21800 1454 21856
rect 1398 17756 1400 17776
rect 1400 17756 1452 17776
rect 1452 17756 1454 17776
rect 1398 17720 1454 17756
rect 1398 16360 1454 16416
rect 1398 10920 1454 10976
rect 1674 25880 1730 25936
rect 1582 9560 1638 9616
rect 1582 8200 1638 8256
rect 1398 4120 1454 4176
rect 1490 2796 1492 2816
rect 1492 2796 1544 2816
rect 1544 2796 1546 2816
rect 1490 2760 1546 2796
rect 10220 27226 10276 27228
rect 10300 27226 10356 27228
rect 10380 27226 10436 27228
rect 10460 27226 10516 27228
rect 10220 27174 10266 27226
rect 10266 27174 10276 27226
rect 10300 27174 10330 27226
rect 10330 27174 10342 27226
rect 10342 27174 10356 27226
rect 10380 27174 10394 27226
rect 10394 27174 10406 27226
rect 10406 27174 10436 27226
rect 10460 27174 10470 27226
rect 10470 27174 10516 27226
rect 10220 27172 10276 27174
rect 10300 27172 10356 27174
rect 10380 27172 10436 27174
rect 10460 27172 10516 27174
rect 5588 26682 5644 26684
rect 5668 26682 5724 26684
rect 5748 26682 5804 26684
rect 5828 26682 5884 26684
rect 5588 26630 5634 26682
rect 5634 26630 5644 26682
rect 5668 26630 5698 26682
rect 5698 26630 5710 26682
rect 5710 26630 5724 26682
rect 5748 26630 5762 26682
rect 5762 26630 5774 26682
rect 5774 26630 5804 26682
rect 5828 26630 5838 26682
rect 5838 26630 5884 26682
rect 5588 26628 5644 26630
rect 5668 26628 5724 26630
rect 5748 26628 5804 26630
rect 5828 26628 5884 26630
rect 10220 26138 10276 26140
rect 10300 26138 10356 26140
rect 10380 26138 10436 26140
rect 10460 26138 10516 26140
rect 10220 26086 10266 26138
rect 10266 26086 10276 26138
rect 10300 26086 10330 26138
rect 10330 26086 10342 26138
rect 10342 26086 10356 26138
rect 10380 26086 10394 26138
rect 10394 26086 10406 26138
rect 10406 26086 10436 26138
rect 10460 26086 10470 26138
rect 10470 26086 10516 26138
rect 10220 26084 10276 26086
rect 10300 26084 10356 26086
rect 10380 26084 10436 26086
rect 10460 26084 10516 26086
rect 5588 25594 5644 25596
rect 5668 25594 5724 25596
rect 5748 25594 5804 25596
rect 5828 25594 5884 25596
rect 5588 25542 5634 25594
rect 5634 25542 5644 25594
rect 5668 25542 5698 25594
rect 5698 25542 5710 25594
rect 5710 25542 5724 25594
rect 5748 25542 5762 25594
rect 5762 25542 5774 25594
rect 5774 25542 5804 25594
rect 5828 25542 5838 25594
rect 5838 25542 5884 25594
rect 5588 25540 5644 25542
rect 5668 25540 5724 25542
rect 5748 25540 5804 25542
rect 5828 25540 5884 25542
rect 10220 25050 10276 25052
rect 10300 25050 10356 25052
rect 10380 25050 10436 25052
rect 10460 25050 10516 25052
rect 10220 24998 10266 25050
rect 10266 24998 10276 25050
rect 10300 24998 10330 25050
rect 10330 24998 10342 25050
rect 10342 24998 10356 25050
rect 10380 24998 10394 25050
rect 10394 24998 10406 25050
rect 10406 24998 10436 25050
rect 10460 24998 10470 25050
rect 10470 24998 10516 25050
rect 10220 24996 10276 24998
rect 10300 24996 10356 24998
rect 10380 24996 10436 24998
rect 10460 24996 10516 24998
rect 5588 24506 5644 24508
rect 5668 24506 5724 24508
rect 5748 24506 5804 24508
rect 5828 24506 5884 24508
rect 5588 24454 5634 24506
rect 5634 24454 5644 24506
rect 5668 24454 5698 24506
rect 5698 24454 5710 24506
rect 5710 24454 5724 24506
rect 5748 24454 5762 24506
rect 5762 24454 5774 24506
rect 5774 24454 5804 24506
rect 5828 24454 5838 24506
rect 5838 24454 5884 24506
rect 5588 24452 5644 24454
rect 5668 24452 5724 24454
rect 5748 24452 5804 24454
rect 5828 24452 5884 24454
rect 10220 23962 10276 23964
rect 10300 23962 10356 23964
rect 10380 23962 10436 23964
rect 10460 23962 10516 23964
rect 10220 23910 10266 23962
rect 10266 23910 10276 23962
rect 10300 23910 10330 23962
rect 10330 23910 10342 23962
rect 10342 23910 10356 23962
rect 10380 23910 10394 23962
rect 10394 23910 10406 23962
rect 10406 23910 10436 23962
rect 10460 23910 10470 23962
rect 10470 23910 10516 23962
rect 10220 23908 10276 23910
rect 10300 23908 10356 23910
rect 10380 23908 10436 23910
rect 10460 23908 10516 23910
rect 5588 23418 5644 23420
rect 5668 23418 5724 23420
rect 5748 23418 5804 23420
rect 5828 23418 5884 23420
rect 5588 23366 5634 23418
rect 5634 23366 5644 23418
rect 5668 23366 5698 23418
rect 5698 23366 5710 23418
rect 5710 23366 5724 23418
rect 5748 23366 5762 23418
rect 5762 23366 5774 23418
rect 5774 23366 5804 23418
rect 5828 23366 5838 23418
rect 5838 23366 5884 23418
rect 5588 23364 5644 23366
rect 5668 23364 5724 23366
rect 5748 23364 5804 23366
rect 5828 23364 5884 23366
rect 10220 22874 10276 22876
rect 10300 22874 10356 22876
rect 10380 22874 10436 22876
rect 10460 22874 10516 22876
rect 10220 22822 10266 22874
rect 10266 22822 10276 22874
rect 10300 22822 10330 22874
rect 10330 22822 10342 22874
rect 10342 22822 10356 22874
rect 10380 22822 10394 22874
rect 10394 22822 10406 22874
rect 10406 22822 10436 22874
rect 10460 22822 10470 22874
rect 10470 22822 10516 22874
rect 10220 22820 10276 22822
rect 10300 22820 10356 22822
rect 10380 22820 10436 22822
rect 10460 22820 10516 22822
rect 5588 22330 5644 22332
rect 5668 22330 5724 22332
rect 5748 22330 5804 22332
rect 5828 22330 5884 22332
rect 5588 22278 5634 22330
rect 5634 22278 5644 22330
rect 5668 22278 5698 22330
rect 5698 22278 5710 22330
rect 5710 22278 5724 22330
rect 5748 22278 5762 22330
rect 5762 22278 5774 22330
rect 5774 22278 5804 22330
rect 5828 22278 5838 22330
rect 5838 22278 5884 22330
rect 5588 22276 5644 22278
rect 5668 22276 5724 22278
rect 5748 22276 5804 22278
rect 5828 22276 5884 22278
rect 10220 21786 10276 21788
rect 10300 21786 10356 21788
rect 10380 21786 10436 21788
rect 10460 21786 10516 21788
rect 10220 21734 10266 21786
rect 10266 21734 10276 21786
rect 10300 21734 10330 21786
rect 10330 21734 10342 21786
rect 10342 21734 10356 21786
rect 10380 21734 10394 21786
rect 10394 21734 10406 21786
rect 10406 21734 10436 21786
rect 10460 21734 10470 21786
rect 10470 21734 10516 21786
rect 10220 21732 10276 21734
rect 10300 21732 10356 21734
rect 10380 21732 10436 21734
rect 10460 21732 10516 21734
rect 5588 21242 5644 21244
rect 5668 21242 5724 21244
rect 5748 21242 5804 21244
rect 5828 21242 5884 21244
rect 5588 21190 5634 21242
rect 5634 21190 5644 21242
rect 5668 21190 5698 21242
rect 5698 21190 5710 21242
rect 5710 21190 5724 21242
rect 5748 21190 5762 21242
rect 5762 21190 5774 21242
rect 5774 21190 5804 21242
rect 5828 21190 5838 21242
rect 5838 21190 5884 21242
rect 5588 21188 5644 21190
rect 5668 21188 5724 21190
rect 5748 21188 5804 21190
rect 5828 21188 5884 21190
rect 10220 20698 10276 20700
rect 10300 20698 10356 20700
rect 10380 20698 10436 20700
rect 10460 20698 10516 20700
rect 10220 20646 10266 20698
rect 10266 20646 10276 20698
rect 10300 20646 10330 20698
rect 10330 20646 10342 20698
rect 10342 20646 10356 20698
rect 10380 20646 10394 20698
rect 10394 20646 10406 20698
rect 10406 20646 10436 20698
rect 10460 20646 10470 20698
rect 10470 20646 10516 20698
rect 10220 20644 10276 20646
rect 10300 20644 10356 20646
rect 10380 20644 10436 20646
rect 10460 20644 10516 20646
rect 5588 20154 5644 20156
rect 5668 20154 5724 20156
rect 5748 20154 5804 20156
rect 5828 20154 5884 20156
rect 5588 20102 5634 20154
rect 5634 20102 5644 20154
rect 5668 20102 5698 20154
rect 5698 20102 5710 20154
rect 5710 20102 5724 20154
rect 5748 20102 5762 20154
rect 5762 20102 5774 20154
rect 5774 20102 5804 20154
rect 5828 20102 5838 20154
rect 5838 20102 5884 20154
rect 5588 20100 5644 20102
rect 5668 20100 5724 20102
rect 5748 20100 5804 20102
rect 5828 20100 5884 20102
rect 5588 19066 5644 19068
rect 5668 19066 5724 19068
rect 5748 19066 5804 19068
rect 5828 19066 5884 19068
rect 5588 19014 5634 19066
rect 5634 19014 5644 19066
rect 5668 19014 5698 19066
rect 5698 19014 5710 19066
rect 5710 19014 5724 19066
rect 5748 19014 5762 19066
rect 5762 19014 5774 19066
rect 5774 19014 5804 19066
rect 5828 19014 5838 19066
rect 5838 19014 5884 19066
rect 5588 19012 5644 19014
rect 5668 19012 5724 19014
rect 5748 19012 5804 19014
rect 5828 19012 5884 19014
rect 5588 17978 5644 17980
rect 5668 17978 5724 17980
rect 5748 17978 5804 17980
rect 5828 17978 5884 17980
rect 5588 17926 5634 17978
rect 5634 17926 5644 17978
rect 5668 17926 5698 17978
rect 5698 17926 5710 17978
rect 5710 17926 5724 17978
rect 5748 17926 5762 17978
rect 5762 17926 5774 17978
rect 5774 17926 5804 17978
rect 5828 17926 5838 17978
rect 5838 17926 5884 17978
rect 5588 17924 5644 17926
rect 5668 17924 5724 17926
rect 5748 17924 5804 17926
rect 5828 17924 5884 17926
rect 5588 16890 5644 16892
rect 5668 16890 5724 16892
rect 5748 16890 5804 16892
rect 5828 16890 5884 16892
rect 5588 16838 5634 16890
rect 5634 16838 5644 16890
rect 5668 16838 5698 16890
rect 5698 16838 5710 16890
rect 5710 16838 5724 16890
rect 5748 16838 5762 16890
rect 5762 16838 5774 16890
rect 5774 16838 5804 16890
rect 5828 16838 5838 16890
rect 5838 16838 5884 16890
rect 5588 16836 5644 16838
rect 5668 16836 5724 16838
rect 5748 16836 5804 16838
rect 5828 16836 5884 16838
rect 5588 15802 5644 15804
rect 5668 15802 5724 15804
rect 5748 15802 5804 15804
rect 5828 15802 5884 15804
rect 5588 15750 5634 15802
rect 5634 15750 5644 15802
rect 5668 15750 5698 15802
rect 5698 15750 5710 15802
rect 5710 15750 5724 15802
rect 5748 15750 5762 15802
rect 5762 15750 5774 15802
rect 5774 15750 5804 15802
rect 5828 15750 5838 15802
rect 5838 15750 5884 15802
rect 5588 15748 5644 15750
rect 5668 15748 5724 15750
rect 5748 15748 5804 15750
rect 5828 15748 5884 15750
rect 4066 15000 4122 15056
rect 5588 14714 5644 14716
rect 5668 14714 5724 14716
rect 5748 14714 5804 14716
rect 5828 14714 5884 14716
rect 5588 14662 5634 14714
rect 5634 14662 5644 14714
rect 5668 14662 5698 14714
rect 5698 14662 5710 14714
rect 5710 14662 5724 14714
rect 5748 14662 5762 14714
rect 5762 14662 5774 14714
rect 5774 14662 5804 14714
rect 5828 14662 5838 14714
rect 5838 14662 5884 14714
rect 5588 14660 5644 14662
rect 5668 14660 5724 14662
rect 5748 14660 5804 14662
rect 5828 14660 5884 14662
rect 6550 14320 6606 14376
rect 5588 13626 5644 13628
rect 5668 13626 5724 13628
rect 5748 13626 5804 13628
rect 5828 13626 5884 13628
rect 5588 13574 5634 13626
rect 5634 13574 5644 13626
rect 5668 13574 5698 13626
rect 5698 13574 5710 13626
rect 5710 13574 5724 13626
rect 5748 13574 5762 13626
rect 5762 13574 5774 13626
rect 5774 13574 5804 13626
rect 5828 13574 5838 13626
rect 5838 13574 5884 13626
rect 5588 13572 5644 13574
rect 5668 13572 5724 13574
rect 5748 13572 5804 13574
rect 5828 13572 5884 13574
rect 10220 19610 10276 19612
rect 10300 19610 10356 19612
rect 10380 19610 10436 19612
rect 10460 19610 10516 19612
rect 10220 19558 10266 19610
rect 10266 19558 10276 19610
rect 10300 19558 10330 19610
rect 10330 19558 10342 19610
rect 10342 19558 10356 19610
rect 10380 19558 10394 19610
rect 10394 19558 10406 19610
rect 10406 19558 10436 19610
rect 10460 19558 10470 19610
rect 10470 19558 10516 19610
rect 10220 19556 10276 19558
rect 10300 19556 10356 19558
rect 10380 19556 10436 19558
rect 10460 19556 10516 19558
rect 10322 19252 10324 19272
rect 10324 19252 10376 19272
rect 10376 19252 10378 19272
rect 10322 19216 10378 19252
rect 9770 16632 9826 16688
rect 5588 12538 5644 12540
rect 5668 12538 5724 12540
rect 5748 12538 5804 12540
rect 5828 12538 5884 12540
rect 5588 12486 5634 12538
rect 5634 12486 5644 12538
rect 5668 12486 5698 12538
rect 5698 12486 5710 12538
rect 5710 12486 5724 12538
rect 5748 12486 5762 12538
rect 5762 12486 5774 12538
rect 5774 12486 5804 12538
rect 5828 12486 5838 12538
rect 5838 12486 5884 12538
rect 5588 12484 5644 12486
rect 5668 12484 5724 12486
rect 5748 12484 5804 12486
rect 5828 12484 5884 12486
rect 1766 12144 1822 12200
rect 8942 13776 8998 13832
rect 10220 18522 10276 18524
rect 10300 18522 10356 18524
rect 10380 18522 10436 18524
rect 10460 18522 10516 18524
rect 10220 18470 10266 18522
rect 10266 18470 10276 18522
rect 10300 18470 10330 18522
rect 10330 18470 10342 18522
rect 10342 18470 10356 18522
rect 10380 18470 10394 18522
rect 10394 18470 10406 18522
rect 10406 18470 10436 18522
rect 10460 18470 10470 18522
rect 10470 18470 10516 18522
rect 10220 18468 10276 18470
rect 10300 18468 10356 18470
rect 10380 18468 10436 18470
rect 10460 18468 10516 18470
rect 10782 18264 10838 18320
rect 10220 17434 10276 17436
rect 10300 17434 10356 17436
rect 10380 17434 10436 17436
rect 10460 17434 10516 17436
rect 10220 17382 10266 17434
rect 10266 17382 10276 17434
rect 10300 17382 10330 17434
rect 10330 17382 10342 17434
rect 10342 17382 10356 17434
rect 10380 17382 10394 17434
rect 10394 17382 10406 17434
rect 10406 17382 10436 17434
rect 10460 17382 10470 17434
rect 10470 17382 10516 17434
rect 10220 17380 10276 17382
rect 10300 17380 10356 17382
rect 10380 17380 10436 17382
rect 10460 17380 10516 17382
rect 10220 16346 10276 16348
rect 10300 16346 10356 16348
rect 10380 16346 10436 16348
rect 10460 16346 10516 16348
rect 10220 16294 10266 16346
rect 10266 16294 10276 16346
rect 10300 16294 10330 16346
rect 10330 16294 10342 16346
rect 10342 16294 10356 16346
rect 10380 16294 10394 16346
rect 10394 16294 10406 16346
rect 10406 16294 10436 16346
rect 10460 16294 10470 16346
rect 10470 16294 10516 16346
rect 10220 16292 10276 16294
rect 10300 16292 10356 16294
rect 10380 16292 10436 16294
rect 10460 16292 10516 16294
rect 10220 15258 10276 15260
rect 10300 15258 10356 15260
rect 10380 15258 10436 15260
rect 10460 15258 10516 15260
rect 10220 15206 10266 15258
rect 10266 15206 10276 15258
rect 10300 15206 10330 15258
rect 10330 15206 10342 15258
rect 10342 15206 10356 15258
rect 10380 15206 10394 15258
rect 10394 15206 10406 15258
rect 10406 15206 10436 15258
rect 10460 15206 10470 15258
rect 10470 15206 10516 15258
rect 10220 15204 10276 15206
rect 10300 15204 10356 15206
rect 10380 15204 10436 15206
rect 10460 15204 10516 15206
rect 10220 14170 10276 14172
rect 10300 14170 10356 14172
rect 10380 14170 10436 14172
rect 10460 14170 10516 14172
rect 10220 14118 10266 14170
rect 10266 14118 10276 14170
rect 10300 14118 10330 14170
rect 10330 14118 10342 14170
rect 10342 14118 10356 14170
rect 10380 14118 10394 14170
rect 10394 14118 10406 14170
rect 10406 14118 10436 14170
rect 10460 14118 10470 14170
rect 10470 14118 10516 14170
rect 10220 14116 10276 14118
rect 10300 14116 10356 14118
rect 10380 14116 10436 14118
rect 10460 14116 10516 14118
rect 10220 13082 10276 13084
rect 10300 13082 10356 13084
rect 10380 13082 10436 13084
rect 10460 13082 10516 13084
rect 10220 13030 10266 13082
rect 10266 13030 10276 13082
rect 10300 13030 10330 13082
rect 10330 13030 10342 13082
rect 10342 13030 10356 13082
rect 10380 13030 10394 13082
rect 10394 13030 10406 13082
rect 10406 13030 10436 13082
rect 10460 13030 10470 13082
rect 10470 13030 10516 13082
rect 10220 13028 10276 13030
rect 10300 13028 10356 13030
rect 10380 13028 10436 13030
rect 10460 13028 10516 13030
rect 5588 11450 5644 11452
rect 5668 11450 5724 11452
rect 5748 11450 5804 11452
rect 5828 11450 5884 11452
rect 5588 11398 5634 11450
rect 5634 11398 5644 11450
rect 5668 11398 5698 11450
rect 5698 11398 5710 11450
rect 5710 11398 5724 11450
rect 5748 11398 5762 11450
rect 5762 11398 5774 11450
rect 5774 11398 5804 11450
rect 5828 11398 5838 11450
rect 5838 11398 5884 11450
rect 5588 11396 5644 11398
rect 5668 11396 5724 11398
rect 5748 11396 5804 11398
rect 5828 11396 5884 11398
rect 5588 10362 5644 10364
rect 5668 10362 5724 10364
rect 5748 10362 5804 10364
rect 5828 10362 5884 10364
rect 5588 10310 5634 10362
rect 5634 10310 5644 10362
rect 5668 10310 5698 10362
rect 5698 10310 5710 10362
rect 5710 10310 5724 10362
rect 5748 10310 5762 10362
rect 5762 10310 5774 10362
rect 5774 10310 5804 10362
rect 5828 10310 5838 10362
rect 5838 10310 5884 10362
rect 5588 10308 5644 10310
rect 5668 10308 5724 10310
rect 5748 10308 5804 10310
rect 5828 10308 5884 10310
rect 5588 9274 5644 9276
rect 5668 9274 5724 9276
rect 5748 9274 5804 9276
rect 5828 9274 5884 9276
rect 5588 9222 5634 9274
rect 5634 9222 5644 9274
rect 5668 9222 5698 9274
rect 5698 9222 5710 9274
rect 5710 9222 5724 9274
rect 5748 9222 5762 9274
rect 5762 9222 5774 9274
rect 5774 9222 5804 9274
rect 5828 9222 5838 9274
rect 5838 9222 5884 9274
rect 5588 9220 5644 9222
rect 5668 9220 5724 9222
rect 5748 9220 5804 9222
rect 5828 9220 5884 9222
rect 9678 11192 9734 11248
rect 10220 11994 10276 11996
rect 10300 11994 10356 11996
rect 10380 11994 10436 11996
rect 10460 11994 10516 11996
rect 10220 11942 10266 11994
rect 10266 11942 10276 11994
rect 10300 11942 10330 11994
rect 10330 11942 10342 11994
rect 10342 11942 10356 11994
rect 10380 11942 10394 11994
rect 10394 11942 10406 11994
rect 10406 11942 10436 11994
rect 10460 11942 10470 11994
rect 10470 11942 10516 11994
rect 10220 11940 10276 11942
rect 10300 11940 10356 11942
rect 10380 11940 10436 11942
rect 10460 11940 10516 11942
rect 10220 10906 10276 10908
rect 10300 10906 10356 10908
rect 10380 10906 10436 10908
rect 10460 10906 10516 10908
rect 10220 10854 10266 10906
rect 10266 10854 10276 10906
rect 10300 10854 10330 10906
rect 10330 10854 10342 10906
rect 10342 10854 10356 10906
rect 10380 10854 10394 10906
rect 10394 10854 10406 10906
rect 10406 10854 10436 10906
rect 10460 10854 10470 10906
rect 10470 10854 10516 10906
rect 10220 10852 10276 10854
rect 10300 10852 10356 10854
rect 10380 10852 10436 10854
rect 10460 10852 10516 10854
rect 1766 8880 1822 8936
rect 5588 8186 5644 8188
rect 5668 8186 5724 8188
rect 5748 8186 5804 8188
rect 5828 8186 5884 8188
rect 5588 8134 5634 8186
rect 5634 8134 5644 8186
rect 5668 8134 5698 8186
rect 5698 8134 5710 8186
rect 5710 8134 5724 8186
rect 5748 8134 5762 8186
rect 5762 8134 5774 8186
rect 5774 8134 5804 8186
rect 5828 8134 5838 8186
rect 5838 8134 5884 8186
rect 5588 8132 5644 8134
rect 5668 8132 5724 8134
rect 5748 8132 5804 8134
rect 5828 8132 5884 8134
rect 5588 7098 5644 7100
rect 5668 7098 5724 7100
rect 5748 7098 5804 7100
rect 5828 7098 5884 7100
rect 5588 7046 5634 7098
rect 5634 7046 5644 7098
rect 5668 7046 5698 7098
rect 5698 7046 5710 7098
rect 5710 7046 5724 7098
rect 5748 7046 5762 7098
rect 5762 7046 5774 7098
rect 5774 7046 5804 7098
rect 5828 7046 5838 7098
rect 5838 7046 5884 7098
rect 5588 7044 5644 7046
rect 5668 7044 5724 7046
rect 5748 7044 5804 7046
rect 5828 7044 5884 7046
rect 5588 6010 5644 6012
rect 5668 6010 5724 6012
rect 5748 6010 5804 6012
rect 5828 6010 5884 6012
rect 5588 5958 5634 6010
rect 5634 5958 5644 6010
rect 5668 5958 5698 6010
rect 5698 5958 5710 6010
rect 5710 5958 5724 6010
rect 5748 5958 5762 6010
rect 5762 5958 5774 6010
rect 5774 5958 5804 6010
rect 5828 5958 5838 6010
rect 5838 5958 5884 6010
rect 5588 5956 5644 5958
rect 5668 5956 5724 5958
rect 5748 5956 5804 5958
rect 5828 5956 5884 5958
rect 5588 4922 5644 4924
rect 5668 4922 5724 4924
rect 5748 4922 5804 4924
rect 5828 4922 5884 4924
rect 5588 4870 5634 4922
rect 5634 4870 5644 4922
rect 5668 4870 5698 4922
rect 5698 4870 5710 4922
rect 5710 4870 5724 4922
rect 5748 4870 5762 4922
rect 5762 4870 5774 4922
rect 5774 4870 5804 4922
rect 5828 4870 5838 4922
rect 5838 4870 5884 4922
rect 5588 4868 5644 4870
rect 5668 4868 5724 4870
rect 5748 4868 5804 4870
rect 5828 4868 5884 4870
rect 5588 3834 5644 3836
rect 5668 3834 5724 3836
rect 5748 3834 5804 3836
rect 5828 3834 5884 3836
rect 5588 3782 5634 3834
rect 5634 3782 5644 3834
rect 5668 3782 5698 3834
rect 5698 3782 5710 3834
rect 5710 3782 5724 3834
rect 5748 3782 5762 3834
rect 5762 3782 5774 3834
rect 5774 3782 5804 3834
rect 5828 3782 5838 3834
rect 5838 3782 5884 3834
rect 5588 3780 5644 3782
rect 5668 3780 5724 3782
rect 5748 3780 5804 3782
rect 5828 3780 5884 3782
rect 5588 2746 5644 2748
rect 5668 2746 5724 2748
rect 5748 2746 5804 2748
rect 5828 2746 5884 2748
rect 5588 2694 5634 2746
rect 5634 2694 5644 2746
rect 5668 2694 5698 2746
rect 5698 2694 5710 2746
rect 5710 2694 5724 2746
rect 5748 2694 5762 2746
rect 5762 2694 5774 2746
rect 5774 2694 5804 2746
rect 5828 2694 5838 2746
rect 5838 2694 5884 2746
rect 5588 2692 5644 2694
rect 5668 2692 5724 2694
rect 5748 2692 5804 2694
rect 5828 2692 5884 2694
rect 10220 9818 10276 9820
rect 10300 9818 10356 9820
rect 10380 9818 10436 9820
rect 10460 9818 10516 9820
rect 10220 9766 10266 9818
rect 10266 9766 10276 9818
rect 10300 9766 10330 9818
rect 10330 9766 10342 9818
rect 10342 9766 10356 9818
rect 10380 9766 10394 9818
rect 10394 9766 10406 9818
rect 10406 9766 10436 9818
rect 10460 9766 10470 9818
rect 10470 9766 10516 9818
rect 10220 9764 10276 9766
rect 10300 9764 10356 9766
rect 10380 9764 10436 9766
rect 10460 9764 10516 9766
rect 12070 19796 12072 19816
rect 12072 19796 12124 19816
rect 12124 19796 12126 19816
rect 12070 19760 12126 19796
rect 11702 18284 11758 18320
rect 11702 18264 11704 18284
rect 11704 18264 11756 18284
rect 11756 18264 11758 18284
rect 11058 17196 11114 17232
rect 11058 17176 11060 17196
rect 11060 17176 11112 17196
rect 11112 17176 11114 17196
rect 11150 16360 11206 16416
rect 11150 13912 11206 13968
rect 11058 12280 11114 12336
rect 11426 16904 11482 16960
rect 11886 16360 11942 16416
rect 11702 15136 11758 15192
rect 12714 19796 12716 19816
rect 12716 19796 12768 19816
rect 12768 19796 12770 19816
rect 12714 19760 12770 19796
rect 12898 20984 12954 21040
rect 12254 13912 12310 13968
rect 11518 12044 11520 12064
rect 11520 12044 11572 12064
rect 11572 12044 11574 12064
rect 11518 12008 11574 12044
rect 10220 8730 10276 8732
rect 10300 8730 10356 8732
rect 10380 8730 10436 8732
rect 10460 8730 10516 8732
rect 10220 8678 10266 8730
rect 10266 8678 10276 8730
rect 10300 8678 10330 8730
rect 10330 8678 10342 8730
rect 10342 8678 10356 8730
rect 10380 8678 10394 8730
rect 10394 8678 10406 8730
rect 10406 8678 10436 8730
rect 10460 8678 10470 8730
rect 10470 8678 10516 8730
rect 10220 8676 10276 8678
rect 10300 8676 10356 8678
rect 10380 8676 10436 8678
rect 10460 8676 10516 8678
rect 10782 8336 10838 8392
rect 10220 7642 10276 7644
rect 10300 7642 10356 7644
rect 10380 7642 10436 7644
rect 10460 7642 10516 7644
rect 10220 7590 10266 7642
rect 10266 7590 10276 7642
rect 10300 7590 10330 7642
rect 10330 7590 10342 7642
rect 10342 7590 10356 7642
rect 10380 7590 10394 7642
rect 10394 7590 10406 7642
rect 10406 7590 10436 7642
rect 10460 7590 10470 7642
rect 10470 7590 10516 7642
rect 10220 7588 10276 7590
rect 10300 7588 10356 7590
rect 10380 7588 10436 7590
rect 10460 7588 10516 7590
rect 14852 26682 14908 26684
rect 14932 26682 14988 26684
rect 15012 26682 15068 26684
rect 15092 26682 15148 26684
rect 14852 26630 14898 26682
rect 14898 26630 14908 26682
rect 14932 26630 14962 26682
rect 14962 26630 14974 26682
rect 14974 26630 14988 26682
rect 15012 26630 15026 26682
rect 15026 26630 15038 26682
rect 15038 26630 15068 26682
rect 15092 26630 15102 26682
rect 15102 26630 15148 26682
rect 14852 26628 14908 26630
rect 14932 26628 14988 26630
rect 15012 26628 15068 26630
rect 15092 26628 15148 26630
rect 14852 25594 14908 25596
rect 14932 25594 14988 25596
rect 15012 25594 15068 25596
rect 15092 25594 15148 25596
rect 14852 25542 14898 25594
rect 14898 25542 14908 25594
rect 14932 25542 14962 25594
rect 14962 25542 14974 25594
rect 14974 25542 14988 25594
rect 15012 25542 15026 25594
rect 15026 25542 15038 25594
rect 15038 25542 15068 25594
rect 15092 25542 15102 25594
rect 15102 25542 15148 25594
rect 14852 25540 14908 25542
rect 14932 25540 14988 25542
rect 15012 25540 15068 25542
rect 15092 25540 15148 25542
rect 14852 24506 14908 24508
rect 14932 24506 14988 24508
rect 15012 24506 15068 24508
rect 15092 24506 15148 24508
rect 14852 24454 14898 24506
rect 14898 24454 14908 24506
rect 14932 24454 14962 24506
rect 14962 24454 14974 24506
rect 14974 24454 14988 24506
rect 15012 24454 15026 24506
rect 15026 24454 15038 24506
rect 15038 24454 15068 24506
rect 15092 24454 15102 24506
rect 15102 24454 15148 24506
rect 14852 24452 14908 24454
rect 14932 24452 14988 24454
rect 15012 24452 15068 24454
rect 15092 24452 15148 24454
rect 14852 23418 14908 23420
rect 14932 23418 14988 23420
rect 15012 23418 15068 23420
rect 15092 23418 15148 23420
rect 14852 23366 14898 23418
rect 14898 23366 14908 23418
rect 14932 23366 14962 23418
rect 14962 23366 14974 23418
rect 14974 23366 14988 23418
rect 15012 23366 15026 23418
rect 15026 23366 15038 23418
rect 15038 23366 15068 23418
rect 15092 23366 15102 23418
rect 15102 23366 15148 23418
rect 14852 23364 14908 23366
rect 14932 23364 14988 23366
rect 15012 23364 15068 23366
rect 15092 23364 15148 23366
rect 14852 22330 14908 22332
rect 14932 22330 14988 22332
rect 15012 22330 15068 22332
rect 15092 22330 15148 22332
rect 14852 22278 14898 22330
rect 14898 22278 14908 22330
rect 14932 22278 14962 22330
rect 14962 22278 14974 22330
rect 14974 22278 14988 22330
rect 15012 22278 15026 22330
rect 15026 22278 15038 22330
rect 15038 22278 15068 22330
rect 15092 22278 15102 22330
rect 15102 22278 15148 22330
rect 14852 22276 14908 22278
rect 14932 22276 14988 22278
rect 15012 22276 15068 22278
rect 15092 22276 15148 22278
rect 12990 16768 13046 16824
rect 12990 15408 13046 15464
rect 12898 15136 12954 15192
rect 13174 15272 13230 15328
rect 13450 15444 13452 15464
rect 13452 15444 13504 15464
rect 13504 15444 13506 15464
rect 13450 15408 13506 15444
rect 14186 20884 14188 20904
rect 14188 20884 14240 20904
rect 14240 20884 14242 20904
rect 14186 20848 14242 20884
rect 14852 21242 14908 21244
rect 14932 21242 14988 21244
rect 15012 21242 15068 21244
rect 15092 21242 15148 21244
rect 14852 21190 14898 21242
rect 14898 21190 14908 21242
rect 14932 21190 14962 21242
rect 14962 21190 14974 21242
rect 14974 21190 14988 21242
rect 15012 21190 15026 21242
rect 15026 21190 15038 21242
rect 15038 21190 15068 21242
rect 15092 21190 15102 21242
rect 15102 21190 15148 21242
rect 14852 21188 14908 21190
rect 14932 21188 14988 21190
rect 15012 21188 15068 21190
rect 15092 21188 15148 21190
rect 14738 20984 14794 21040
rect 14852 20154 14908 20156
rect 14932 20154 14988 20156
rect 15012 20154 15068 20156
rect 15092 20154 15148 20156
rect 14852 20102 14898 20154
rect 14898 20102 14908 20154
rect 14932 20102 14962 20154
rect 14962 20102 14974 20154
rect 14974 20102 14988 20154
rect 15012 20102 15026 20154
rect 15026 20102 15038 20154
rect 15038 20102 15068 20154
rect 15092 20102 15102 20154
rect 15102 20102 15148 20154
rect 14852 20100 14908 20102
rect 14932 20100 14988 20102
rect 15012 20100 15068 20102
rect 15092 20100 15148 20102
rect 13082 14884 13138 14920
rect 13082 14864 13084 14884
rect 13084 14864 13136 14884
rect 13136 14864 13138 14884
rect 12714 12044 12716 12064
rect 12716 12044 12768 12064
rect 12768 12044 12770 12064
rect 12714 12008 12770 12044
rect 12714 9596 12716 9616
rect 12716 9596 12768 9616
rect 12768 9596 12770 9616
rect 12714 9560 12770 9596
rect 10220 6554 10276 6556
rect 10300 6554 10356 6556
rect 10380 6554 10436 6556
rect 10460 6554 10516 6556
rect 10220 6502 10266 6554
rect 10266 6502 10276 6554
rect 10300 6502 10330 6554
rect 10330 6502 10342 6554
rect 10342 6502 10356 6554
rect 10380 6502 10394 6554
rect 10394 6502 10406 6554
rect 10406 6502 10436 6554
rect 10460 6502 10470 6554
rect 10470 6502 10516 6554
rect 10220 6500 10276 6502
rect 10300 6500 10356 6502
rect 10380 6500 10436 6502
rect 10460 6500 10516 6502
rect 10220 5466 10276 5468
rect 10300 5466 10356 5468
rect 10380 5466 10436 5468
rect 10460 5466 10516 5468
rect 10220 5414 10266 5466
rect 10266 5414 10276 5466
rect 10300 5414 10330 5466
rect 10330 5414 10342 5466
rect 10342 5414 10356 5466
rect 10380 5414 10394 5466
rect 10394 5414 10406 5466
rect 10406 5414 10436 5466
rect 10460 5414 10470 5466
rect 10470 5414 10516 5466
rect 10220 5412 10276 5414
rect 10300 5412 10356 5414
rect 10380 5412 10436 5414
rect 10460 5412 10516 5414
rect 10220 4378 10276 4380
rect 10300 4378 10356 4380
rect 10380 4378 10436 4380
rect 10460 4378 10516 4380
rect 10220 4326 10266 4378
rect 10266 4326 10276 4378
rect 10300 4326 10330 4378
rect 10330 4326 10342 4378
rect 10342 4326 10356 4378
rect 10380 4326 10394 4378
rect 10394 4326 10406 4378
rect 10406 4326 10436 4378
rect 10460 4326 10470 4378
rect 10470 4326 10516 4378
rect 10220 4324 10276 4326
rect 10300 4324 10356 4326
rect 10380 4324 10436 4326
rect 10460 4324 10516 4326
rect 10220 3290 10276 3292
rect 10300 3290 10356 3292
rect 10380 3290 10436 3292
rect 10460 3290 10516 3292
rect 10220 3238 10266 3290
rect 10266 3238 10276 3290
rect 10300 3238 10330 3290
rect 10330 3238 10342 3290
rect 10342 3238 10356 3290
rect 10380 3238 10394 3290
rect 10394 3238 10406 3290
rect 10406 3238 10436 3290
rect 10460 3238 10470 3290
rect 10470 3238 10516 3290
rect 10220 3236 10276 3238
rect 10300 3236 10356 3238
rect 10380 3236 10436 3238
rect 10460 3236 10516 3238
rect 13818 14492 13820 14512
rect 13820 14492 13872 14512
rect 13872 14492 13874 14512
rect 13818 14456 13874 14492
rect 14852 19066 14908 19068
rect 14932 19066 14988 19068
rect 15012 19066 15068 19068
rect 15092 19066 15148 19068
rect 14852 19014 14898 19066
rect 14898 19014 14908 19066
rect 14932 19014 14962 19066
rect 14962 19014 14974 19066
rect 14974 19014 14988 19066
rect 15012 19014 15026 19066
rect 15026 19014 15038 19066
rect 15038 19014 15068 19066
rect 15092 19014 15102 19066
rect 15102 19014 15148 19066
rect 14852 19012 14908 19014
rect 14932 19012 14988 19014
rect 15012 19012 15068 19014
rect 15092 19012 15148 19014
rect 19484 27226 19540 27228
rect 19564 27226 19620 27228
rect 19644 27226 19700 27228
rect 19724 27226 19780 27228
rect 19484 27174 19530 27226
rect 19530 27174 19540 27226
rect 19564 27174 19594 27226
rect 19594 27174 19606 27226
rect 19606 27174 19620 27226
rect 19644 27174 19658 27226
rect 19658 27174 19670 27226
rect 19670 27174 19700 27226
rect 19724 27174 19734 27226
rect 19734 27174 19780 27226
rect 19484 27172 19540 27174
rect 19564 27172 19620 27174
rect 19644 27172 19700 27174
rect 19724 27172 19780 27174
rect 16302 24928 16358 24984
rect 15750 24112 15806 24168
rect 17314 25336 17370 25392
rect 14646 16904 14702 16960
rect 14094 14864 14150 14920
rect 14370 15020 14426 15056
rect 14370 15000 14372 15020
rect 14372 15000 14424 15020
rect 14424 15000 14426 15020
rect 14462 14476 14518 14512
rect 14462 14456 14464 14476
rect 14464 14456 14516 14476
rect 14516 14456 14518 14476
rect 14852 17978 14908 17980
rect 14932 17978 14988 17980
rect 15012 17978 15068 17980
rect 15092 17978 15148 17980
rect 14852 17926 14898 17978
rect 14898 17926 14908 17978
rect 14932 17926 14962 17978
rect 14962 17926 14974 17978
rect 14974 17926 14988 17978
rect 15012 17926 15026 17978
rect 15026 17926 15038 17978
rect 15038 17926 15068 17978
rect 15092 17926 15102 17978
rect 15102 17926 15148 17978
rect 14852 17924 14908 17926
rect 14932 17924 14988 17926
rect 15012 17924 15068 17926
rect 15092 17924 15148 17926
rect 14852 16890 14908 16892
rect 14932 16890 14988 16892
rect 15012 16890 15068 16892
rect 15092 16890 15148 16892
rect 14852 16838 14898 16890
rect 14898 16838 14908 16890
rect 14932 16838 14962 16890
rect 14962 16838 14974 16890
rect 14974 16838 14988 16890
rect 15012 16838 15026 16890
rect 15026 16838 15038 16890
rect 15038 16838 15068 16890
rect 15092 16838 15102 16890
rect 15102 16838 15148 16890
rect 14852 16836 14908 16838
rect 14932 16836 14988 16838
rect 15012 16836 15068 16838
rect 15092 16836 15148 16838
rect 15842 19780 15898 19816
rect 15842 19760 15844 19780
rect 15844 19760 15896 19780
rect 15896 19760 15898 19780
rect 15566 17740 15622 17776
rect 15566 17720 15568 17740
rect 15568 17720 15620 17740
rect 15620 17720 15622 17740
rect 14852 15802 14908 15804
rect 14932 15802 14988 15804
rect 15012 15802 15068 15804
rect 15092 15802 15148 15804
rect 14852 15750 14898 15802
rect 14898 15750 14908 15802
rect 14932 15750 14962 15802
rect 14962 15750 14974 15802
rect 14974 15750 14988 15802
rect 15012 15750 15026 15802
rect 15026 15750 15038 15802
rect 15038 15750 15068 15802
rect 15092 15750 15102 15802
rect 15102 15750 15148 15802
rect 14852 15748 14908 15750
rect 14932 15748 14988 15750
rect 15012 15748 15068 15750
rect 15092 15748 15148 15750
rect 14738 15000 14794 15056
rect 14646 13776 14702 13832
rect 14852 14714 14908 14716
rect 14932 14714 14988 14716
rect 15012 14714 15068 14716
rect 15092 14714 15148 14716
rect 14852 14662 14898 14714
rect 14898 14662 14908 14714
rect 14932 14662 14962 14714
rect 14962 14662 14974 14714
rect 14974 14662 14988 14714
rect 15012 14662 15026 14714
rect 15026 14662 15038 14714
rect 15038 14662 15068 14714
rect 15092 14662 15102 14714
rect 15102 14662 15148 14714
rect 14852 14660 14908 14662
rect 14932 14660 14988 14662
rect 15012 14660 15068 14662
rect 15092 14660 15148 14662
rect 15290 14320 15346 14376
rect 14852 13626 14908 13628
rect 14932 13626 14988 13628
rect 15012 13626 15068 13628
rect 15092 13626 15148 13628
rect 14852 13574 14898 13626
rect 14898 13574 14908 13626
rect 14932 13574 14962 13626
rect 14962 13574 14974 13626
rect 14974 13574 14988 13626
rect 15012 13574 15026 13626
rect 15026 13574 15038 13626
rect 15038 13574 15068 13626
rect 15092 13574 15102 13626
rect 15102 13574 15148 13626
rect 14852 13572 14908 13574
rect 14932 13572 14988 13574
rect 15012 13572 15068 13574
rect 15092 13572 15148 13574
rect 14852 12538 14908 12540
rect 14932 12538 14988 12540
rect 15012 12538 15068 12540
rect 15092 12538 15148 12540
rect 14852 12486 14898 12538
rect 14898 12486 14908 12538
rect 14932 12486 14962 12538
rect 14962 12486 14974 12538
rect 14974 12486 14988 12538
rect 15012 12486 15026 12538
rect 15026 12486 15038 12538
rect 15038 12486 15068 12538
rect 15092 12486 15102 12538
rect 15102 12486 15148 12538
rect 14852 12484 14908 12486
rect 14932 12484 14988 12486
rect 15012 12484 15068 12486
rect 15092 12484 15148 12486
rect 14278 12280 14334 12336
rect 13634 8628 13690 8664
rect 13634 8608 13636 8628
rect 13636 8608 13688 8628
rect 13688 8608 13690 8628
rect 14852 11450 14908 11452
rect 14932 11450 14988 11452
rect 15012 11450 15068 11452
rect 15092 11450 15148 11452
rect 14852 11398 14898 11450
rect 14898 11398 14908 11450
rect 14932 11398 14962 11450
rect 14962 11398 14974 11450
rect 14974 11398 14988 11450
rect 15012 11398 15026 11450
rect 15026 11398 15038 11450
rect 15038 11398 15068 11450
rect 15092 11398 15102 11450
rect 15102 11398 15148 11450
rect 14852 11396 14908 11398
rect 14932 11396 14988 11398
rect 15012 11396 15068 11398
rect 15092 11396 15148 11398
rect 14852 10362 14908 10364
rect 14932 10362 14988 10364
rect 15012 10362 15068 10364
rect 15092 10362 15148 10364
rect 14852 10310 14898 10362
rect 14898 10310 14908 10362
rect 14932 10310 14962 10362
rect 14962 10310 14974 10362
rect 14974 10310 14988 10362
rect 15012 10310 15026 10362
rect 15026 10310 15038 10362
rect 15038 10310 15068 10362
rect 15092 10310 15102 10362
rect 15102 10310 15148 10362
rect 14852 10308 14908 10310
rect 14932 10308 14988 10310
rect 15012 10308 15068 10310
rect 15092 10308 15148 10310
rect 14852 9274 14908 9276
rect 14932 9274 14988 9276
rect 15012 9274 15068 9276
rect 15092 9274 15148 9276
rect 14852 9222 14898 9274
rect 14898 9222 14908 9274
rect 14932 9222 14962 9274
rect 14962 9222 14974 9274
rect 14974 9222 14988 9274
rect 15012 9222 15026 9274
rect 15026 9222 15038 9274
rect 15038 9222 15068 9274
rect 15092 9222 15102 9274
rect 15102 9222 15148 9274
rect 14852 9220 14908 9222
rect 14932 9220 14988 9222
rect 15012 9220 15068 9222
rect 15092 9220 15148 9222
rect 15566 9596 15568 9616
rect 15568 9596 15620 9616
rect 15620 9596 15622 9616
rect 15566 9560 15622 9596
rect 16118 12144 16174 12200
rect 16854 18420 16910 18456
rect 16854 18400 16856 18420
rect 16856 18400 16908 18420
rect 16908 18400 16910 18420
rect 17590 18284 17646 18320
rect 17590 18264 17592 18284
rect 17592 18264 17644 18284
rect 17644 18264 17646 18284
rect 18418 19896 18474 19952
rect 19484 26138 19540 26140
rect 19564 26138 19620 26140
rect 19644 26138 19700 26140
rect 19724 26138 19780 26140
rect 19484 26086 19530 26138
rect 19530 26086 19540 26138
rect 19564 26086 19594 26138
rect 19594 26086 19606 26138
rect 19606 26086 19620 26138
rect 19644 26086 19658 26138
rect 19658 26086 19670 26138
rect 19670 26086 19700 26138
rect 19724 26086 19734 26138
rect 19734 26086 19780 26138
rect 19484 26084 19540 26086
rect 19564 26084 19620 26086
rect 19644 26084 19700 26086
rect 19724 26084 19780 26086
rect 19484 25050 19540 25052
rect 19564 25050 19620 25052
rect 19644 25050 19700 25052
rect 19724 25050 19780 25052
rect 19484 24998 19530 25050
rect 19530 24998 19540 25050
rect 19564 24998 19594 25050
rect 19594 24998 19606 25050
rect 19606 24998 19620 25050
rect 19644 24998 19658 25050
rect 19658 24998 19670 25050
rect 19670 24998 19700 25050
rect 19724 24998 19734 25050
rect 19734 24998 19780 25050
rect 19484 24996 19540 24998
rect 19564 24996 19620 24998
rect 19644 24996 19700 24998
rect 19724 24996 19780 24998
rect 19484 23962 19540 23964
rect 19564 23962 19620 23964
rect 19644 23962 19700 23964
rect 19724 23962 19780 23964
rect 19484 23910 19530 23962
rect 19530 23910 19540 23962
rect 19564 23910 19594 23962
rect 19594 23910 19606 23962
rect 19606 23910 19620 23962
rect 19644 23910 19658 23962
rect 19658 23910 19670 23962
rect 19670 23910 19700 23962
rect 19724 23910 19734 23962
rect 19734 23910 19780 23962
rect 19484 23908 19540 23910
rect 19564 23908 19620 23910
rect 19644 23908 19700 23910
rect 19724 23908 19780 23910
rect 24116 27770 24172 27772
rect 24196 27770 24252 27772
rect 24276 27770 24332 27772
rect 24356 27770 24412 27772
rect 24116 27718 24162 27770
rect 24162 27718 24172 27770
rect 24196 27718 24226 27770
rect 24226 27718 24238 27770
rect 24238 27718 24252 27770
rect 24276 27718 24290 27770
rect 24290 27718 24302 27770
rect 24302 27718 24332 27770
rect 24356 27718 24366 27770
rect 24366 27718 24412 27770
rect 24116 27716 24172 27718
rect 24196 27716 24252 27718
rect 24276 27716 24332 27718
rect 24356 27716 24412 27718
rect 27526 28600 27582 28656
rect 21086 25336 21142 25392
rect 20718 24112 20774 24168
rect 19484 22874 19540 22876
rect 19564 22874 19620 22876
rect 19644 22874 19700 22876
rect 19724 22874 19780 22876
rect 19484 22822 19530 22874
rect 19530 22822 19540 22874
rect 19564 22822 19594 22874
rect 19594 22822 19606 22874
rect 19606 22822 19620 22874
rect 19644 22822 19658 22874
rect 19658 22822 19670 22874
rect 19670 22822 19700 22874
rect 19724 22822 19734 22874
rect 19734 22822 19780 22874
rect 19484 22820 19540 22822
rect 19564 22820 19620 22822
rect 19644 22820 19700 22822
rect 19724 22820 19780 22822
rect 19484 21786 19540 21788
rect 19564 21786 19620 21788
rect 19644 21786 19700 21788
rect 19724 21786 19780 21788
rect 19484 21734 19530 21786
rect 19530 21734 19540 21786
rect 19564 21734 19594 21786
rect 19594 21734 19606 21786
rect 19606 21734 19620 21786
rect 19644 21734 19658 21786
rect 19658 21734 19670 21786
rect 19670 21734 19700 21786
rect 19724 21734 19734 21786
rect 19734 21734 19780 21786
rect 19484 21732 19540 21734
rect 19564 21732 19620 21734
rect 19644 21732 19700 21734
rect 19724 21732 19780 21734
rect 18878 20440 18934 20496
rect 18878 19896 18934 19952
rect 17130 16632 17186 16688
rect 17130 16108 17186 16144
rect 17130 16088 17132 16108
rect 17132 16088 17184 16108
rect 17184 16088 17186 16108
rect 17958 17196 18014 17232
rect 17958 17176 17960 17196
rect 17960 17176 18012 17196
rect 18012 17176 18014 17196
rect 17958 16360 18014 16416
rect 16302 11736 16358 11792
rect 16210 11228 16212 11248
rect 16212 11228 16264 11248
rect 16264 11228 16266 11248
rect 16210 11192 16266 11228
rect 15382 8336 15438 8392
rect 14852 8186 14908 8188
rect 14932 8186 14988 8188
rect 15012 8186 15068 8188
rect 15092 8186 15148 8188
rect 14852 8134 14898 8186
rect 14898 8134 14908 8186
rect 14932 8134 14962 8186
rect 14962 8134 14974 8186
rect 14974 8134 14988 8186
rect 15012 8134 15026 8186
rect 15026 8134 15038 8186
rect 15038 8134 15068 8186
rect 15092 8134 15102 8186
rect 15102 8134 15148 8186
rect 14852 8132 14908 8134
rect 14932 8132 14988 8134
rect 15012 8132 15068 8134
rect 15092 8132 15148 8134
rect 13450 6840 13506 6896
rect 14852 7098 14908 7100
rect 14932 7098 14988 7100
rect 15012 7098 15068 7100
rect 15092 7098 15148 7100
rect 14852 7046 14898 7098
rect 14898 7046 14908 7098
rect 14932 7046 14962 7098
rect 14962 7046 14974 7098
rect 14974 7046 14988 7098
rect 15012 7046 15026 7098
rect 15026 7046 15038 7098
rect 15038 7046 15068 7098
rect 15092 7046 15102 7098
rect 15102 7046 15148 7098
rect 14852 7044 14908 7046
rect 14932 7044 14988 7046
rect 15012 7044 15068 7046
rect 15092 7044 15148 7046
rect 14852 6010 14908 6012
rect 14932 6010 14988 6012
rect 15012 6010 15068 6012
rect 15092 6010 15148 6012
rect 14852 5958 14898 6010
rect 14898 5958 14908 6010
rect 14932 5958 14962 6010
rect 14962 5958 14974 6010
rect 14974 5958 14988 6010
rect 15012 5958 15026 6010
rect 15026 5958 15038 6010
rect 15038 5958 15068 6010
rect 15092 5958 15102 6010
rect 15102 5958 15148 6010
rect 14852 5956 14908 5958
rect 14932 5956 14988 5958
rect 15012 5956 15068 5958
rect 15092 5956 15148 5958
rect 14852 4922 14908 4924
rect 14932 4922 14988 4924
rect 15012 4922 15068 4924
rect 15092 4922 15148 4924
rect 14852 4870 14898 4922
rect 14898 4870 14908 4922
rect 14932 4870 14962 4922
rect 14962 4870 14974 4922
rect 14974 4870 14988 4922
rect 15012 4870 15026 4922
rect 15026 4870 15038 4922
rect 15038 4870 15068 4922
rect 15092 4870 15102 4922
rect 15102 4870 15148 4922
rect 14852 4868 14908 4870
rect 14932 4868 14988 4870
rect 15012 4868 15068 4870
rect 15092 4868 15148 4870
rect 14852 3834 14908 3836
rect 14932 3834 14988 3836
rect 15012 3834 15068 3836
rect 15092 3834 15148 3836
rect 14852 3782 14898 3834
rect 14898 3782 14908 3834
rect 14932 3782 14962 3834
rect 14962 3782 14974 3834
rect 14974 3782 14988 3834
rect 15012 3782 15026 3834
rect 15026 3782 15038 3834
rect 15038 3782 15068 3834
rect 15092 3782 15102 3834
rect 15102 3782 15148 3834
rect 14852 3780 14908 3782
rect 14932 3780 14988 3782
rect 15012 3780 15068 3782
rect 15092 3780 15148 3782
rect 14852 2746 14908 2748
rect 14932 2746 14988 2748
rect 15012 2746 15068 2748
rect 15092 2746 15148 2748
rect 1490 1400 1546 1456
rect 14852 2694 14898 2746
rect 14898 2694 14908 2746
rect 14932 2694 14962 2746
rect 14962 2694 14974 2746
rect 14974 2694 14988 2746
rect 15012 2694 15026 2746
rect 15026 2694 15038 2746
rect 15038 2694 15068 2746
rect 15092 2694 15102 2746
rect 15102 2694 15148 2746
rect 14852 2692 14908 2694
rect 14932 2692 14988 2694
rect 15012 2692 15068 2694
rect 15092 2692 15148 2694
rect 17130 11636 17132 11656
rect 17132 11636 17184 11656
rect 17184 11636 17186 11656
rect 17130 11600 17186 11636
rect 17958 15428 18014 15464
rect 17958 15408 17960 15428
rect 17960 15408 18012 15428
rect 18012 15408 18014 15428
rect 17682 13912 17738 13968
rect 18602 17584 18658 17640
rect 18602 16360 18658 16416
rect 18878 16088 18934 16144
rect 16670 8608 16726 8664
rect 18694 14356 18696 14376
rect 18696 14356 18748 14376
rect 18748 14356 18750 14376
rect 18694 14320 18750 14356
rect 18142 8880 18198 8936
rect 19484 20698 19540 20700
rect 19564 20698 19620 20700
rect 19644 20698 19700 20700
rect 19724 20698 19780 20700
rect 19484 20646 19530 20698
rect 19530 20646 19540 20698
rect 19564 20646 19594 20698
rect 19594 20646 19606 20698
rect 19606 20646 19620 20698
rect 19644 20646 19658 20698
rect 19658 20646 19670 20698
rect 19670 20646 19700 20698
rect 19724 20646 19734 20698
rect 19734 20646 19780 20698
rect 19484 20644 19540 20646
rect 19564 20644 19620 20646
rect 19644 20644 19700 20646
rect 19724 20644 19780 20646
rect 19484 19610 19540 19612
rect 19564 19610 19620 19612
rect 19644 19610 19700 19612
rect 19724 19610 19780 19612
rect 19484 19558 19530 19610
rect 19530 19558 19540 19610
rect 19564 19558 19594 19610
rect 19594 19558 19606 19610
rect 19606 19558 19620 19610
rect 19644 19558 19658 19610
rect 19658 19558 19670 19610
rect 19670 19558 19700 19610
rect 19724 19558 19734 19610
rect 19734 19558 19780 19610
rect 19484 19556 19540 19558
rect 19564 19556 19620 19558
rect 19644 19556 19700 19558
rect 19724 19556 19780 19558
rect 19484 18522 19540 18524
rect 19564 18522 19620 18524
rect 19644 18522 19700 18524
rect 19724 18522 19780 18524
rect 19484 18470 19530 18522
rect 19530 18470 19540 18522
rect 19564 18470 19594 18522
rect 19594 18470 19606 18522
rect 19606 18470 19620 18522
rect 19644 18470 19658 18522
rect 19658 18470 19670 18522
rect 19670 18470 19700 18522
rect 19724 18470 19734 18522
rect 19734 18470 19780 18522
rect 19484 18468 19540 18470
rect 19564 18468 19620 18470
rect 19644 18468 19700 18470
rect 19724 18468 19780 18470
rect 19982 18400 20038 18456
rect 19484 17434 19540 17436
rect 19564 17434 19620 17436
rect 19644 17434 19700 17436
rect 19724 17434 19780 17436
rect 19484 17382 19530 17434
rect 19530 17382 19540 17434
rect 19564 17382 19594 17434
rect 19594 17382 19606 17434
rect 19606 17382 19620 17434
rect 19644 17382 19658 17434
rect 19658 17382 19670 17434
rect 19670 17382 19700 17434
rect 19724 17382 19734 17434
rect 19734 17382 19780 17434
rect 19484 17380 19540 17382
rect 19564 17380 19620 17382
rect 19644 17380 19700 17382
rect 19724 17380 19780 17382
rect 19484 16346 19540 16348
rect 19564 16346 19620 16348
rect 19644 16346 19700 16348
rect 19724 16346 19780 16348
rect 19484 16294 19530 16346
rect 19530 16294 19540 16346
rect 19564 16294 19594 16346
rect 19594 16294 19606 16346
rect 19606 16294 19620 16346
rect 19644 16294 19658 16346
rect 19658 16294 19670 16346
rect 19670 16294 19700 16346
rect 19724 16294 19734 16346
rect 19734 16294 19780 16346
rect 19484 16292 19540 16294
rect 19564 16292 19620 16294
rect 19644 16292 19700 16294
rect 19724 16292 19780 16294
rect 19484 15258 19540 15260
rect 19564 15258 19620 15260
rect 19644 15258 19700 15260
rect 19724 15258 19780 15260
rect 19484 15206 19530 15258
rect 19530 15206 19540 15258
rect 19564 15206 19594 15258
rect 19594 15206 19606 15258
rect 19606 15206 19620 15258
rect 19644 15206 19658 15258
rect 19658 15206 19670 15258
rect 19670 15206 19700 15258
rect 19724 15206 19734 15258
rect 19734 15206 19780 15258
rect 19484 15204 19540 15206
rect 19564 15204 19620 15206
rect 19644 15204 19700 15206
rect 19724 15204 19780 15206
rect 19484 14170 19540 14172
rect 19564 14170 19620 14172
rect 19644 14170 19700 14172
rect 19724 14170 19780 14172
rect 19484 14118 19530 14170
rect 19530 14118 19540 14170
rect 19564 14118 19594 14170
rect 19594 14118 19606 14170
rect 19606 14118 19620 14170
rect 19644 14118 19658 14170
rect 19658 14118 19670 14170
rect 19670 14118 19700 14170
rect 19724 14118 19734 14170
rect 19734 14118 19780 14170
rect 19484 14116 19540 14118
rect 19564 14116 19620 14118
rect 19644 14116 19700 14118
rect 19724 14116 19780 14118
rect 19798 13232 19854 13288
rect 19484 13082 19540 13084
rect 19564 13082 19620 13084
rect 19644 13082 19700 13084
rect 19724 13082 19780 13084
rect 19484 13030 19530 13082
rect 19530 13030 19540 13082
rect 19564 13030 19594 13082
rect 19594 13030 19606 13082
rect 19606 13030 19620 13082
rect 19644 13030 19658 13082
rect 19658 13030 19670 13082
rect 19670 13030 19700 13082
rect 19724 13030 19734 13082
rect 19734 13030 19780 13082
rect 19484 13028 19540 13030
rect 19564 13028 19620 13030
rect 19644 13028 19700 13030
rect 19724 13028 19780 13030
rect 19484 11994 19540 11996
rect 19564 11994 19620 11996
rect 19644 11994 19700 11996
rect 19724 11994 19780 11996
rect 19484 11942 19530 11994
rect 19530 11942 19540 11994
rect 19564 11942 19594 11994
rect 19594 11942 19606 11994
rect 19606 11942 19620 11994
rect 19644 11942 19658 11994
rect 19658 11942 19670 11994
rect 19670 11942 19700 11994
rect 19724 11942 19734 11994
rect 19734 11942 19780 11994
rect 19484 11940 19540 11942
rect 19564 11940 19620 11942
rect 19644 11940 19700 11942
rect 19724 11940 19780 11942
rect 19798 11756 19854 11792
rect 19798 11736 19800 11756
rect 19800 11736 19852 11756
rect 19852 11736 19854 11756
rect 19484 10906 19540 10908
rect 19564 10906 19620 10908
rect 19644 10906 19700 10908
rect 19724 10906 19780 10908
rect 19484 10854 19530 10906
rect 19530 10854 19540 10906
rect 19564 10854 19594 10906
rect 19594 10854 19606 10906
rect 19606 10854 19620 10906
rect 19644 10854 19658 10906
rect 19658 10854 19670 10906
rect 19670 10854 19700 10906
rect 19724 10854 19734 10906
rect 19734 10854 19780 10906
rect 19484 10852 19540 10854
rect 19564 10852 19620 10854
rect 19644 10852 19700 10854
rect 19724 10852 19780 10854
rect 24116 26682 24172 26684
rect 24196 26682 24252 26684
rect 24276 26682 24332 26684
rect 24356 26682 24412 26684
rect 24116 26630 24162 26682
rect 24162 26630 24172 26682
rect 24196 26630 24226 26682
rect 24226 26630 24238 26682
rect 24238 26630 24252 26682
rect 24276 26630 24290 26682
rect 24290 26630 24302 26682
rect 24302 26630 24332 26682
rect 24356 26630 24366 26682
rect 24366 26630 24412 26682
rect 24116 26628 24172 26630
rect 24196 26628 24252 26630
rect 24276 26628 24332 26630
rect 24356 26628 24412 26630
rect 24116 25594 24172 25596
rect 24196 25594 24252 25596
rect 24276 25594 24332 25596
rect 24356 25594 24412 25596
rect 24116 25542 24162 25594
rect 24162 25542 24172 25594
rect 24196 25542 24226 25594
rect 24226 25542 24238 25594
rect 24238 25542 24252 25594
rect 24276 25542 24290 25594
rect 24290 25542 24302 25594
rect 24302 25542 24332 25594
rect 24356 25542 24366 25594
rect 24366 25542 24412 25594
rect 24116 25540 24172 25542
rect 24196 25540 24252 25542
rect 24276 25540 24332 25542
rect 24356 25540 24412 25542
rect 24116 24506 24172 24508
rect 24196 24506 24252 24508
rect 24276 24506 24332 24508
rect 24356 24506 24412 24508
rect 24116 24454 24162 24506
rect 24162 24454 24172 24506
rect 24196 24454 24226 24506
rect 24226 24454 24238 24506
rect 24238 24454 24252 24506
rect 24276 24454 24290 24506
rect 24290 24454 24302 24506
rect 24302 24454 24332 24506
rect 24356 24454 24366 24506
rect 24366 24454 24412 24506
rect 24116 24452 24172 24454
rect 24196 24452 24252 24454
rect 24276 24452 24332 24454
rect 24356 24452 24412 24454
rect 24116 23418 24172 23420
rect 24196 23418 24252 23420
rect 24276 23418 24332 23420
rect 24356 23418 24412 23420
rect 24116 23366 24162 23418
rect 24162 23366 24172 23418
rect 24196 23366 24226 23418
rect 24226 23366 24238 23418
rect 24238 23366 24252 23418
rect 24276 23366 24290 23418
rect 24290 23366 24302 23418
rect 24302 23366 24332 23418
rect 24356 23366 24366 23418
rect 24366 23366 24412 23418
rect 24116 23364 24172 23366
rect 24196 23364 24252 23366
rect 24276 23364 24332 23366
rect 24356 23364 24412 23366
rect 22926 21392 22982 21448
rect 21454 19624 21510 19680
rect 20994 14356 20996 14376
rect 20996 14356 21048 14376
rect 21048 14356 21050 14376
rect 20994 14320 21050 14356
rect 20902 14048 20958 14104
rect 21362 14048 21418 14104
rect 20534 12960 20590 13016
rect 19982 10104 20038 10160
rect 19484 9818 19540 9820
rect 19564 9818 19620 9820
rect 19644 9818 19700 9820
rect 19724 9818 19780 9820
rect 19484 9766 19530 9818
rect 19530 9766 19540 9818
rect 19564 9766 19594 9818
rect 19594 9766 19606 9818
rect 19606 9766 19620 9818
rect 19644 9766 19658 9818
rect 19658 9766 19670 9818
rect 19670 9766 19700 9818
rect 19724 9766 19734 9818
rect 19734 9766 19780 9818
rect 19484 9764 19540 9766
rect 19564 9764 19620 9766
rect 19644 9764 19700 9766
rect 19724 9764 19780 9766
rect 22282 19624 22338 19680
rect 22190 19216 22246 19272
rect 23294 18400 23350 18456
rect 21454 13368 21510 13424
rect 20626 12708 20682 12744
rect 20626 12688 20628 12708
rect 20628 12688 20680 12708
rect 20680 12688 20682 12708
rect 22558 12980 22614 13016
rect 22558 12960 22560 12980
rect 22560 12960 22612 12980
rect 22612 12960 22614 12980
rect 22098 12416 22154 12472
rect 22282 11600 22338 11656
rect 19484 8730 19540 8732
rect 19564 8730 19620 8732
rect 19644 8730 19700 8732
rect 19724 8730 19780 8732
rect 19484 8678 19530 8730
rect 19530 8678 19540 8730
rect 19564 8678 19594 8730
rect 19594 8678 19606 8730
rect 19606 8678 19620 8730
rect 19644 8678 19658 8730
rect 19658 8678 19670 8730
rect 19670 8678 19700 8730
rect 19724 8678 19734 8730
rect 19734 8678 19780 8730
rect 19484 8676 19540 8678
rect 19564 8676 19620 8678
rect 19644 8676 19700 8678
rect 19724 8676 19780 8678
rect 19484 7642 19540 7644
rect 19564 7642 19620 7644
rect 19644 7642 19700 7644
rect 19724 7642 19780 7644
rect 19484 7590 19530 7642
rect 19530 7590 19540 7642
rect 19564 7590 19594 7642
rect 19594 7590 19606 7642
rect 19606 7590 19620 7642
rect 19644 7590 19658 7642
rect 19658 7590 19670 7642
rect 19670 7590 19700 7642
rect 19724 7590 19734 7642
rect 19734 7590 19780 7642
rect 19484 7588 19540 7590
rect 19564 7588 19620 7590
rect 19644 7588 19700 7590
rect 19724 7588 19780 7590
rect 19484 6554 19540 6556
rect 19564 6554 19620 6556
rect 19644 6554 19700 6556
rect 19724 6554 19780 6556
rect 19484 6502 19530 6554
rect 19530 6502 19540 6554
rect 19564 6502 19594 6554
rect 19594 6502 19606 6554
rect 19606 6502 19620 6554
rect 19644 6502 19658 6554
rect 19658 6502 19670 6554
rect 19670 6502 19700 6554
rect 19724 6502 19734 6554
rect 19734 6502 19780 6554
rect 19484 6500 19540 6502
rect 19564 6500 19620 6502
rect 19644 6500 19700 6502
rect 19724 6500 19780 6502
rect 24116 22330 24172 22332
rect 24196 22330 24252 22332
rect 24276 22330 24332 22332
rect 24356 22330 24412 22332
rect 24116 22278 24162 22330
rect 24162 22278 24172 22330
rect 24196 22278 24226 22330
rect 24226 22278 24238 22330
rect 24238 22278 24252 22330
rect 24276 22278 24290 22330
rect 24290 22278 24302 22330
rect 24302 22278 24332 22330
rect 24356 22278 24366 22330
rect 24366 22278 24412 22330
rect 24116 22276 24172 22278
rect 24196 22276 24252 22278
rect 24276 22276 24332 22278
rect 24356 22276 24412 22278
rect 24306 22092 24362 22128
rect 24306 22072 24308 22092
rect 24308 22072 24360 22092
rect 24360 22072 24362 22092
rect 24306 21956 24362 21992
rect 24306 21936 24308 21956
rect 24308 21936 24360 21956
rect 24360 21936 24362 21956
rect 24116 21242 24172 21244
rect 24196 21242 24252 21244
rect 24276 21242 24332 21244
rect 24356 21242 24412 21244
rect 24116 21190 24162 21242
rect 24162 21190 24172 21242
rect 24196 21190 24226 21242
rect 24226 21190 24238 21242
rect 24238 21190 24252 21242
rect 24276 21190 24290 21242
rect 24290 21190 24302 21242
rect 24302 21190 24332 21242
rect 24356 21190 24366 21242
rect 24366 21190 24412 21242
rect 24116 21188 24172 21190
rect 24196 21188 24252 21190
rect 24276 21188 24332 21190
rect 24356 21188 24412 21190
rect 25134 26308 25190 26344
rect 25134 26288 25136 26308
rect 25136 26288 25188 26308
rect 25188 26288 25190 26308
rect 25502 26288 25558 26344
rect 25042 21936 25098 21992
rect 24116 20154 24172 20156
rect 24196 20154 24252 20156
rect 24276 20154 24332 20156
rect 24356 20154 24412 20156
rect 24116 20102 24162 20154
rect 24162 20102 24172 20154
rect 24196 20102 24226 20154
rect 24226 20102 24238 20154
rect 24238 20102 24252 20154
rect 24276 20102 24290 20154
rect 24290 20102 24302 20154
rect 24302 20102 24332 20154
rect 24356 20102 24366 20154
rect 24366 20102 24412 20154
rect 24116 20100 24172 20102
rect 24196 20100 24252 20102
rect 24276 20100 24332 20102
rect 24356 20100 24412 20102
rect 23938 19372 23994 19408
rect 23938 19352 23940 19372
rect 23940 19352 23992 19372
rect 23992 19352 23994 19372
rect 24950 21392 25006 21448
rect 24116 19066 24172 19068
rect 24196 19066 24252 19068
rect 24276 19066 24332 19068
rect 24356 19066 24412 19068
rect 24116 19014 24162 19066
rect 24162 19014 24172 19066
rect 24196 19014 24226 19066
rect 24226 19014 24238 19066
rect 24238 19014 24252 19066
rect 24276 19014 24290 19066
rect 24290 19014 24302 19066
rect 24302 19014 24332 19066
rect 24356 19014 24366 19066
rect 24366 19014 24412 19066
rect 24116 19012 24172 19014
rect 24196 19012 24252 19014
rect 24276 19012 24332 19014
rect 24356 19012 24412 19014
rect 23938 18400 23994 18456
rect 24858 18944 24914 19000
rect 25502 22072 25558 22128
rect 25778 20440 25834 20496
rect 24116 17978 24172 17980
rect 24196 17978 24252 17980
rect 24276 17978 24332 17980
rect 24356 17978 24412 17980
rect 24116 17926 24162 17978
rect 24162 17926 24172 17978
rect 24196 17926 24226 17978
rect 24226 17926 24238 17978
rect 24238 17926 24252 17978
rect 24276 17926 24290 17978
rect 24290 17926 24302 17978
rect 24302 17926 24332 17978
rect 24356 17926 24366 17978
rect 24366 17926 24412 17978
rect 24116 17924 24172 17926
rect 24196 17924 24252 17926
rect 24276 17924 24332 17926
rect 24356 17924 24412 17926
rect 23294 14456 23350 14512
rect 23294 14068 23350 14104
rect 23294 14048 23296 14068
rect 23296 14048 23348 14068
rect 23348 14048 23350 14068
rect 23018 11600 23074 11656
rect 24116 16890 24172 16892
rect 24196 16890 24252 16892
rect 24276 16890 24332 16892
rect 24356 16890 24412 16892
rect 24116 16838 24162 16890
rect 24162 16838 24172 16890
rect 24196 16838 24226 16890
rect 24226 16838 24238 16890
rect 24238 16838 24252 16890
rect 24276 16838 24290 16890
rect 24290 16838 24302 16890
rect 24302 16838 24332 16890
rect 24356 16838 24366 16890
rect 24366 16838 24412 16890
rect 24116 16836 24172 16838
rect 24196 16836 24252 16838
rect 24276 16836 24332 16838
rect 24356 16836 24412 16838
rect 24116 15802 24172 15804
rect 24196 15802 24252 15804
rect 24276 15802 24332 15804
rect 24356 15802 24412 15804
rect 24116 15750 24162 15802
rect 24162 15750 24172 15802
rect 24196 15750 24226 15802
rect 24226 15750 24238 15802
rect 24238 15750 24252 15802
rect 24276 15750 24290 15802
rect 24290 15750 24302 15802
rect 24302 15750 24332 15802
rect 24356 15750 24366 15802
rect 24366 15750 24412 15802
rect 24116 15748 24172 15750
rect 24196 15748 24252 15750
rect 24276 15748 24332 15750
rect 24356 15748 24412 15750
rect 24116 14714 24172 14716
rect 24196 14714 24252 14716
rect 24276 14714 24332 14716
rect 24356 14714 24412 14716
rect 24116 14662 24162 14714
rect 24162 14662 24172 14714
rect 24196 14662 24226 14714
rect 24226 14662 24238 14714
rect 24238 14662 24252 14714
rect 24276 14662 24290 14714
rect 24290 14662 24302 14714
rect 24302 14662 24332 14714
rect 24356 14662 24366 14714
rect 24366 14662 24412 14714
rect 24116 14660 24172 14662
rect 24196 14660 24252 14662
rect 24276 14660 24332 14662
rect 24356 14660 24412 14662
rect 23754 14184 23810 14240
rect 24766 14456 24822 14512
rect 24116 13626 24172 13628
rect 24196 13626 24252 13628
rect 24276 13626 24332 13628
rect 24356 13626 24412 13628
rect 24116 13574 24162 13626
rect 24162 13574 24172 13626
rect 24196 13574 24226 13626
rect 24226 13574 24238 13626
rect 24238 13574 24252 13626
rect 24276 13574 24290 13626
rect 24290 13574 24302 13626
rect 24302 13574 24332 13626
rect 24356 13574 24366 13626
rect 24366 13574 24412 13626
rect 24116 13572 24172 13574
rect 24196 13572 24252 13574
rect 24276 13572 24332 13574
rect 24356 13572 24412 13574
rect 24398 13368 24454 13424
rect 23386 12416 23442 12472
rect 24116 12538 24172 12540
rect 24196 12538 24252 12540
rect 24276 12538 24332 12540
rect 24356 12538 24412 12540
rect 24116 12486 24162 12538
rect 24162 12486 24172 12538
rect 24196 12486 24226 12538
rect 24226 12486 24238 12538
rect 24238 12486 24252 12538
rect 24276 12486 24290 12538
rect 24290 12486 24302 12538
rect 24302 12486 24332 12538
rect 24356 12486 24366 12538
rect 24366 12486 24412 12538
rect 24116 12484 24172 12486
rect 24196 12484 24252 12486
rect 24276 12484 24332 12486
rect 24356 12484 24412 12486
rect 26698 19760 26754 19816
rect 26514 19372 26570 19408
rect 26514 19352 26516 19372
rect 26516 19352 26568 19372
rect 26568 19352 26570 19372
rect 25410 14456 25466 14512
rect 25502 14220 25504 14240
rect 25504 14220 25556 14240
rect 25556 14220 25558 14240
rect 25502 14184 25558 14220
rect 25686 13252 25742 13288
rect 25686 13232 25688 13252
rect 25688 13232 25740 13252
rect 25740 13232 25742 13252
rect 23662 11600 23718 11656
rect 19484 5466 19540 5468
rect 19564 5466 19620 5468
rect 19644 5466 19700 5468
rect 19724 5466 19780 5468
rect 19484 5414 19530 5466
rect 19530 5414 19540 5466
rect 19564 5414 19594 5466
rect 19594 5414 19606 5466
rect 19606 5414 19620 5466
rect 19644 5414 19658 5466
rect 19658 5414 19670 5466
rect 19670 5414 19700 5466
rect 19724 5414 19734 5466
rect 19734 5414 19780 5466
rect 19484 5412 19540 5414
rect 19564 5412 19620 5414
rect 19644 5412 19700 5414
rect 19724 5412 19780 5414
rect 24116 11450 24172 11452
rect 24196 11450 24252 11452
rect 24276 11450 24332 11452
rect 24356 11450 24412 11452
rect 24116 11398 24162 11450
rect 24162 11398 24172 11450
rect 24196 11398 24226 11450
rect 24226 11398 24238 11450
rect 24238 11398 24252 11450
rect 24276 11398 24290 11450
rect 24290 11398 24302 11450
rect 24302 11398 24332 11450
rect 24356 11398 24366 11450
rect 24366 11398 24412 11450
rect 24116 11396 24172 11398
rect 24196 11396 24252 11398
rect 24276 11396 24332 11398
rect 24356 11396 24412 11398
rect 24116 10362 24172 10364
rect 24196 10362 24252 10364
rect 24276 10362 24332 10364
rect 24356 10362 24412 10364
rect 24116 10310 24162 10362
rect 24162 10310 24172 10362
rect 24196 10310 24226 10362
rect 24226 10310 24238 10362
rect 24238 10310 24252 10362
rect 24276 10310 24290 10362
rect 24290 10310 24302 10362
rect 24302 10310 24332 10362
rect 24356 10310 24366 10362
rect 24366 10310 24412 10362
rect 24116 10308 24172 10310
rect 24196 10308 24252 10310
rect 24276 10308 24332 10310
rect 24356 10308 24412 10310
rect 24116 9274 24172 9276
rect 24196 9274 24252 9276
rect 24276 9274 24332 9276
rect 24356 9274 24412 9276
rect 24116 9222 24162 9274
rect 24162 9222 24172 9274
rect 24196 9222 24226 9274
rect 24226 9222 24238 9274
rect 24238 9222 24252 9274
rect 24276 9222 24290 9274
rect 24290 9222 24302 9274
rect 24302 9222 24332 9274
rect 24356 9222 24366 9274
rect 24366 9222 24412 9274
rect 24116 9220 24172 9222
rect 24196 9220 24252 9222
rect 24276 9220 24332 9222
rect 24356 9220 24412 9222
rect 24116 8186 24172 8188
rect 24196 8186 24252 8188
rect 24276 8186 24332 8188
rect 24356 8186 24412 8188
rect 24116 8134 24162 8186
rect 24162 8134 24172 8186
rect 24196 8134 24226 8186
rect 24226 8134 24238 8186
rect 24238 8134 24252 8186
rect 24276 8134 24290 8186
rect 24290 8134 24302 8186
rect 24302 8134 24332 8186
rect 24356 8134 24366 8186
rect 24366 8134 24412 8186
rect 24116 8132 24172 8134
rect 24196 8132 24252 8134
rect 24276 8132 24332 8134
rect 24356 8132 24412 8134
rect 24116 7098 24172 7100
rect 24196 7098 24252 7100
rect 24276 7098 24332 7100
rect 24356 7098 24412 7100
rect 24116 7046 24162 7098
rect 24162 7046 24172 7098
rect 24196 7046 24226 7098
rect 24226 7046 24238 7098
rect 24238 7046 24252 7098
rect 24276 7046 24290 7098
rect 24290 7046 24302 7098
rect 24302 7046 24332 7098
rect 24356 7046 24366 7098
rect 24366 7046 24412 7098
rect 24116 7044 24172 7046
rect 24196 7044 24252 7046
rect 24276 7044 24332 7046
rect 24356 7044 24412 7046
rect 28262 24520 28318 24576
rect 27802 18964 27858 19000
rect 27802 18944 27804 18964
rect 27804 18944 27856 18964
rect 27856 18944 27858 18964
rect 28262 23160 28318 23216
rect 28354 21800 28410 21856
rect 28354 20440 28410 20496
rect 28354 19080 28410 19136
rect 28170 17720 28226 17776
rect 28170 17584 28226 17640
rect 28354 16360 28410 16416
rect 27986 14048 28042 14104
rect 27066 12688 27122 12744
rect 28262 13640 28318 13696
rect 28354 12300 28410 12336
rect 28354 12280 28356 12300
rect 28356 12280 28408 12300
rect 28408 12280 28410 12300
rect 28354 10920 28410 10976
rect 24116 6010 24172 6012
rect 24196 6010 24252 6012
rect 24276 6010 24332 6012
rect 24356 6010 24412 6012
rect 24116 5958 24162 6010
rect 24162 5958 24172 6010
rect 24196 5958 24226 6010
rect 24226 5958 24238 6010
rect 24238 5958 24252 6010
rect 24276 5958 24290 6010
rect 24290 5958 24302 6010
rect 24302 5958 24332 6010
rect 24356 5958 24366 6010
rect 24366 5958 24412 6010
rect 24116 5956 24172 5958
rect 24196 5956 24252 5958
rect 24276 5956 24332 5958
rect 24356 5956 24412 5958
rect 28262 9580 28318 9616
rect 28262 9560 28264 9580
rect 28264 9560 28316 9580
rect 28316 9560 28318 9580
rect 28354 8200 28410 8256
rect 28354 6840 28410 6896
rect 28262 5516 28264 5536
rect 28264 5516 28316 5536
rect 28316 5516 28318 5536
rect 28262 5480 28318 5516
rect 24116 4922 24172 4924
rect 24196 4922 24252 4924
rect 24276 4922 24332 4924
rect 24356 4922 24412 4924
rect 24116 4870 24162 4922
rect 24162 4870 24172 4922
rect 24196 4870 24226 4922
rect 24226 4870 24238 4922
rect 24238 4870 24252 4922
rect 24276 4870 24290 4922
rect 24290 4870 24302 4922
rect 24302 4870 24332 4922
rect 24356 4870 24366 4922
rect 24366 4870 24412 4922
rect 24116 4868 24172 4870
rect 24196 4868 24252 4870
rect 24276 4868 24332 4870
rect 24356 4868 24412 4870
rect 19484 4378 19540 4380
rect 19564 4378 19620 4380
rect 19644 4378 19700 4380
rect 19724 4378 19780 4380
rect 19484 4326 19530 4378
rect 19530 4326 19540 4378
rect 19564 4326 19594 4378
rect 19594 4326 19606 4378
rect 19606 4326 19620 4378
rect 19644 4326 19658 4378
rect 19658 4326 19670 4378
rect 19670 4326 19700 4378
rect 19724 4326 19734 4378
rect 19734 4326 19780 4378
rect 19484 4324 19540 4326
rect 19564 4324 19620 4326
rect 19644 4324 19700 4326
rect 19724 4324 19780 4326
rect 28354 4120 28410 4176
rect 24116 3834 24172 3836
rect 24196 3834 24252 3836
rect 24276 3834 24332 3836
rect 24356 3834 24412 3836
rect 24116 3782 24162 3834
rect 24162 3782 24172 3834
rect 24196 3782 24226 3834
rect 24226 3782 24238 3834
rect 24238 3782 24252 3834
rect 24276 3782 24290 3834
rect 24290 3782 24302 3834
rect 24302 3782 24332 3834
rect 24356 3782 24366 3834
rect 24366 3782 24412 3834
rect 24116 3780 24172 3782
rect 24196 3780 24252 3782
rect 24276 3780 24332 3782
rect 24356 3780 24412 3782
rect 19484 3290 19540 3292
rect 19564 3290 19620 3292
rect 19644 3290 19700 3292
rect 19724 3290 19780 3292
rect 19484 3238 19530 3290
rect 19530 3238 19540 3290
rect 19564 3238 19594 3290
rect 19594 3238 19606 3290
rect 19606 3238 19620 3290
rect 19644 3238 19658 3290
rect 19658 3238 19670 3290
rect 19670 3238 19700 3290
rect 19724 3238 19734 3290
rect 19734 3238 19780 3290
rect 19484 3236 19540 3238
rect 19564 3236 19620 3238
rect 19644 3236 19700 3238
rect 19724 3236 19780 3238
rect 24116 2746 24172 2748
rect 24196 2746 24252 2748
rect 24276 2746 24332 2748
rect 24356 2746 24412 2748
rect 24116 2694 24162 2746
rect 24162 2694 24172 2746
rect 24196 2694 24226 2746
rect 24226 2694 24238 2746
rect 24238 2694 24252 2746
rect 24276 2694 24290 2746
rect 24290 2694 24302 2746
rect 24302 2694 24332 2746
rect 24356 2694 24366 2746
rect 24366 2694 24412 2746
rect 24116 2692 24172 2694
rect 24196 2692 24252 2694
rect 24276 2692 24332 2694
rect 24356 2692 24412 2694
rect 28354 2796 28356 2816
rect 28356 2796 28408 2816
rect 28408 2796 28410 2816
rect 28354 2760 28410 2796
rect 10220 2202 10276 2204
rect 10300 2202 10356 2204
rect 10380 2202 10436 2204
rect 10460 2202 10516 2204
rect 10220 2150 10266 2202
rect 10266 2150 10276 2202
rect 10300 2150 10330 2202
rect 10330 2150 10342 2202
rect 10342 2150 10356 2202
rect 10380 2150 10394 2202
rect 10394 2150 10406 2202
rect 10406 2150 10436 2202
rect 10460 2150 10470 2202
rect 10470 2150 10516 2202
rect 10220 2148 10276 2150
rect 10300 2148 10356 2150
rect 10380 2148 10436 2150
rect 10460 2148 10516 2150
rect 19484 2202 19540 2204
rect 19564 2202 19620 2204
rect 19644 2202 19700 2204
rect 19724 2202 19780 2204
rect 19484 2150 19530 2202
rect 19530 2150 19540 2202
rect 19564 2150 19594 2202
rect 19594 2150 19606 2202
rect 19606 2150 19620 2202
rect 19644 2150 19658 2202
rect 19658 2150 19670 2202
rect 19670 2150 19700 2202
rect 19724 2150 19734 2202
rect 19734 2150 19780 2202
rect 19484 2148 19540 2150
rect 19564 2148 19620 2150
rect 19644 2148 19700 2150
rect 19724 2148 19780 2150
rect 27526 40 27582 96
<< metal3 >>
rect 0 28658 800 28688
rect 1393 28658 1459 28661
rect 0 28656 1459 28658
rect 0 28600 1398 28656
rect 1454 28600 1459 28656
rect 0 28598 1459 28600
rect 0 28568 800 28598
rect 1393 28595 1459 28598
rect 27521 28658 27587 28661
rect 29200 28658 30000 28688
rect 27521 28656 30000 28658
rect 27521 28600 27526 28656
rect 27582 28600 30000 28656
rect 27521 28598 30000 28600
rect 27521 28595 27587 28598
rect 29200 28568 30000 28598
rect 5576 27776 5896 27777
rect 5576 27712 5584 27776
rect 5648 27712 5664 27776
rect 5728 27712 5744 27776
rect 5808 27712 5824 27776
rect 5888 27712 5896 27776
rect 5576 27711 5896 27712
rect 14840 27776 15160 27777
rect 14840 27712 14848 27776
rect 14912 27712 14928 27776
rect 14992 27712 15008 27776
rect 15072 27712 15088 27776
rect 15152 27712 15160 27776
rect 14840 27711 15160 27712
rect 24104 27776 24424 27777
rect 24104 27712 24112 27776
rect 24176 27712 24192 27776
rect 24256 27712 24272 27776
rect 24336 27712 24352 27776
rect 24416 27712 24424 27776
rect 24104 27711 24424 27712
rect 0 27298 800 27328
rect 1393 27298 1459 27301
rect 0 27296 1459 27298
rect 0 27240 1398 27296
rect 1454 27240 1459 27296
rect 0 27238 1459 27240
rect 0 27208 800 27238
rect 1393 27235 1459 27238
rect 10208 27232 10528 27233
rect 10208 27168 10216 27232
rect 10280 27168 10296 27232
rect 10360 27168 10376 27232
rect 10440 27168 10456 27232
rect 10520 27168 10528 27232
rect 10208 27167 10528 27168
rect 19472 27232 19792 27233
rect 19472 27168 19480 27232
rect 19544 27168 19560 27232
rect 19624 27168 19640 27232
rect 19704 27168 19720 27232
rect 19784 27168 19792 27232
rect 29200 27208 30000 27328
rect 19472 27167 19792 27168
rect 5576 26688 5896 26689
rect 5576 26624 5584 26688
rect 5648 26624 5664 26688
rect 5728 26624 5744 26688
rect 5808 26624 5824 26688
rect 5888 26624 5896 26688
rect 5576 26623 5896 26624
rect 14840 26688 15160 26689
rect 14840 26624 14848 26688
rect 14912 26624 14928 26688
rect 14992 26624 15008 26688
rect 15072 26624 15088 26688
rect 15152 26624 15160 26688
rect 14840 26623 15160 26624
rect 24104 26688 24424 26689
rect 24104 26624 24112 26688
rect 24176 26624 24192 26688
rect 24256 26624 24272 26688
rect 24336 26624 24352 26688
rect 24416 26624 24424 26688
rect 24104 26623 24424 26624
rect 25129 26346 25195 26349
rect 25497 26346 25563 26349
rect 25630 26346 25636 26348
rect 25129 26344 25636 26346
rect 25129 26288 25134 26344
rect 25190 26288 25502 26344
rect 25558 26288 25636 26344
rect 25129 26286 25636 26288
rect 25129 26283 25195 26286
rect 25497 26283 25563 26286
rect 25630 26284 25636 26286
rect 25700 26284 25706 26348
rect 10208 26144 10528 26145
rect 10208 26080 10216 26144
rect 10280 26080 10296 26144
rect 10360 26080 10376 26144
rect 10440 26080 10456 26144
rect 10520 26080 10528 26144
rect 10208 26079 10528 26080
rect 19472 26144 19792 26145
rect 19472 26080 19480 26144
rect 19544 26080 19560 26144
rect 19624 26080 19640 26144
rect 19704 26080 19720 26144
rect 19784 26080 19792 26144
rect 19472 26079 19792 26080
rect 0 25938 800 25968
rect 1669 25938 1735 25941
rect 0 25936 1735 25938
rect 0 25880 1674 25936
rect 1730 25880 1735 25936
rect 0 25878 1735 25880
rect 0 25848 800 25878
rect 1669 25875 1735 25878
rect 29200 25848 30000 25968
rect 5576 25600 5896 25601
rect 5576 25536 5584 25600
rect 5648 25536 5664 25600
rect 5728 25536 5744 25600
rect 5808 25536 5824 25600
rect 5888 25536 5896 25600
rect 5576 25535 5896 25536
rect 14840 25600 15160 25601
rect 14840 25536 14848 25600
rect 14912 25536 14928 25600
rect 14992 25536 15008 25600
rect 15072 25536 15088 25600
rect 15152 25536 15160 25600
rect 14840 25535 15160 25536
rect 24104 25600 24424 25601
rect 24104 25536 24112 25600
rect 24176 25536 24192 25600
rect 24256 25536 24272 25600
rect 24336 25536 24352 25600
rect 24416 25536 24424 25600
rect 24104 25535 24424 25536
rect 17309 25394 17375 25397
rect 21081 25394 21147 25397
rect 17309 25392 21147 25394
rect 17309 25336 17314 25392
rect 17370 25336 21086 25392
rect 21142 25336 21147 25392
rect 17309 25334 21147 25336
rect 17309 25331 17375 25334
rect 21081 25331 21147 25334
rect 10208 25056 10528 25057
rect 10208 24992 10216 25056
rect 10280 24992 10296 25056
rect 10360 24992 10376 25056
rect 10440 24992 10456 25056
rect 10520 24992 10528 25056
rect 10208 24991 10528 24992
rect 19472 25056 19792 25057
rect 19472 24992 19480 25056
rect 19544 24992 19560 25056
rect 19624 24992 19640 25056
rect 19704 24992 19720 25056
rect 19784 24992 19792 25056
rect 19472 24991 19792 24992
rect 16297 24986 16363 24989
rect 16430 24986 16436 24988
rect 16297 24984 16436 24986
rect 16297 24928 16302 24984
rect 16358 24928 16436 24984
rect 16297 24926 16436 24928
rect 16297 24923 16363 24926
rect 16430 24924 16436 24926
rect 16500 24924 16506 24988
rect 0 24488 800 24608
rect 28257 24578 28323 24581
rect 29200 24578 30000 24608
rect 28257 24576 30000 24578
rect 28257 24520 28262 24576
rect 28318 24520 30000 24576
rect 28257 24518 30000 24520
rect 28257 24515 28323 24518
rect 5576 24512 5896 24513
rect 5576 24448 5584 24512
rect 5648 24448 5664 24512
rect 5728 24448 5744 24512
rect 5808 24448 5824 24512
rect 5888 24448 5896 24512
rect 5576 24447 5896 24448
rect 14840 24512 15160 24513
rect 14840 24448 14848 24512
rect 14912 24448 14928 24512
rect 14992 24448 15008 24512
rect 15072 24448 15088 24512
rect 15152 24448 15160 24512
rect 14840 24447 15160 24448
rect 24104 24512 24424 24513
rect 24104 24448 24112 24512
rect 24176 24448 24192 24512
rect 24256 24448 24272 24512
rect 24336 24448 24352 24512
rect 24416 24448 24424 24512
rect 29200 24488 30000 24518
rect 24104 24447 24424 24448
rect 15745 24170 15811 24173
rect 20713 24170 20779 24173
rect 15745 24168 20779 24170
rect 15745 24112 15750 24168
rect 15806 24112 20718 24168
rect 20774 24112 20779 24168
rect 15745 24110 20779 24112
rect 15745 24107 15811 24110
rect 20713 24107 20779 24110
rect 10208 23968 10528 23969
rect 10208 23904 10216 23968
rect 10280 23904 10296 23968
rect 10360 23904 10376 23968
rect 10440 23904 10456 23968
rect 10520 23904 10528 23968
rect 10208 23903 10528 23904
rect 19472 23968 19792 23969
rect 19472 23904 19480 23968
rect 19544 23904 19560 23968
rect 19624 23904 19640 23968
rect 19704 23904 19720 23968
rect 19784 23904 19792 23968
rect 19472 23903 19792 23904
rect 5576 23424 5896 23425
rect 5576 23360 5584 23424
rect 5648 23360 5664 23424
rect 5728 23360 5744 23424
rect 5808 23360 5824 23424
rect 5888 23360 5896 23424
rect 5576 23359 5896 23360
rect 14840 23424 15160 23425
rect 14840 23360 14848 23424
rect 14912 23360 14928 23424
rect 14992 23360 15008 23424
rect 15072 23360 15088 23424
rect 15152 23360 15160 23424
rect 14840 23359 15160 23360
rect 24104 23424 24424 23425
rect 24104 23360 24112 23424
rect 24176 23360 24192 23424
rect 24256 23360 24272 23424
rect 24336 23360 24352 23424
rect 24416 23360 24424 23424
rect 24104 23359 24424 23360
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 28257 23218 28323 23221
rect 29200 23218 30000 23248
rect 28257 23216 30000 23218
rect 28257 23160 28262 23216
rect 28318 23160 30000 23216
rect 28257 23158 30000 23160
rect 28257 23155 28323 23158
rect 29200 23128 30000 23158
rect 10208 22880 10528 22881
rect 10208 22816 10216 22880
rect 10280 22816 10296 22880
rect 10360 22816 10376 22880
rect 10440 22816 10456 22880
rect 10520 22816 10528 22880
rect 10208 22815 10528 22816
rect 19472 22880 19792 22881
rect 19472 22816 19480 22880
rect 19544 22816 19560 22880
rect 19624 22816 19640 22880
rect 19704 22816 19720 22880
rect 19784 22816 19792 22880
rect 19472 22815 19792 22816
rect 5576 22336 5896 22337
rect 5576 22272 5584 22336
rect 5648 22272 5664 22336
rect 5728 22272 5744 22336
rect 5808 22272 5824 22336
rect 5888 22272 5896 22336
rect 5576 22271 5896 22272
rect 14840 22336 15160 22337
rect 14840 22272 14848 22336
rect 14912 22272 14928 22336
rect 14992 22272 15008 22336
rect 15072 22272 15088 22336
rect 15152 22272 15160 22336
rect 14840 22271 15160 22272
rect 24104 22336 24424 22337
rect 24104 22272 24112 22336
rect 24176 22272 24192 22336
rect 24256 22272 24272 22336
rect 24336 22272 24352 22336
rect 24416 22272 24424 22336
rect 24104 22271 24424 22272
rect 24301 22130 24367 22133
rect 25497 22130 25563 22133
rect 24301 22128 25563 22130
rect 24301 22072 24306 22128
rect 24362 22072 25502 22128
rect 25558 22072 25563 22128
rect 24301 22070 25563 22072
rect 24301 22067 24367 22070
rect 25497 22067 25563 22070
rect 24301 21994 24367 21997
rect 25037 21994 25103 21997
rect 24301 21992 25103 21994
rect 24301 21936 24306 21992
rect 24362 21936 25042 21992
rect 25098 21936 25103 21992
rect 24301 21934 25103 21936
rect 24301 21931 24367 21934
rect 25037 21931 25103 21934
rect 0 21858 800 21888
rect 1393 21858 1459 21861
rect 0 21856 1459 21858
rect 0 21800 1398 21856
rect 1454 21800 1459 21856
rect 0 21798 1459 21800
rect 0 21768 800 21798
rect 1393 21795 1459 21798
rect 28349 21858 28415 21861
rect 29200 21858 30000 21888
rect 28349 21856 30000 21858
rect 28349 21800 28354 21856
rect 28410 21800 30000 21856
rect 28349 21798 30000 21800
rect 28349 21795 28415 21798
rect 10208 21792 10528 21793
rect 10208 21728 10216 21792
rect 10280 21728 10296 21792
rect 10360 21728 10376 21792
rect 10440 21728 10456 21792
rect 10520 21728 10528 21792
rect 10208 21727 10528 21728
rect 19472 21792 19792 21793
rect 19472 21728 19480 21792
rect 19544 21728 19560 21792
rect 19624 21728 19640 21792
rect 19704 21728 19720 21792
rect 19784 21728 19792 21792
rect 29200 21768 30000 21798
rect 19472 21727 19792 21728
rect 22921 21450 22987 21453
rect 24945 21450 25011 21453
rect 22921 21448 25011 21450
rect 22921 21392 22926 21448
rect 22982 21392 24950 21448
rect 25006 21392 25011 21448
rect 22921 21390 25011 21392
rect 22921 21387 22987 21390
rect 24945 21387 25011 21390
rect 5576 21248 5896 21249
rect 5576 21184 5584 21248
rect 5648 21184 5664 21248
rect 5728 21184 5744 21248
rect 5808 21184 5824 21248
rect 5888 21184 5896 21248
rect 5576 21183 5896 21184
rect 14840 21248 15160 21249
rect 14840 21184 14848 21248
rect 14912 21184 14928 21248
rect 14992 21184 15008 21248
rect 15072 21184 15088 21248
rect 15152 21184 15160 21248
rect 14840 21183 15160 21184
rect 24104 21248 24424 21249
rect 24104 21184 24112 21248
rect 24176 21184 24192 21248
rect 24256 21184 24272 21248
rect 24336 21184 24352 21248
rect 24416 21184 24424 21248
rect 24104 21183 24424 21184
rect 12893 21042 12959 21045
rect 14733 21042 14799 21045
rect 12893 21040 14799 21042
rect 12893 20984 12898 21040
rect 12954 20984 14738 21040
rect 14794 20984 14799 21040
rect 12893 20982 14799 20984
rect 12893 20979 12959 20982
rect 14733 20979 14799 20982
rect 14181 20906 14247 20909
rect 14590 20906 14596 20908
rect 14181 20904 14596 20906
rect 14181 20848 14186 20904
rect 14242 20848 14596 20904
rect 14181 20846 14596 20848
rect 14181 20843 14247 20846
rect 14590 20844 14596 20846
rect 14660 20844 14666 20908
rect 10208 20704 10528 20705
rect 10208 20640 10216 20704
rect 10280 20640 10296 20704
rect 10360 20640 10376 20704
rect 10440 20640 10456 20704
rect 10520 20640 10528 20704
rect 10208 20639 10528 20640
rect 19472 20704 19792 20705
rect 19472 20640 19480 20704
rect 19544 20640 19560 20704
rect 19624 20640 19640 20704
rect 19704 20640 19720 20704
rect 19784 20640 19792 20704
rect 19472 20639 19792 20640
rect 0 20408 800 20528
rect 18873 20498 18939 20501
rect 25773 20498 25839 20501
rect 18873 20496 25839 20498
rect 18873 20440 18878 20496
rect 18934 20440 25778 20496
rect 25834 20440 25839 20496
rect 18873 20438 25839 20440
rect 18873 20435 18939 20438
rect 25773 20435 25839 20438
rect 28349 20498 28415 20501
rect 29200 20498 30000 20528
rect 28349 20496 30000 20498
rect 28349 20440 28354 20496
rect 28410 20440 30000 20496
rect 28349 20438 30000 20440
rect 28349 20435 28415 20438
rect 29200 20408 30000 20438
rect 5576 20160 5896 20161
rect 5576 20096 5584 20160
rect 5648 20096 5664 20160
rect 5728 20096 5744 20160
rect 5808 20096 5824 20160
rect 5888 20096 5896 20160
rect 5576 20095 5896 20096
rect 14840 20160 15160 20161
rect 14840 20096 14848 20160
rect 14912 20096 14928 20160
rect 14992 20096 15008 20160
rect 15072 20096 15088 20160
rect 15152 20096 15160 20160
rect 14840 20095 15160 20096
rect 24104 20160 24424 20161
rect 24104 20096 24112 20160
rect 24176 20096 24192 20160
rect 24256 20096 24272 20160
rect 24336 20096 24352 20160
rect 24416 20096 24424 20160
rect 24104 20095 24424 20096
rect 18413 19954 18479 19957
rect 18873 19954 18939 19957
rect 15702 19952 18939 19954
rect 15702 19896 18418 19952
rect 18474 19896 18878 19952
rect 18934 19896 18939 19952
rect 15702 19894 18939 19896
rect 12065 19818 12131 19821
rect 12709 19818 12775 19821
rect 15702 19818 15762 19894
rect 18413 19891 18479 19894
rect 18873 19891 18939 19894
rect 12065 19816 15762 19818
rect 12065 19760 12070 19816
rect 12126 19760 12714 19816
rect 12770 19760 15762 19816
rect 12065 19758 15762 19760
rect 15837 19818 15903 19821
rect 26693 19818 26759 19821
rect 15837 19816 26759 19818
rect 15837 19760 15842 19816
rect 15898 19760 26698 19816
rect 26754 19760 26759 19816
rect 15837 19758 26759 19760
rect 12065 19755 12131 19758
rect 12709 19755 12775 19758
rect 15837 19755 15903 19758
rect 26693 19755 26759 19758
rect 21449 19682 21515 19685
rect 22277 19682 22343 19685
rect 21449 19680 22343 19682
rect 21449 19624 21454 19680
rect 21510 19624 22282 19680
rect 22338 19624 22343 19680
rect 21449 19622 22343 19624
rect 21449 19619 21515 19622
rect 22277 19619 22343 19622
rect 10208 19616 10528 19617
rect 10208 19552 10216 19616
rect 10280 19552 10296 19616
rect 10360 19552 10376 19616
rect 10440 19552 10456 19616
rect 10520 19552 10528 19616
rect 10208 19551 10528 19552
rect 19472 19616 19792 19617
rect 19472 19552 19480 19616
rect 19544 19552 19560 19616
rect 19624 19552 19640 19616
rect 19704 19552 19720 19616
rect 19784 19552 19792 19616
rect 19472 19551 19792 19552
rect 23933 19410 23999 19413
rect 26509 19410 26575 19413
rect 23933 19408 26575 19410
rect 23933 19352 23938 19408
rect 23994 19352 26514 19408
rect 26570 19352 26575 19408
rect 23933 19350 26575 19352
rect 23933 19347 23999 19350
rect 26509 19347 26575 19350
rect 10317 19274 10383 19277
rect 22185 19274 22251 19277
rect 10317 19272 22251 19274
rect 10317 19216 10322 19272
rect 10378 19216 22190 19272
rect 22246 19216 22251 19272
rect 10317 19214 22251 19216
rect 10317 19211 10383 19214
rect 22185 19211 22251 19214
rect 0 19048 800 19168
rect 28349 19138 28415 19141
rect 29200 19138 30000 19168
rect 28349 19136 30000 19138
rect 28349 19080 28354 19136
rect 28410 19080 30000 19136
rect 28349 19078 30000 19080
rect 28349 19075 28415 19078
rect 5576 19072 5896 19073
rect 5576 19008 5584 19072
rect 5648 19008 5664 19072
rect 5728 19008 5744 19072
rect 5808 19008 5824 19072
rect 5888 19008 5896 19072
rect 5576 19007 5896 19008
rect 14840 19072 15160 19073
rect 14840 19008 14848 19072
rect 14912 19008 14928 19072
rect 14992 19008 15008 19072
rect 15072 19008 15088 19072
rect 15152 19008 15160 19072
rect 14840 19007 15160 19008
rect 24104 19072 24424 19073
rect 24104 19008 24112 19072
rect 24176 19008 24192 19072
rect 24256 19008 24272 19072
rect 24336 19008 24352 19072
rect 24416 19008 24424 19072
rect 29200 19048 30000 19078
rect 24104 19007 24424 19008
rect 24853 19002 24919 19005
rect 27797 19002 27863 19005
rect 24853 19000 27863 19002
rect 24853 18944 24858 19000
rect 24914 18944 27802 19000
rect 27858 18944 27863 19000
rect 24853 18942 27863 18944
rect 24853 18939 24919 18942
rect 27797 18939 27863 18942
rect 10208 18528 10528 18529
rect 10208 18464 10216 18528
rect 10280 18464 10296 18528
rect 10360 18464 10376 18528
rect 10440 18464 10456 18528
rect 10520 18464 10528 18528
rect 10208 18463 10528 18464
rect 19472 18528 19792 18529
rect 19472 18464 19480 18528
rect 19544 18464 19560 18528
rect 19624 18464 19640 18528
rect 19704 18464 19720 18528
rect 19784 18464 19792 18528
rect 19472 18463 19792 18464
rect 16430 18396 16436 18460
rect 16500 18458 16506 18460
rect 16849 18458 16915 18461
rect 16500 18456 16915 18458
rect 16500 18400 16854 18456
rect 16910 18400 16915 18456
rect 16500 18398 16915 18400
rect 16500 18396 16506 18398
rect 16849 18395 16915 18398
rect 19977 18458 20043 18461
rect 23289 18458 23355 18461
rect 23933 18458 23999 18461
rect 19977 18456 23999 18458
rect 19977 18400 19982 18456
rect 20038 18400 23294 18456
rect 23350 18400 23938 18456
rect 23994 18400 23999 18456
rect 19977 18398 23999 18400
rect 19977 18395 20043 18398
rect 23289 18395 23355 18398
rect 23933 18395 23999 18398
rect 10777 18322 10843 18325
rect 11697 18322 11763 18325
rect 17585 18322 17651 18325
rect 10777 18320 17651 18322
rect 10777 18264 10782 18320
rect 10838 18264 11702 18320
rect 11758 18264 17590 18320
rect 17646 18264 17651 18320
rect 10777 18262 17651 18264
rect 10777 18259 10843 18262
rect 11697 18259 11763 18262
rect 17585 18259 17651 18262
rect 5576 17984 5896 17985
rect 5576 17920 5584 17984
rect 5648 17920 5664 17984
rect 5728 17920 5744 17984
rect 5808 17920 5824 17984
rect 5888 17920 5896 17984
rect 5576 17919 5896 17920
rect 14840 17984 15160 17985
rect 14840 17920 14848 17984
rect 14912 17920 14928 17984
rect 14992 17920 15008 17984
rect 15072 17920 15088 17984
rect 15152 17920 15160 17984
rect 14840 17919 15160 17920
rect 24104 17984 24424 17985
rect 24104 17920 24112 17984
rect 24176 17920 24192 17984
rect 24256 17920 24272 17984
rect 24336 17920 24352 17984
rect 24416 17920 24424 17984
rect 24104 17919 24424 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 15561 17778 15627 17781
rect 25630 17778 25636 17780
rect 15561 17776 25636 17778
rect 15561 17720 15566 17776
rect 15622 17720 25636 17776
rect 15561 17718 25636 17720
rect 15561 17715 15627 17718
rect 25630 17716 25636 17718
rect 25700 17716 25706 17780
rect 28165 17778 28231 17781
rect 29200 17778 30000 17808
rect 28165 17776 30000 17778
rect 28165 17720 28170 17776
rect 28226 17720 30000 17776
rect 28165 17718 30000 17720
rect 28165 17715 28231 17718
rect 29200 17688 30000 17718
rect 18597 17642 18663 17645
rect 28165 17642 28231 17645
rect 18597 17640 28231 17642
rect 18597 17584 18602 17640
rect 18658 17584 28170 17640
rect 28226 17584 28231 17640
rect 18597 17582 28231 17584
rect 18597 17579 18663 17582
rect 28165 17579 28231 17582
rect 10208 17440 10528 17441
rect 10208 17376 10216 17440
rect 10280 17376 10296 17440
rect 10360 17376 10376 17440
rect 10440 17376 10456 17440
rect 10520 17376 10528 17440
rect 10208 17375 10528 17376
rect 19472 17440 19792 17441
rect 19472 17376 19480 17440
rect 19544 17376 19560 17440
rect 19624 17376 19640 17440
rect 19704 17376 19720 17440
rect 19784 17376 19792 17440
rect 19472 17375 19792 17376
rect 11053 17234 11119 17237
rect 17953 17234 18019 17237
rect 11053 17232 18019 17234
rect 11053 17176 11058 17232
rect 11114 17176 17958 17232
rect 18014 17176 18019 17232
rect 11053 17174 18019 17176
rect 11053 17171 11119 17174
rect 17953 17171 18019 17174
rect 11421 16962 11487 16965
rect 14641 16962 14707 16965
rect 11421 16960 14707 16962
rect 11421 16904 11426 16960
rect 11482 16904 14646 16960
rect 14702 16904 14707 16960
rect 11421 16902 14707 16904
rect 11421 16899 11487 16902
rect 14641 16899 14707 16902
rect 5576 16896 5896 16897
rect 5576 16832 5584 16896
rect 5648 16832 5664 16896
rect 5728 16832 5744 16896
rect 5808 16832 5824 16896
rect 5888 16832 5896 16896
rect 5576 16831 5896 16832
rect 14840 16896 15160 16897
rect 14840 16832 14848 16896
rect 14912 16832 14928 16896
rect 14992 16832 15008 16896
rect 15072 16832 15088 16896
rect 15152 16832 15160 16896
rect 14840 16831 15160 16832
rect 24104 16896 24424 16897
rect 24104 16832 24112 16896
rect 24176 16832 24192 16896
rect 24256 16832 24272 16896
rect 24336 16832 24352 16896
rect 24416 16832 24424 16896
rect 24104 16831 24424 16832
rect 12985 16826 13051 16829
rect 12985 16824 14106 16826
rect 12985 16768 12990 16824
rect 13046 16768 14106 16824
rect 12985 16766 14106 16768
rect 12985 16763 13051 16766
rect 9765 16690 9831 16693
rect 13854 16690 13860 16692
rect 9765 16688 13860 16690
rect 9765 16632 9770 16688
rect 9826 16632 13860 16688
rect 9765 16630 13860 16632
rect 9765 16627 9831 16630
rect 13854 16628 13860 16630
rect 13924 16628 13930 16692
rect 14046 16690 14106 16766
rect 17125 16690 17191 16693
rect 14046 16688 17191 16690
rect 14046 16632 17130 16688
rect 17186 16632 17191 16688
rect 14046 16630 17191 16632
rect 17125 16627 17191 16630
rect 0 16418 800 16448
rect 1393 16418 1459 16421
rect 0 16416 1459 16418
rect 0 16360 1398 16416
rect 1454 16360 1459 16416
rect 0 16358 1459 16360
rect 0 16328 800 16358
rect 1393 16355 1459 16358
rect 11145 16418 11211 16421
rect 11881 16418 11947 16421
rect 17953 16418 18019 16421
rect 18597 16418 18663 16421
rect 11145 16416 18663 16418
rect 11145 16360 11150 16416
rect 11206 16360 11886 16416
rect 11942 16360 17958 16416
rect 18014 16360 18602 16416
rect 18658 16360 18663 16416
rect 11145 16358 18663 16360
rect 11145 16355 11211 16358
rect 11881 16355 11947 16358
rect 17953 16355 18019 16358
rect 18597 16355 18663 16358
rect 28349 16418 28415 16421
rect 29200 16418 30000 16448
rect 28349 16416 30000 16418
rect 28349 16360 28354 16416
rect 28410 16360 30000 16416
rect 28349 16358 30000 16360
rect 28349 16355 28415 16358
rect 10208 16352 10528 16353
rect 10208 16288 10216 16352
rect 10280 16288 10296 16352
rect 10360 16288 10376 16352
rect 10440 16288 10456 16352
rect 10520 16288 10528 16352
rect 10208 16287 10528 16288
rect 19472 16352 19792 16353
rect 19472 16288 19480 16352
rect 19544 16288 19560 16352
rect 19624 16288 19640 16352
rect 19704 16288 19720 16352
rect 19784 16288 19792 16352
rect 29200 16328 30000 16358
rect 19472 16287 19792 16288
rect 17125 16146 17191 16149
rect 18873 16146 18939 16149
rect 17125 16144 18939 16146
rect 17125 16088 17130 16144
rect 17186 16088 18878 16144
rect 18934 16088 18939 16144
rect 17125 16086 18939 16088
rect 17125 16083 17191 16086
rect 18873 16083 18939 16086
rect 5576 15808 5896 15809
rect 5576 15744 5584 15808
rect 5648 15744 5664 15808
rect 5728 15744 5744 15808
rect 5808 15744 5824 15808
rect 5888 15744 5896 15808
rect 5576 15743 5896 15744
rect 14840 15808 15160 15809
rect 14840 15744 14848 15808
rect 14912 15744 14928 15808
rect 14992 15744 15008 15808
rect 15072 15744 15088 15808
rect 15152 15744 15160 15808
rect 14840 15743 15160 15744
rect 24104 15808 24424 15809
rect 24104 15744 24112 15808
rect 24176 15744 24192 15808
rect 24256 15744 24272 15808
rect 24336 15744 24352 15808
rect 24416 15744 24424 15808
rect 24104 15743 24424 15744
rect 12985 15466 13051 15469
rect 13445 15466 13511 15469
rect 12985 15464 13511 15466
rect 12985 15408 12990 15464
rect 13046 15408 13450 15464
rect 13506 15408 13511 15464
rect 12985 15406 13511 15408
rect 12985 15403 13051 15406
rect 13445 15403 13511 15406
rect 17953 15466 18019 15469
rect 19926 15466 19932 15468
rect 17953 15464 19932 15466
rect 17953 15408 17958 15464
rect 18014 15408 19932 15464
rect 17953 15406 19932 15408
rect 17953 15403 18019 15406
rect 19926 15404 19932 15406
rect 19996 15404 20002 15468
rect 13169 15330 13235 15333
rect 13486 15330 13492 15332
rect 13169 15328 13492 15330
rect 13169 15272 13174 15328
rect 13230 15272 13492 15328
rect 13169 15270 13492 15272
rect 13169 15267 13235 15270
rect 13486 15268 13492 15270
rect 13556 15268 13562 15332
rect 10208 15264 10528 15265
rect 10208 15200 10216 15264
rect 10280 15200 10296 15264
rect 10360 15200 10376 15264
rect 10440 15200 10456 15264
rect 10520 15200 10528 15264
rect 10208 15199 10528 15200
rect 19472 15264 19792 15265
rect 19472 15200 19480 15264
rect 19544 15200 19560 15264
rect 19624 15200 19640 15264
rect 19704 15200 19720 15264
rect 19784 15200 19792 15264
rect 19472 15199 19792 15200
rect 11697 15194 11763 15197
rect 12893 15194 12959 15197
rect 11697 15192 14658 15194
rect 11697 15136 11702 15192
rect 11758 15136 12898 15192
rect 12954 15136 14658 15192
rect 11697 15134 14658 15136
rect 11697 15131 11763 15134
rect 12893 15131 12959 15134
rect 0 15058 800 15088
rect 4061 15058 4127 15061
rect 0 15056 4127 15058
rect 0 15000 4066 15056
rect 4122 15000 4127 15056
rect 0 14998 4127 15000
rect 0 14968 800 14998
rect 4061 14995 4127 14998
rect 13854 14996 13860 15060
rect 13924 15058 13930 15060
rect 14365 15058 14431 15061
rect 13924 15056 14431 15058
rect 13924 15000 14370 15056
rect 14426 15000 14431 15056
rect 13924 14998 14431 15000
rect 14598 15058 14658 15134
rect 14733 15058 14799 15061
rect 14598 15056 14799 15058
rect 14598 15000 14738 15056
rect 14794 15000 14799 15056
rect 14598 14998 14799 15000
rect 13924 14996 13930 14998
rect 14365 14995 14431 14998
rect 14733 14995 14799 14998
rect 29200 14968 30000 15088
rect 13077 14922 13143 14925
rect 14089 14922 14155 14925
rect 13077 14920 14155 14922
rect 13077 14864 13082 14920
rect 13138 14864 14094 14920
rect 14150 14864 14155 14920
rect 13077 14862 14155 14864
rect 13077 14859 13143 14862
rect 14089 14859 14155 14862
rect 5576 14720 5896 14721
rect 5576 14656 5584 14720
rect 5648 14656 5664 14720
rect 5728 14656 5744 14720
rect 5808 14656 5824 14720
rect 5888 14656 5896 14720
rect 5576 14655 5896 14656
rect 14840 14720 15160 14721
rect 14840 14656 14848 14720
rect 14912 14656 14928 14720
rect 14992 14656 15008 14720
rect 15072 14656 15088 14720
rect 15152 14656 15160 14720
rect 14840 14655 15160 14656
rect 24104 14720 24424 14721
rect 24104 14656 24112 14720
rect 24176 14656 24192 14720
rect 24256 14656 24272 14720
rect 24336 14656 24352 14720
rect 24416 14656 24424 14720
rect 24104 14655 24424 14656
rect 13813 14514 13879 14517
rect 14457 14514 14523 14517
rect 13813 14512 14523 14514
rect 13813 14456 13818 14512
rect 13874 14456 14462 14512
rect 14518 14456 14523 14512
rect 13813 14454 14523 14456
rect 13813 14451 13879 14454
rect 14457 14451 14523 14454
rect 23289 14514 23355 14517
rect 24761 14514 24827 14517
rect 25405 14514 25471 14517
rect 23289 14512 25471 14514
rect 23289 14456 23294 14512
rect 23350 14456 24766 14512
rect 24822 14456 25410 14512
rect 25466 14456 25471 14512
rect 23289 14454 25471 14456
rect 23289 14451 23355 14454
rect 24761 14451 24827 14454
rect 25405 14451 25471 14454
rect 6545 14378 6611 14381
rect 15285 14378 15351 14381
rect 6545 14376 15351 14378
rect 6545 14320 6550 14376
rect 6606 14320 15290 14376
rect 15346 14320 15351 14376
rect 6545 14318 15351 14320
rect 6545 14315 6611 14318
rect 15285 14315 15351 14318
rect 18689 14378 18755 14381
rect 20989 14378 21055 14381
rect 18689 14376 21055 14378
rect 18689 14320 18694 14376
rect 18750 14320 20994 14376
rect 21050 14320 21055 14376
rect 18689 14318 21055 14320
rect 18689 14315 18755 14318
rect 20989 14315 21055 14318
rect 23749 14242 23815 14245
rect 25497 14242 25563 14245
rect 23749 14240 25563 14242
rect 23749 14184 23754 14240
rect 23810 14184 25502 14240
rect 25558 14184 25563 14240
rect 23749 14182 25563 14184
rect 23749 14179 23815 14182
rect 25497 14179 25563 14182
rect 10208 14176 10528 14177
rect 10208 14112 10216 14176
rect 10280 14112 10296 14176
rect 10360 14112 10376 14176
rect 10440 14112 10456 14176
rect 10520 14112 10528 14176
rect 10208 14111 10528 14112
rect 19472 14176 19792 14177
rect 19472 14112 19480 14176
rect 19544 14112 19560 14176
rect 19624 14112 19640 14176
rect 19704 14112 19720 14176
rect 19784 14112 19792 14176
rect 19472 14111 19792 14112
rect 20897 14106 20963 14109
rect 21357 14106 21423 14109
rect 23289 14106 23355 14109
rect 27981 14106 28047 14109
rect 20897 14104 28047 14106
rect 20897 14048 20902 14104
rect 20958 14048 21362 14104
rect 21418 14048 23294 14104
rect 23350 14048 27986 14104
rect 28042 14048 28047 14104
rect 20897 14046 28047 14048
rect 20897 14043 20963 14046
rect 21357 14043 21423 14046
rect 23289 14043 23355 14046
rect 27981 14043 28047 14046
rect 11145 13970 11211 13973
rect 12249 13970 12315 13973
rect 17677 13970 17743 13973
rect 11145 13968 17743 13970
rect 11145 13912 11150 13968
rect 11206 13912 12254 13968
rect 12310 13912 17682 13968
rect 17738 13912 17743 13968
rect 11145 13910 17743 13912
rect 11145 13907 11211 13910
rect 12249 13907 12315 13910
rect 17677 13907 17743 13910
rect 8937 13834 9003 13837
rect 14641 13834 14707 13837
rect 8937 13832 14707 13834
rect 8937 13776 8942 13832
rect 8998 13776 14646 13832
rect 14702 13776 14707 13832
rect 8937 13774 14707 13776
rect 8937 13771 9003 13774
rect 14641 13771 14707 13774
rect 0 13608 800 13728
rect 28257 13698 28323 13701
rect 29200 13698 30000 13728
rect 28257 13696 30000 13698
rect 28257 13640 28262 13696
rect 28318 13640 30000 13696
rect 28257 13638 30000 13640
rect 28257 13635 28323 13638
rect 5576 13632 5896 13633
rect 5576 13568 5584 13632
rect 5648 13568 5664 13632
rect 5728 13568 5744 13632
rect 5808 13568 5824 13632
rect 5888 13568 5896 13632
rect 5576 13567 5896 13568
rect 14840 13632 15160 13633
rect 14840 13568 14848 13632
rect 14912 13568 14928 13632
rect 14992 13568 15008 13632
rect 15072 13568 15088 13632
rect 15152 13568 15160 13632
rect 14840 13567 15160 13568
rect 24104 13632 24424 13633
rect 24104 13568 24112 13632
rect 24176 13568 24192 13632
rect 24256 13568 24272 13632
rect 24336 13568 24352 13632
rect 24416 13568 24424 13632
rect 29200 13608 30000 13638
rect 24104 13567 24424 13568
rect 21449 13426 21515 13429
rect 24393 13426 24459 13429
rect 21449 13424 24459 13426
rect 21449 13368 21454 13424
rect 21510 13368 24398 13424
rect 24454 13368 24459 13424
rect 21449 13366 24459 13368
rect 21449 13363 21515 13366
rect 24393 13363 24459 13366
rect 19793 13290 19859 13293
rect 25681 13290 25747 13293
rect 19793 13288 25747 13290
rect 19793 13232 19798 13288
rect 19854 13232 25686 13288
rect 25742 13232 25747 13288
rect 19793 13230 25747 13232
rect 19793 13227 19859 13230
rect 25681 13227 25747 13230
rect 10208 13088 10528 13089
rect 10208 13024 10216 13088
rect 10280 13024 10296 13088
rect 10360 13024 10376 13088
rect 10440 13024 10456 13088
rect 10520 13024 10528 13088
rect 10208 13023 10528 13024
rect 19472 13088 19792 13089
rect 19472 13024 19480 13088
rect 19544 13024 19560 13088
rect 19624 13024 19640 13088
rect 19704 13024 19720 13088
rect 19784 13024 19792 13088
rect 19472 13023 19792 13024
rect 20529 13018 20595 13021
rect 22553 13018 22619 13021
rect 20529 13016 22619 13018
rect 20529 12960 20534 13016
rect 20590 12960 22558 13016
rect 22614 12960 22619 13016
rect 20529 12958 22619 12960
rect 20529 12955 20595 12958
rect 22553 12955 22619 12958
rect 20621 12746 20687 12749
rect 27061 12746 27127 12749
rect 20621 12744 27127 12746
rect 20621 12688 20626 12744
rect 20682 12688 27066 12744
rect 27122 12688 27127 12744
rect 20621 12686 27127 12688
rect 20621 12683 20687 12686
rect 27061 12683 27127 12686
rect 5576 12544 5896 12545
rect 5576 12480 5584 12544
rect 5648 12480 5664 12544
rect 5728 12480 5744 12544
rect 5808 12480 5824 12544
rect 5888 12480 5896 12544
rect 5576 12479 5896 12480
rect 14840 12544 15160 12545
rect 14840 12480 14848 12544
rect 14912 12480 14928 12544
rect 14992 12480 15008 12544
rect 15072 12480 15088 12544
rect 15152 12480 15160 12544
rect 14840 12479 15160 12480
rect 24104 12544 24424 12545
rect 24104 12480 24112 12544
rect 24176 12480 24192 12544
rect 24256 12480 24272 12544
rect 24336 12480 24352 12544
rect 24416 12480 24424 12544
rect 24104 12479 24424 12480
rect 22093 12474 22159 12477
rect 23381 12474 23447 12477
rect 22093 12472 23447 12474
rect 22093 12416 22098 12472
rect 22154 12416 23386 12472
rect 23442 12416 23447 12472
rect 22093 12414 23447 12416
rect 22093 12411 22159 12414
rect 23381 12411 23447 12414
rect 0 12248 800 12368
rect 11053 12338 11119 12341
rect 14273 12338 14339 12341
rect 11053 12336 14339 12338
rect 11053 12280 11058 12336
rect 11114 12280 14278 12336
rect 14334 12280 14339 12336
rect 11053 12278 14339 12280
rect 11053 12275 11119 12278
rect 14273 12275 14339 12278
rect 28349 12338 28415 12341
rect 29200 12338 30000 12368
rect 28349 12336 30000 12338
rect 28349 12280 28354 12336
rect 28410 12280 30000 12336
rect 28349 12278 30000 12280
rect 28349 12275 28415 12278
rect 29200 12248 30000 12278
rect 1761 12202 1827 12205
rect 16113 12202 16179 12205
rect 1761 12200 16179 12202
rect 1761 12144 1766 12200
rect 1822 12144 16118 12200
rect 16174 12144 16179 12200
rect 1761 12142 16179 12144
rect 1761 12139 1827 12142
rect 16113 12139 16179 12142
rect 11513 12066 11579 12069
rect 12709 12066 12775 12069
rect 13670 12066 13676 12068
rect 11513 12064 13676 12066
rect 11513 12008 11518 12064
rect 11574 12008 12714 12064
rect 12770 12008 13676 12064
rect 11513 12006 13676 12008
rect 11513 12003 11579 12006
rect 12709 12003 12775 12006
rect 13670 12004 13676 12006
rect 13740 12066 13746 12068
rect 14590 12066 14596 12068
rect 13740 12006 14596 12066
rect 13740 12004 13746 12006
rect 14590 12004 14596 12006
rect 14660 12004 14666 12068
rect 10208 12000 10528 12001
rect 10208 11936 10216 12000
rect 10280 11936 10296 12000
rect 10360 11936 10376 12000
rect 10440 11936 10456 12000
rect 10520 11936 10528 12000
rect 10208 11935 10528 11936
rect 19472 12000 19792 12001
rect 19472 11936 19480 12000
rect 19544 11936 19560 12000
rect 19624 11936 19640 12000
rect 19704 11936 19720 12000
rect 19784 11936 19792 12000
rect 19472 11935 19792 11936
rect 16297 11794 16363 11797
rect 19793 11794 19859 11797
rect 16297 11792 19859 11794
rect 16297 11736 16302 11792
rect 16358 11736 19798 11792
rect 19854 11736 19859 11792
rect 16297 11734 19859 11736
rect 16297 11731 16363 11734
rect 19793 11731 19859 11734
rect 17125 11658 17191 11661
rect 22277 11658 22343 11661
rect 17125 11656 22343 11658
rect 17125 11600 17130 11656
rect 17186 11600 22282 11656
rect 22338 11600 22343 11656
rect 17125 11598 22343 11600
rect 17125 11595 17191 11598
rect 22277 11595 22343 11598
rect 23013 11658 23079 11661
rect 23657 11658 23723 11661
rect 23013 11656 23723 11658
rect 23013 11600 23018 11656
rect 23074 11600 23662 11656
rect 23718 11600 23723 11656
rect 23013 11598 23723 11600
rect 23013 11595 23079 11598
rect 23657 11595 23723 11598
rect 5576 11456 5896 11457
rect 5576 11392 5584 11456
rect 5648 11392 5664 11456
rect 5728 11392 5744 11456
rect 5808 11392 5824 11456
rect 5888 11392 5896 11456
rect 5576 11391 5896 11392
rect 14840 11456 15160 11457
rect 14840 11392 14848 11456
rect 14912 11392 14928 11456
rect 14992 11392 15008 11456
rect 15072 11392 15088 11456
rect 15152 11392 15160 11456
rect 14840 11391 15160 11392
rect 24104 11456 24424 11457
rect 24104 11392 24112 11456
rect 24176 11392 24192 11456
rect 24256 11392 24272 11456
rect 24336 11392 24352 11456
rect 24416 11392 24424 11456
rect 24104 11391 24424 11392
rect 9673 11250 9739 11253
rect 16205 11250 16271 11253
rect 9673 11248 16271 11250
rect 9673 11192 9678 11248
rect 9734 11192 16210 11248
rect 16266 11192 16271 11248
rect 9673 11190 16271 11192
rect 9673 11187 9739 11190
rect 16205 11187 16271 11190
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 28349 10978 28415 10981
rect 29200 10978 30000 11008
rect 28349 10976 30000 10978
rect 28349 10920 28354 10976
rect 28410 10920 30000 10976
rect 28349 10918 30000 10920
rect 28349 10915 28415 10918
rect 10208 10912 10528 10913
rect 10208 10848 10216 10912
rect 10280 10848 10296 10912
rect 10360 10848 10376 10912
rect 10440 10848 10456 10912
rect 10520 10848 10528 10912
rect 10208 10847 10528 10848
rect 19472 10912 19792 10913
rect 19472 10848 19480 10912
rect 19544 10848 19560 10912
rect 19624 10848 19640 10912
rect 19704 10848 19720 10912
rect 19784 10848 19792 10912
rect 29200 10888 30000 10918
rect 19472 10847 19792 10848
rect 5576 10368 5896 10369
rect 5576 10304 5584 10368
rect 5648 10304 5664 10368
rect 5728 10304 5744 10368
rect 5808 10304 5824 10368
rect 5888 10304 5896 10368
rect 5576 10303 5896 10304
rect 14840 10368 15160 10369
rect 14840 10304 14848 10368
rect 14912 10304 14928 10368
rect 14992 10304 15008 10368
rect 15072 10304 15088 10368
rect 15152 10304 15160 10368
rect 14840 10303 15160 10304
rect 24104 10368 24424 10369
rect 24104 10304 24112 10368
rect 24176 10304 24192 10368
rect 24256 10304 24272 10368
rect 24336 10304 24352 10368
rect 24416 10304 24424 10368
rect 24104 10303 24424 10304
rect 19977 10164 20043 10165
rect 19926 10100 19932 10164
rect 19996 10162 20043 10164
rect 19996 10160 20088 10162
rect 20038 10104 20088 10160
rect 19996 10102 20088 10104
rect 19996 10100 20043 10102
rect 19977 10099 20043 10100
rect 10208 9824 10528 9825
rect 10208 9760 10216 9824
rect 10280 9760 10296 9824
rect 10360 9760 10376 9824
rect 10440 9760 10456 9824
rect 10520 9760 10528 9824
rect 10208 9759 10528 9760
rect 19472 9824 19792 9825
rect 19472 9760 19480 9824
rect 19544 9760 19560 9824
rect 19624 9760 19640 9824
rect 19704 9760 19720 9824
rect 19784 9760 19792 9824
rect 19472 9759 19792 9760
rect 0 9618 800 9648
rect 1577 9618 1643 9621
rect 0 9616 1643 9618
rect 0 9560 1582 9616
rect 1638 9560 1643 9616
rect 0 9558 1643 9560
rect 0 9528 800 9558
rect 1577 9555 1643 9558
rect 12709 9618 12775 9621
rect 15561 9618 15627 9621
rect 12709 9616 15627 9618
rect 12709 9560 12714 9616
rect 12770 9560 15566 9616
rect 15622 9560 15627 9616
rect 12709 9558 15627 9560
rect 12709 9555 12775 9558
rect 15561 9555 15627 9558
rect 28257 9618 28323 9621
rect 29200 9618 30000 9648
rect 28257 9616 30000 9618
rect 28257 9560 28262 9616
rect 28318 9560 30000 9616
rect 28257 9558 30000 9560
rect 28257 9555 28323 9558
rect 29200 9528 30000 9558
rect 5576 9280 5896 9281
rect 5576 9216 5584 9280
rect 5648 9216 5664 9280
rect 5728 9216 5744 9280
rect 5808 9216 5824 9280
rect 5888 9216 5896 9280
rect 5576 9215 5896 9216
rect 14840 9280 15160 9281
rect 14840 9216 14848 9280
rect 14912 9216 14928 9280
rect 14992 9216 15008 9280
rect 15072 9216 15088 9280
rect 15152 9216 15160 9280
rect 14840 9215 15160 9216
rect 24104 9280 24424 9281
rect 24104 9216 24112 9280
rect 24176 9216 24192 9280
rect 24256 9216 24272 9280
rect 24336 9216 24352 9280
rect 24416 9216 24424 9280
rect 24104 9215 24424 9216
rect 1761 8938 1827 8941
rect 18137 8938 18203 8941
rect 1761 8936 18203 8938
rect 1761 8880 1766 8936
rect 1822 8880 18142 8936
rect 18198 8880 18203 8936
rect 1761 8878 18203 8880
rect 1761 8875 1827 8878
rect 18137 8875 18203 8878
rect 10208 8736 10528 8737
rect 10208 8672 10216 8736
rect 10280 8672 10296 8736
rect 10360 8672 10376 8736
rect 10440 8672 10456 8736
rect 10520 8672 10528 8736
rect 10208 8671 10528 8672
rect 19472 8736 19792 8737
rect 19472 8672 19480 8736
rect 19544 8672 19560 8736
rect 19624 8672 19640 8736
rect 19704 8672 19720 8736
rect 19784 8672 19792 8736
rect 19472 8671 19792 8672
rect 13629 8668 13695 8669
rect 13629 8666 13676 8668
rect 13584 8664 13676 8666
rect 13740 8666 13746 8668
rect 16665 8666 16731 8669
rect 13740 8664 16731 8666
rect 13584 8608 13634 8664
rect 13740 8608 16670 8664
rect 16726 8608 16731 8664
rect 13584 8606 13676 8608
rect 13629 8604 13676 8606
rect 13740 8606 16731 8608
rect 13740 8604 13746 8606
rect 13629 8603 13695 8604
rect 16665 8603 16731 8606
rect 10777 8394 10843 8397
rect 15377 8394 15443 8397
rect 10777 8392 15443 8394
rect 10777 8336 10782 8392
rect 10838 8336 15382 8392
rect 15438 8336 15443 8392
rect 10777 8334 15443 8336
rect 10777 8331 10843 8334
rect 15377 8331 15443 8334
rect 0 8258 800 8288
rect 1577 8258 1643 8261
rect 0 8256 1643 8258
rect 0 8200 1582 8256
rect 1638 8200 1643 8256
rect 0 8198 1643 8200
rect 0 8168 800 8198
rect 1577 8195 1643 8198
rect 28349 8258 28415 8261
rect 29200 8258 30000 8288
rect 28349 8256 30000 8258
rect 28349 8200 28354 8256
rect 28410 8200 30000 8256
rect 28349 8198 30000 8200
rect 28349 8195 28415 8198
rect 5576 8192 5896 8193
rect 5576 8128 5584 8192
rect 5648 8128 5664 8192
rect 5728 8128 5744 8192
rect 5808 8128 5824 8192
rect 5888 8128 5896 8192
rect 5576 8127 5896 8128
rect 14840 8192 15160 8193
rect 14840 8128 14848 8192
rect 14912 8128 14928 8192
rect 14992 8128 15008 8192
rect 15072 8128 15088 8192
rect 15152 8128 15160 8192
rect 14840 8127 15160 8128
rect 24104 8192 24424 8193
rect 24104 8128 24112 8192
rect 24176 8128 24192 8192
rect 24256 8128 24272 8192
rect 24336 8128 24352 8192
rect 24416 8128 24424 8192
rect 29200 8168 30000 8198
rect 24104 8127 24424 8128
rect 10208 7648 10528 7649
rect 10208 7584 10216 7648
rect 10280 7584 10296 7648
rect 10360 7584 10376 7648
rect 10440 7584 10456 7648
rect 10520 7584 10528 7648
rect 10208 7583 10528 7584
rect 19472 7648 19792 7649
rect 19472 7584 19480 7648
rect 19544 7584 19560 7648
rect 19624 7584 19640 7648
rect 19704 7584 19720 7648
rect 19784 7584 19792 7648
rect 19472 7583 19792 7584
rect 5576 7104 5896 7105
rect 5576 7040 5584 7104
rect 5648 7040 5664 7104
rect 5728 7040 5744 7104
rect 5808 7040 5824 7104
rect 5888 7040 5896 7104
rect 5576 7039 5896 7040
rect 14840 7104 15160 7105
rect 14840 7040 14848 7104
rect 14912 7040 14928 7104
rect 14992 7040 15008 7104
rect 15072 7040 15088 7104
rect 15152 7040 15160 7104
rect 14840 7039 15160 7040
rect 24104 7104 24424 7105
rect 24104 7040 24112 7104
rect 24176 7040 24192 7104
rect 24256 7040 24272 7104
rect 24336 7040 24352 7104
rect 24416 7040 24424 7104
rect 24104 7039 24424 7040
rect 0 6808 800 6928
rect 13445 6900 13511 6901
rect 13445 6896 13492 6900
rect 13556 6898 13562 6900
rect 28349 6898 28415 6901
rect 29200 6898 30000 6928
rect 13445 6840 13450 6896
rect 13445 6836 13492 6840
rect 13556 6838 13602 6898
rect 28349 6896 30000 6898
rect 28349 6840 28354 6896
rect 28410 6840 30000 6896
rect 28349 6838 30000 6840
rect 13556 6836 13562 6838
rect 13445 6835 13511 6836
rect 28349 6835 28415 6838
rect 29200 6808 30000 6838
rect 10208 6560 10528 6561
rect 10208 6496 10216 6560
rect 10280 6496 10296 6560
rect 10360 6496 10376 6560
rect 10440 6496 10456 6560
rect 10520 6496 10528 6560
rect 10208 6495 10528 6496
rect 19472 6560 19792 6561
rect 19472 6496 19480 6560
rect 19544 6496 19560 6560
rect 19624 6496 19640 6560
rect 19704 6496 19720 6560
rect 19784 6496 19792 6560
rect 19472 6495 19792 6496
rect 5576 6016 5896 6017
rect 5576 5952 5584 6016
rect 5648 5952 5664 6016
rect 5728 5952 5744 6016
rect 5808 5952 5824 6016
rect 5888 5952 5896 6016
rect 5576 5951 5896 5952
rect 14840 6016 15160 6017
rect 14840 5952 14848 6016
rect 14912 5952 14928 6016
rect 14992 5952 15008 6016
rect 15072 5952 15088 6016
rect 15152 5952 15160 6016
rect 14840 5951 15160 5952
rect 24104 6016 24424 6017
rect 24104 5952 24112 6016
rect 24176 5952 24192 6016
rect 24256 5952 24272 6016
rect 24336 5952 24352 6016
rect 24416 5952 24424 6016
rect 24104 5951 24424 5952
rect 0 5448 800 5568
rect 28257 5538 28323 5541
rect 29200 5538 30000 5568
rect 28257 5536 30000 5538
rect 28257 5480 28262 5536
rect 28318 5480 30000 5536
rect 28257 5478 30000 5480
rect 28257 5475 28323 5478
rect 10208 5472 10528 5473
rect 10208 5408 10216 5472
rect 10280 5408 10296 5472
rect 10360 5408 10376 5472
rect 10440 5408 10456 5472
rect 10520 5408 10528 5472
rect 10208 5407 10528 5408
rect 19472 5472 19792 5473
rect 19472 5408 19480 5472
rect 19544 5408 19560 5472
rect 19624 5408 19640 5472
rect 19704 5408 19720 5472
rect 19784 5408 19792 5472
rect 29200 5448 30000 5478
rect 19472 5407 19792 5408
rect 5576 4928 5896 4929
rect 5576 4864 5584 4928
rect 5648 4864 5664 4928
rect 5728 4864 5744 4928
rect 5808 4864 5824 4928
rect 5888 4864 5896 4928
rect 5576 4863 5896 4864
rect 14840 4928 15160 4929
rect 14840 4864 14848 4928
rect 14912 4864 14928 4928
rect 14992 4864 15008 4928
rect 15072 4864 15088 4928
rect 15152 4864 15160 4928
rect 14840 4863 15160 4864
rect 24104 4928 24424 4929
rect 24104 4864 24112 4928
rect 24176 4864 24192 4928
rect 24256 4864 24272 4928
rect 24336 4864 24352 4928
rect 24416 4864 24424 4928
rect 24104 4863 24424 4864
rect 10208 4384 10528 4385
rect 10208 4320 10216 4384
rect 10280 4320 10296 4384
rect 10360 4320 10376 4384
rect 10440 4320 10456 4384
rect 10520 4320 10528 4384
rect 10208 4319 10528 4320
rect 19472 4384 19792 4385
rect 19472 4320 19480 4384
rect 19544 4320 19560 4384
rect 19624 4320 19640 4384
rect 19704 4320 19720 4384
rect 19784 4320 19792 4384
rect 19472 4319 19792 4320
rect 0 4178 800 4208
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4088 800 4118
rect 1393 4115 1459 4118
rect 28349 4178 28415 4181
rect 29200 4178 30000 4208
rect 28349 4176 30000 4178
rect 28349 4120 28354 4176
rect 28410 4120 30000 4176
rect 28349 4118 30000 4120
rect 28349 4115 28415 4118
rect 29200 4088 30000 4118
rect 5576 3840 5896 3841
rect 5576 3776 5584 3840
rect 5648 3776 5664 3840
rect 5728 3776 5744 3840
rect 5808 3776 5824 3840
rect 5888 3776 5896 3840
rect 5576 3775 5896 3776
rect 14840 3840 15160 3841
rect 14840 3776 14848 3840
rect 14912 3776 14928 3840
rect 14992 3776 15008 3840
rect 15072 3776 15088 3840
rect 15152 3776 15160 3840
rect 14840 3775 15160 3776
rect 24104 3840 24424 3841
rect 24104 3776 24112 3840
rect 24176 3776 24192 3840
rect 24256 3776 24272 3840
rect 24336 3776 24352 3840
rect 24416 3776 24424 3840
rect 24104 3775 24424 3776
rect 10208 3296 10528 3297
rect 10208 3232 10216 3296
rect 10280 3232 10296 3296
rect 10360 3232 10376 3296
rect 10440 3232 10456 3296
rect 10520 3232 10528 3296
rect 10208 3231 10528 3232
rect 19472 3296 19792 3297
rect 19472 3232 19480 3296
rect 19544 3232 19560 3296
rect 19624 3232 19640 3296
rect 19704 3232 19720 3296
rect 19784 3232 19792 3296
rect 19472 3231 19792 3232
rect 0 2818 800 2848
rect 1485 2818 1551 2821
rect 0 2816 1551 2818
rect 0 2760 1490 2816
rect 1546 2760 1551 2816
rect 0 2758 1551 2760
rect 0 2728 800 2758
rect 1485 2755 1551 2758
rect 28349 2818 28415 2821
rect 29200 2818 30000 2848
rect 28349 2816 30000 2818
rect 28349 2760 28354 2816
rect 28410 2760 30000 2816
rect 28349 2758 30000 2760
rect 28349 2755 28415 2758
rect 5576 2752 5896 2753
rect 5576 2688 5584 2752
rect 5648 2688 5664 2752
rect 5728 2688 5744 2752
rect 5808 2688 5824 2752
rect 5888 2688 5896 2752
rect 5576 2687 5896 2688
rect 14840 2752 15160 2753
rect 14840 2688 14848 2752
rect 14912 2688 14928 2752
rect 14992 2688 15008 2752
rect 15072 2688 15088 2752
rect 15152 2688 15160 2752
rect 14840 2687 15160 2688
rect 24104 2752 24424 2753
rect 24104 2688 24112 2752
rect 24176 2688 24192 2752
rect 24256 2688 24272 2752
rect 24336 2688 24352 2752
rect 24416 2688 24424 2752
rect 29200 2728 30000 2758
rect 24104 2687 24424 2688
rect 10208 2208 10528 2209
rect 10208 2144 10216 2208
rect 10280 2144 10296 2208
rect 10360 2144 10376 2208
rect 10440 2144 10456 2208
rect 10520 2144 10528 2208
rect 10208 2143 10528 2144
rect 19472 2208 19792 2209
rect 19472 2144 19480 2208
rect 19544 2144 19560 2208
rect 19624 2144 19640 2208
rect 19704 2144 19720 2208
rect 19784 2144 19792 2208
rect 19472 2143 19792 2144
rect 0 1458 800 1488
rect 1485 1458 1551 1461
rect 0 1456 1551 1458
rect 0 1400 1490 1456
rect 1546 1400 1551 1456
rect 0 1398 1551 1400
rect 0 1368 800 1398
rect 1485 1395 1551 1398
rect 29200 1368 30000 1488
rect 27521 98 27587 101
rect 29200 98 30000 128
rect 27521 96 30000 98
rect 27521 40 27526 96
rect 27582 40 30000 96
rect 27521 38 30000 40
rect 27521 35 27587 38
rect 29200 8 30000 38
<< via3 >>
rect 5584 27772 5648 27776
rect 5584 27716 5588 27772
rect 5588 27716 5644 27772
rect 5644 27716 5648 27772
rect 5584 27712 5648 27716
rect 5664 27772 5728 27776
rect 5664 27716 5668 27772
rect 5668 27716 5724 27772
rect 5724 27716 5728 27772
rect 5664 27712 5728 27716
rect 5744 27772 5808 27776
rect 5744 27716 5748 27772
rect 5748 27716 5804 27772
rect 5804 27716 5808 27772
rect 5744 27712 5808 27716
rect 5824 27772 5888 27776
rect 5824 27716 5828 27772
rect 5828 27716 5884 27772
rect 5884 27716 5888 27772
rect 5824 27712 5888 27716
rect 14848 27772 14912 27776
rect 14848 27716 14852 27772
rect 14852 27716 14908 27772
rect 14908 27716 14912 27772
rect 14848 27712 14912 27716
rect 14928 27772 14992 27776
rect 14928 27716 14932 27772
rect 14932 27716 14988 27772
rect 14988 27716 14992 27772
rect 14928 27712 14992 27716
rect 15008 27772 15072 27776
rect 15008 27716 15012 27772
rect 15012 27716 15068 27772
rect 15068 27716 15072 27772
rect 15008 27712 15072 27716
rect 15088 27772 15152 27776
rect 15088 27716 15092 27772
rect 15092 27716 15148 27772
rect 15148 27716 15152 27772
rect 15088 27712 15152 27716
rect 24112 27772 24176 27776
rect 24112 27716 24116 27772
rect 24116 27716 24172 27772
rect 24172 27716 24176 27772
rect 24112 27712 24176 27716
rect 24192 27772 24256 27776
rect 24192 27716 24196 27772
rect 24196 27716 24252 27772
rect 24252 27716 24256 27772
rect 24192 27712 24256 27716
rect 24272 27772 24336 27776
rect 24272 27716 24276 27772
rect 24276 27716 24332 27772
rect 24332 27716 24336 27772
rect 24272 27712 24336 27716
rect 24352 27772 24416 27776
rect 24352 27716 24356 27772
rect 24356 27716 24412 27772
rect 24412 27716 24416 27772
rect 24352 27712 24416 27716
rect 10216 27228 10280 27232
rect 10216 27172 10220 27228
rect 10220 27172 10276 27228
rect 10276 27172 10280 27228
rect 10216 27168 10280 27172
rect 10296 27228 10360 27232
rect 10296 27172 10300 27228
rect 10300 27172 10356 27228
rect 10356 27172 10360 27228
rect 10296 27168 10360 27172
rect 10376 27228 10440 27232
rect 10376 27172 10380 27228
rect 10380 27172 10436 27228
rect 10436 27172 10440 27228
rect 10376 27168 10440 27172
rect 10456 27228 10520 27232
rect 10456 27172 10460 27228
rect 10460 27172 10516 27228
rect 10516 27172 10520 27228
rect 10456 27168 10520 27172
rect 19480 27228 19544 27232
rect 19480 27172 19484 27228
rect 19484 27172 19540 27228
rect 19540 27172 19544 27228
rect 19480 27168 19544 27172
rect 19560 27228 19624 27232
rect 19560 27172 19564 27228
rect 19564 27172 19620 27228
rect 19620 27172 19624 27228
rect 19560 27168 19624 27172
rect 19640 27228 19704 27232
rect 19640 27172 19644 27228
rect 19644 27172 19700 27228
rect 19700 27172 19704 27228
rect 19640 27168 19704 27172
rect 19720 27228 19784 27232
rect 19720 27172 19724 27228
rect 19724 27172 19780 27228
rect 19780 27172 19784 27228
rect 19720 27168 19784 27172
rect 5584 26684 5648 26688
rect 5584 26628 5588 26684
rect 5588 26628 5644 26684
rect 5644 26628 5648 26684
rect 5584 26624 5648 26628
rect 5664 26684 5728 26688
rect 5664 26628 5668 26684
rect 5668 26628 5724 26684
rect 5724 26628 5728 26684
rect 5664 26624 5728 26628
rect 5744 26684 5808 26688
rect 5744 26628 5748 26684
rect 5748 26628 5804 26684
rect 5804 26628 5808 26684
rect 5744 26624 5808 26628
rect 5824 26684 5888 26688
rect 5824 26628 5828 26684
rect 5828 26628 5884 26684
rect 5884 26628 5888 26684
rect 5824 26624 5888 26628
rect 14848 26684 14912 26688
rect 14848 26628 14852 26684
rect 14852 26628 14908 26684
rect 14908 26628 14912 26684
rect 14848 26624 14912 26628
rect 14928 26684 14992 26688
rect 14928 26628 14932 26684
rect 14932 26628 14988 26684
rect 14988 26628 14992 26684
rect 14928 26624 14992 26628
rect 15008 26684 15072 26688
rect 15008 26628 15012 26684
rect 15012 26628 15068 26684
rect 15068 26628 15072 26684
rect 15008 26624 15072 26628
rect 15088 26684 15152 26688
rect 15088 26628 15092 26684
rect 15092 26628 15148 26684
rect 15148 26628 15152 26684
rect 15088 26624 15152 26628
rect 24112 26684 24176 26688
rect 24112 26628 24116 26684
rect 24116 26628 24172 26684
rect 24172 26628 24176 26684
rect 24112 26624 24176 26628
rect 24192 26684 24256 26688
rect 24192 26628 24196 26684
rect 24196 26628 24252 26684
rect 24252 26628 24256 26684
rect 24192 26624 24256 26628
rect 24272 26684 24336 26688
rect 24272 26628 24276 26684
rect 24276 26628 24332 26684
rect 24332 26628 24336 26684
rect 24272 26624 24336 26628
rect 24352 26684 24416 26688
rect 24352 26628 24356 26684
rect 24356 26628 24412 26684
rect 24412 26628 24416 26684
rect 24352 26624 24416 26628
rect 25636 26284 25700 26348
rect 10216 26140 10280 26144
rect 10216 26084 10220 26140
rect 10220 26084 10276 26140
rect 10276 26084 10280 26140
rect 10216 26080 10280 26084
rect 10296 26140 10360 26144
rect 10296 26084 10300 26140
rect 10300 26084 10356 26140
rect 10356 26084 10360 26140
rect 10296 26080 10360 26084
rect 10376 26140 10440 26144
rect 10376 26084 10380 26140
rect 10380 26084 10436 26140
rect 10436 26084 10440 26140
rect 10376 26080 10440 26084
rect 10456 26140 10520 26144
rect 10456 26084 10460 26140
rect 10460 26084 10516 26140
rect 10516 26084 10520 26140
rect 10456 26080 10520 26084
rect 19480 26140 19544 26144
rect 19480 26084 19484 26140
rect 19484 26084 19540 26140
rect 19540 26084 19544 26140
rect 19480 26080 19544 26084
rect 19560 26140 19624 26144
rect 19560 26084 19564 26140
rect 19564 26084 19620 26140
rect 19620 26084 19624 26140
rect 19560 26080 19624 26084
rect 19640 26140 19704 26144
rect 19640 26084 19644 26140
rect 19644 26084 19700 26140
rect 19700 26084 19704 26140
rect 19640 26080 19704 26084
rect 19720 26140 19784 26144
rect 19720 26084 19724 26140
rect 19724 26084 19780 26140
rect 19780 26084 19784 26140
rect 19720 26080 19784 26084
rect 5584 25596 5648 25600
rect 5584 25540 5588 25596
rect 5588 25540 5644 25596
rect 5644 25540 5648 25596
rect 5584 25536 5648 25540
rect 5664 25596 5728 25600
rect 5664 25540 5668 25596
rect 5668 25540 5724 25596
rect 5724 25540 5728 25596
rect 5664 25536 5728 25540
rect 5744 25596 5808 25600
rect 5744 25540 5748 25596
rect 5748 25540 5804 25596
rect 5804 25540 5808 25596
rect 5744 25536 5808 25540
rect 5824 25596 5888 25600
rect 5824 25540 5828 25596
rect 5828 25540 5884 25596
rect 5884 25540 5888 25596
rect 5824 25536 5888 25540
rect 14848 25596 14912 25600
rect 14848 25540 14852 25596
rect 14852 25540 14908 25596
rect 14908 25540 14912 25596
rect 14848 25536 14912 25540
rect 14928 25596 14992 25600
rect 14928 25540 14932 25596
rect 14932 25540 14988 25596
rect 14988 25540 14992 25596
rect 14928 25536 14992 25540
rect 15008 25596 15072 25600
rect 15008 25540 15012 25596
rect 15012 25540 15068 25596
rect 15068 25540 15072 25596
rect 15008 25536 15072 25540
rect 15088 25596 15152 25600
rect 15088 25540 15092 25596
rect 15092 25540 15148 25596
rect 15148 25540 15152 25596
rect 15088 25536 15152 25540
rect 24112 25596 24176 25600
rect 24112 25540 24116 25596
rect 24116 25540 24172 25596
rect 24172 25540 24176 25596
rect 24112 25536 24176 25540
rect 24192 25596 24256 25600
rect 24192 25540 24196 25596
rect 24196 25540 24252 25596
rect 24252 25540 24256 25596
rect 24192 25536 24256 25540
rect 24272 25596 24336 25600
rect 24272 25540 24276 25596
rect 24276 25540 24332 25596
rect 24332 25540 24336 25596
rect 24272 25536 24336 25540
rect 24352 25596 24416 25600
rect 24352 25540 24356 25596
rect 24356 25540 24412 25596
rect 24412 25540 24416 25596
rect 24352 25536 24416 25540
rect 10216 25052 10280 25056
rect 10216 24996 10220 25052
rect 10220 24996 10276 25052
rect 10276 24996 10280 25052
rect 10216 24992 10280 24996
rect 10296 25052 10360 25056
rect 10296 24996 10300 25052
rect 10300 24996 10356 25052
rect 10356 24996 10360 25052
rect 10296 24992 10360 24996
rect 10376 25052 10440 25056
rect 10376 24996 10380 25052
rect 10380 24996 10436 25052
rect 10436 24996 10440 25052
rect 10376 24992 10440 24996
rect 10456 25052 10520 25056
rect 10456 24996 10460 25052
rect 10460 24996 10516 25052
rect 10516 24996 10520 25052
rect 10456 24992 10520 24996
rect 19480 25052 19544 25056
rect 19480 24996 19484 25052
rect 19484 24996 19540 25052
rect 19540 24996 19544 25052
rect 19480 24992 19544 24996
rect 19560 25052 19624 25056
rect 19560 24996 19564 25052
rect 19564 24996 19620 25052
rect 19620 24996 19624 25052
rect 19560 24992 19624 24996
rect 19640 25052 19704 25056
rect 19640 24996 19644 25052
rect 19644 24996 19700 25052
rect 19700 24996 19704 25052
rect 19640 24992 19704 24996
rect 19720 25052 19784 25056
rect 19720 24996 19724 25052
rect 19724 24996 19780 25052
rect 19780 24996 19784 25052
rect 19720 24992 19784 24996
rect 16436 24924 16500 24988
rect 5584 24508 5648 24512
rect 5584 24452 5588 24508
rect 5588 24452 5644 24508
rect 5644 24452 5648 24508
rect 5584 24448 5648 24452
rect 5664 24508 5728 24512
rect 5664 24452 5668 24508
rect 5668 24452 5724 24508
rect 5724 24452 5728 24508
rect 5664 24448 5728 24452
rect 5744 24508 5808 24512
rect 5744 24452 5748 24508
rect 5748 24452 5804 24508
rect 5804 24452 5808 24508
rect 5744 24448 5808 24452
rect 5824 24508 5888 24512
rect 5824 24452 5828 24508
rect 5828 24452 5884 24508
rect 5884 24452 5888 24508
rect 5824 24448 5888 24452
rect 14848 24508 14912 24512
rect 14848 24452 14852 24508
rect 14852 24452 14908 24508
rect 14908 24452 14912 24508
rect 14848 24448 14912 24452
rect 14928 24508 14992 24512
rect 14928 24452 14932 24508
rect 14932 24452 14988 24508
rect 14988 24452 14992 24508
rect 14928 24448 14992 24452
rect 15008 24508 15072 24512
rect 15008 24452 15012 24508
rect 15012 24452 15068 24508
rect 15068 24452 15072 24508
rect 15008 24448 15072 24452
rect 15088 24508 15152 24512
rect 15088 24452 15092 24508
rect 15092 24452 15148 24508
rect 15148 24452 15152 24508
rect 15088 24448 15152 24452
rect 24112 24508 24176 24512
rect 24112 24452 24116 24508
rect 24116 24452 24172 24508
rect 24172 24452 24176 24508
rect 24112 24448 24176 24452
rect 24192 24508 24256 24512
rect 24192 24452 24196 24508
rect 24196 24452 24252 24508
rect 24252 24452 24256 24508
rect 24192 24448 24256 24452
rect 24272 24508 24336 24512
rect 24272 24452 24276 24508
rect 24276 24452 24332 24508
rect 24332 24452 24336 24508
rect 24272 24448 24336 24452
rect 24352 24508 24416 24512
rect 24352 24452 24356 24508
rect 24356 24452 24412 24508
rect 24412 24452 24416 24508
rect 24352 24448 24416 24452
rect 10216 23964 10280 23968
rect 10216 23908 10220 23964
rect 10220 23908 10276 23964
rect 10276 23908 10280 23964
rect 10216 23904 10280 23908
rect 10296 23964 10360 23968
rect 10296 23908 10300 23964
rect 10300 23908 10356 23964
rect 10356 23908 10360 23964
rect 10296 23904 10360 23908
rect 10376 23964 10440 23968
rect 10376 23908 10380 23964
rect 10380 23908 10436 23964
rect 10436 23908 10440 23964
rect 10376 23904 10440 23908
rect 10456 23964 10520 23968
rect 10456 23908 10460 23964
rect 10460 23908 10516 23964
rect 10516 23908 10520 23964
rect 10456 23904 10520 23908
rect 19480 23964 19544 23968
rect 19480 23908 19484 23964
rect 19484 23908 19540 23964
rect 19540 23908 19544 23964
rect 19480 23904 19544 23908
rect 19560 23964 19624 23968
rect 19560 23908 19564 23964
rect 19564 23908 19620 23964
rect 19620 23908 19624 23964
rect 19560 23904 19624 23908
rect 19640 23964 19704 23968
rect 19640 23908 19644 23964
rect 19644 23908 19700 23964
rect 19700 23908 19704 23964
rect 19640 23904 19704 23908
rect 19720 23964 19784 23968
rect 19720 23908 19724 23964
rect 19724 23908 19780 23964
rect 19780 23908 19784 23964
rect 19720 23904 19784 23908
rect 5584 23420 5648 23424
rect 5584 23364 5588 23420
rect 5588 23364 5644 23420
rect 5644 23364 5648 23420
rect 5584 23360 5648 23364
rect 5664 23420 5728 23424
rect 5664 23364 5668 23420
rect 5668 23364 5724 23420
rect 5724 23364 5728 23420
rect 5664 23360 5728 23364
rect 5744 23420 5808 23424
rect 5744 23364 5748 23420
rect 5748 23364 5804 23420
rect 5804 23364 5808 23420
rect 5744 23360 5808 23364
rect 5824 23420 5888 23424
rect 5824 23364 5828 23420
rect 5828 23364 5884 23420
rect 5884 23364 5888 23420
rect 5824 23360 5888 23364
rect 14848 23420 14912 23424
rect 14848 23364 14852 23420
rect 14852 23364 14908 23420
rect 14908 23364 14912 23420
rect 14848 23360 14912 23364
rect 14928 23420 14992 23424
rect 14928 23364 14932 23420
rect 14932 23364 14988 23420
rect 14988 23364 14992 23420
rect 14928 23360 14992 23364
rect 15008 23420 15072 23424
rect 15008 23364 15012 23420
rect 15012 23364 15068 23420
rect 15068 23364 15072 23420
rect 15008 23360 15072 23364
rect 15088 23420 15152 23424
rect 15088 23364 15092 23420
rect 15092 23364 15148 23420
rect 15148 23364 15152 23420
rect 15088 23360 15152 23364
rect 24112 23420 24176 23424
rect 24112 23364 24116 23420
rect 24116 23364 24172 23420
rect 24172 23364 24176 23420
rect 24112 23360 24176 23364
rect 24192 23420 24256 23424
rect 24192 23364 24196 23420
rect 24196 23364 24252 23420
rect 24252 23364 24256 23420
rect 24192 23360 24256 23364
rect 24272 23420 24336 23424
rect 24272 23364 24276 23420
rect 24276 23364 24332 23420
rect 24332 23364 24336 23420
rect 24272 23360 24336 23364
rect 24352 23420 24416 23424
rect 24352 23364 24356 23420
rect 24356 23364 24412 23420
rect 24412 23364 24416 23420
rect 24352 23360 24416 23364
rect 10216 22876 10280 22880
rect 10216 22820 10220 22876
rect 10220 22820 10276 22876
rect 10276 22820 10280 22876
rect 10216 22816 10280 22820
rect 10296 22876 10360 22880
rect 10296 22820 10300 22876
rect 10300 22820 10356 22876
rect 10356 22820 10360 22876
rect 10296 22816 10360 22820
rect 10376 22876 10440 22880
rect 10376 22820 10380 22876
rect 10380 22820 10436 22876
rect 10436 22820 10440 22876
rect 10376 22816 10440 22820
rect 10456 22876 10520 22880
rect 10456 22820 10460 22876
rect 10460 22820 10516 22876
rect 10516 22820 10520 22876
rect 10456 22816 10520 22820
rect 19480 22876 19544 22880
rect 19480 22820 19484 22876
rect 19484 22820 19540 22876
rect 19540 22820 19544 22876
rect 19480 22816 19544 22820
rect 19560 22876 19624 22880
rect 19560 22820 19564 22876
rect 19564 22820 19620 22876
rect 19620 22820 19624 22876
rect 19560 22816 19624 22820
rect 19640 22876 19704 22880
rect 19640 22820 19644 22876
rect 19644 22820 19700 22876
rect 19700 22820 19704 22876
rect 19640 22816 19704 22820
rect 19720 22876 19784 22880
rect 19720 22820 19724 22876
rect 19724 22820 19780 22876
rect 19780 22820 19784 22876
rect 19720 22816 19784 22820
rect 5584 22332 5648 22336
rect 5584 22276 5588 22332
rect 5588 22276 5644 22332
rect 5644 22276 5648 22332
rect 5584 22272 5648 22276
rect 5664 22332 5728 22336
rect 5664 22276 5668 22332
rect 5668 22276 5724 22332
rect 5724 22276 5728 22332
rect 5664 22272 5728 22276
rect 5744 22332 5808 22336
rect 5744 22276 5748 22332
rect 5748 22276 5804 22332
rect 5804 22276 5808 22332
rect 5744 22272 5808 22276
rect 5824 22332 5888 22336
rect 5824 22276 5828 22332
rect 5828 22276 5884 22332
rect 5884 22276 5888 22332
rect 5824 22272 5888 22276
rect 14848 22332 14912 22336
rect 14848 22276 14852 22332
rect 14852 22276 14908 22332
rect 14908 22276 14912 22332
rect 14848 22272 14912 22276
rect 14928 22332 14992 22336
rect 14928 22276 14932 22332
rect 14932 22276 14988 22332
rect 14988 22276 14992 22332
rect 14928 22272 14992 22276
rect 15008 22332 15072 22336
rect 15008 22276 15012 22332
rect 15012 22276 15068 22332
rect 15068 22276 15072 22332
rect 15008 22272 15072 22276
rect 15088 22332 15152 22336
rect 15088 22276 15092 22332
rect 15092 22276 15148 22332
rect 15148 22276 15152 22332
rect 15088 22272 15152 22276
rect 24112 22332 24176 22336
rect 24112 22276 24116 22332
rect 24116 22276 24172 22332
rect 24172 22276 24176 22332
rect 24112 22272 24176 22276
rect 24192 22332 24256 22336
rect 24192 22276 24196 22332
rect 24196 22276 24252 22332
rect 24252 22276 24256 22332
rect 24192 22272 24256 22276
rect 24272 22332 24336 22336
rect 24272 22276 24276 22332
rect 24276 22276 24332 22332
rect 24332 22276 24336 22332
rect 24272 22272 24336 22276
rect 24352 22332 24416 22336
rect 24352 22276 24356 22332
rect 24356 22276 24412 22332
rect 24412 22276 24416 22332
rect 24352 22272 24416 22276
rect 10216 21788 10280 21792
rect 10216 21732 10220 21788
rect 10220 21732 10276 21788
rect 10276 21732 10280 21788
rect 10216 21728 10280 21732
rect 10296 21788 10360 21792
rect 10296 21732 10300 21788
rect 10300 21732 10356 21788
rect 10356 21732 10360 21788
rect 10296 21728 10360 21732
rect 10376 21788 10440 21792
rect 10376 21732 10380 21788
rect 10380 21732 10436 21788
rect 10436 21732 10440 21788
rect 10376 21728 10440 21732
rect 10456 21788 10520 21792
rect 10456 21732 10460 21788
rect 10460 21732 10516 21788
rect 10516 21732 10520 21788
rect 10456 21728 10520 21732
rect 19480 21788 19544 21792
rect 19480 21732 19484 21788
rect 19484 21732 19540 21788
rect 19540 21732 19544 21788
rect 19480 21728 19544 21732
rect 19560 21788 19624 21792
rect 19560 21732 19564 21788
rect 19564 21732 19620 21788
rect 19620 21732 19624 21788
rect 19560 21728 19624 21732
rect 19640 21788 19704 21792
rect 19640 21732 19644 21788
rect 19644 21732 19700 21788
rect 19700 21732 19704 21788
rect 19640 21728 19704 21732
rect 19720 21788 19784 21792
rect 19720 21732 19724 21788
rect 19724 21732 19780 21788
rect 19780 21732 19784 21788
rect 19720 21728 19784 21732
rect 5584 21244 5648 21248
rect 5584 21188 5588 21244
rect 5588 21188 5644 21244
rect 5644 21188 5648 21244
rect 5584 21184 5648 21188
rect 5664 21244 5728 21248
rect 5664 21188 5668 21244
rect 5668 21188 5724 21244
rect 5724 21188 5728 21244
rect 5664 21184 5728 21188
rect 5744 21244 5808 21248
rect 5744 21188 5748 21244
rect 5748 21188 5804 21244
rect 5804 21188 5808 21244
rect 5744 21184 5808 21188
rect 5824 21244 5888 21248
rect 5824 21188 5828 21244
rect 5828 21188 5884 21244
rect 5884 21188 5888 21244
rect 5824 21184 5888 21188
rect 14848 21244 14912 21248
rect 14848 21188 14852 21244
rect 14852 21188 14908 21244
rect 14908 21188 14912 21244
rect 14848 21184 14912 21188
rect 14928 21244 14992 21248
rect 14928 21188 14932 21244
rect 14932 21188 14988 21244
rect 14988 21188 14992 21244
rect 14928 21184 14992 21188
rect 15008 21244 15072 21248
rect 15008 21188 15012 21244
rect 15012 21188 15068 21244
rect 15068 21188 15072 21244
rect 15008 21184 15072 21188
rect 15088 21244 15152 21248
rect 15088 21188 15092 21244
rect 15092 21188 15148 21244
rect 15148 21188 15152 21244
rect 15088 21184 15152 21188
rect 24112 21244 24176 21248
rect 24112 21188 24116 21244
rect 24116 21188 24172 21244
rect 24172 21188 24176 21244
rect 24112 21184 24176 21188
rect 24192 21244 24256 21248
rect 24192 21188 24196 21244
rect 24196 21188 24252 21244
rect 24252 21188 24256 21244
rect 24192 21184 24256 21188
rect 24272 21244 24336 21248
rect 24272 21188 24276 21244
rect 24276 21188 24332 21244
rect 24332 21188 24336 21244
rect 24272 21184 24336 21188
rect 24352 21244 24416 21248
rect 24352 21188 24356 21244
rect 24356 21188 24412 21244
rect 24412 21188 24416 21244
rect 24352 21184 24416 21188
rect 14596 20844 14660 20908
rect 10216 20700 10280 20704
rect 10216 20644 10220 20700
rect 10220 20644 10276 20700
rect 10276 20644 10280 20700
rect 10216 20640 10280 20644
rect 10296 20700 10360 20704
rect 10296 20644 10300 20700
rect 10300 20644 10356 20700
rect 10356 20644 10360 20700
rect 10296 20640 10360 20644
rect 10376 20700 10440 20704
rect 10376 20644 10380 20700
rect 10380 20644 10436 20700
rect 10436 20644 10440 20700
rect 10376 20640 10440 20644
rect 10456 20700 10520 20704
rect 10456 20644 10460 20700
rect 10460 20644 10516 20700
rect 10516 20644 10520 20700
rect 10456 20640 10520 20644
rect 19480 20700 19544 20704
rect 19480 20644 19484 20700
rect 19484 20644 19540 20700
rect 19540 20644 19544 20700
rect 19480 20640 19544 20644
rect 19560 20700 19624 20704
rect 19560 20644 19564 20700
rect 19564 20644 19620 20700
rect 19620 20644 19624 20700
rect 19560 20640 19624 20644
rect 19640 20700 19704 20704
rect 19640 20644 19644 20700
rect 19644 20644 19700 20700
rect 19700 20644 19704 20700
rect 19640 20640 19704 20644
rect 19720 20700 19784 20704
rect 19720 20644 19724 20700
rect 19724 20644 19780 20700
rect 19780 20644 19784 20700
rect 19720 20640 19784 20644
rect 5584 20156 5648 20160
rect 5584 20100 5588 20156
rect 5588 20100 5644 20156
rect 5644 20100 5648 20156
rect 5584 20096 5648 20100
rect 5664 20156 5728 20160
rect 5664 20100 5668 20156
rect 5668 20100 5724 20156
rect 5724 20100 5728 20156
rect 5664 20096 5728 20100
rect 5744 20156 5808 20160
rect 5744 20100 5748 20156
rect 5748 20100 5804 20156
rect 5804 20100 5808 20156
rect 5744 20096 5808 20100
rect 5824 20156 5888 20160
rect 5824 20100 5828 20156
rect 5828 20100 5884 20156
rect 5884 20100 5888 20156
rect 5824 20096 5888 20100
rect 14848 20156 14912 20160
rect 14848 20100 14852 20156
rect 14852 20100 14908 20156
rect 14908 20100 14912 20156
rect 14848 20096 14912 20100
rect 14928 20156 14992 20160
rect 14928 20100 14932 20156
rect 14932 20100 14988 20156
rect 14988 20100 14992 20156
rect 14928 20096 14992 20100
rect 15008 20156 15072 20160
rect 15008 20100 15012 20156
rect 15012 20100 15068 20156
rect 15068 20100 15072 20156
rect 15008 20096 15072 20100
rect 15088 20156 15152 20160
rect 15088 20100 15092 20156
rect 15092 20100 15148 20156
rect 15148 20100 15152 20156
rect 15088 20096 15152 20100
rect 24112 20156 24176 20160
rect 24112 20100 24116 20156
rect 24116 20100 24172 20156
rect 24172 20100 24176 20156
rect 24112 20096 24176 20100
rect 24192 20156 24256 20160
rect 24192 20100 24196 20156
rect 24196 20100 24252 20156
rect 24252 20100 24256 20156
rect 24192 20096 24256 20100
rect 24272 20156 24336 20160
rect 24272 20100 24276 20156
rect 24276 20100 24332 20156
rect 24332 20100 24336 20156
rect 24272 20096 24336 20100
rect 24352 20156 24416 20160
rect 24352 20100 24356 20156
rect 24356 20100 24412 20156
rect 24412 20100 24416 20156
rect 24352 20096 24416 20100
rect 10216 19612 10280 19616
rect 10216 19556 10220 19612
rect 10220 19556 10276 19612
rect 10276 19556 10280 19612
rect 10216 19552 10280 19556
rect 10296 19612 10360 19616
rect 10296 19556 10300 19612
rect 10300 19556 10356 19612
rect 10356 19556 10360 19612
rect 10296 19552 10360 19556
rect 10376 19612 10440 19616
rect 10376 19556 10380 19612
rect 10380 19556 10436 19612
rect 10436 19556 10440 19612
rect 10376 19552 10440 19556
rect 10456 19612 10520 19616
rect 10456 19556 10460 19612
rect 10460 19556 10516 19612
rect 10516 19556 10520 19612
rect 10456 19552 10520 19556
rect 19480 19612 19544 19616
rect 19480 19556 19484 19612
rect 19484 19556 19540 19612
rect 19540 19556 19544 19612
rect 19480 19552 19544 19556
rect 19560 19612 19624 19616
rect 19560 19556 19564 19612
rect 19564 19556 19620 19612
rect 19620 19556 19624 19612
rect 19560 19552 19624 19556
rect 19640 19612 19704 19616
rect 19640 19556 19644 19612
rect 19644 19556 19700 19612
rect 19700 19556 19704 19612
rect 19640 19552 19704 19556
rect 19720 19612 19784 19616
rect 19720 19556 19724 19612
rect 19724 19556 19780 19612
rect 19780 19556 19784 19612
rect 19720 19552 19784 19556
rect 5584 19068 5648 19072
rect 5584 19012 5588 19068
rect 5588 19012 5644 19068
rect 5644 19012 5648 19068
rect 5584 19008 5648 19012
rect 5664 19068 5728 19072
rect 5664 19012 5668 19068
rect 5668 19012 5724 19068
rect 5724 19012 5728 19068
rect 5664 19008 5728 19012
rect 5744 19068 5808 19072
rect 5744 19012 5748 19068
rect 5748 19012 5804 19068
rect 5804 19012 5808 19068
rect 5744 19008 5808 19012
rect 5824 19068 5888 19072
rect 5824 19012 5828 19068
rect 5828 19012 5884 19068
rect 5884 19012 5888 19068
rect 5824 19008 5888 19012
rect 14848 19068 14912 19072
rect 14848 19012 14852 19068
rect 14852 19012 14908 19068
rect 14908 19012 14912 19068
rect 14848 19008 14912 19012
rect 14928 19068 14992 19072
rect 14928 19012 14932 19068
rect 14932 19012 14988 19068
rect 14988 19012 14992 19068
rect 14928 19008 14992 19012
rect 15008 19068 15072 19072
rect 15008 19012 15012 19068
rect 15012 19012 15068 19068
rect 15068 19012 15072 19068
rect 15008 19008 15072 19012
rect 15088 19068 15152 19072
rect 15088 19012 15092 19068
rect 15092 19012 15148 19068
rect 15148 19012 15152 19068
rect 15088 19008 15152 19012
rect 24112 19068 24176 19072
rect 24112 19012 24116 19068
rect 24116 19012 24172 19068
rect 24172 19012 24176 19068
rect 24112 19008 24176 19012
rect 24192 19068 24256 19072
rect 24192 19012 24196 19068
rect 24196 19012 24252 19068
rect 24252 19012 24256 19068
rect 24192 19008 24256 19012
rect 24272 19068 24336 19072
rect 24272 19012 24276 19068
rect 24276 19012 24332 19068
rect 24332 19012 24336 19068
rect 24272 19008 24336 19012
rect 24352 19068 24416 19072
rect 24352 19012 24356 19068
rect 24356 19012 24412 19068
rect 24412 19012 24416 19068
rect 24352 19008 24416 19012
rect 10216 18524 10280 18528
rect 10216 18468 10220 18524
rect 10220 18468 10276 18524
rect 10276 18468 10280 18524
rect 10216 18464 10280 18468
rect 10296 18524 10360 18528
rect 10296 18468 10300 18524
rect 10300 18468 10356 18524
rect 10356 18468 10360 18524
rect 10296 18464 10360 18468
rect 10376 18524 10440 18528
rect 10376 18468 10380 18524
rect 10380 18468 10436 18524
rect 10436 18468 10440 18524
rect 10376 18464 10440 18468
rect 10456 18524 10520 18528
rect 10456 18468 10460 18524
rect 10460 18468 10516 18524
rect 10516 18468 10520 18524
rect 10456 18464 10520 18468
rect 19480 18524 19544 18528
rect 19480 18468 19484 18524
rect 19484 18468 19540 18524
rect 19540 18468 19544 18524
rect 19480 18464 19544 18468
rect 19560 18524 19624 18528
rect 19560 18468 19564 18524
rect 19564 18468 19620 18524
rect 19620 18468 19624 18524
rect 19560 18464 19624 18468
rect 19640 18524 19704 18528
rect 19640 18468 19644 18524
rect 19644 18468 19700 18524
rect 19700 18468 19704 18524
rect 19640 18464 19704 18468
rect 19720 18524 19784 18528
rect 19720 18468 19724 18524
rect 19724 18468 19780 18524
rect 19780 18468 19784 18524
rect 19720 18464 19784 18468
rect 16436 18396 16500 18460
rect 5584 17980 5648 17984
rect 5584 17924 5588 17980
rect 5588 17924 5644 17980
rect 5644 17924 5648 17980
rect 5584 17920 5648 17924
rect 5664 17980 5728 17984
rect 5664 17924 5668 17980
rect 5668 17924 5724 17980
rect 5724 17924 5728 17980
rect 5664 17920 5728 17924
rect 5744 17980 5808 17984
rect 5744 17924 5748 17980
rect 5748 17924 5804 17980
rect 5804 17924 5808 17980
rect 5744 17920 5808 17924
rect 5824 17980 5888 17984
rect 5824 17924 5828 17980
rect 5828 17924 5884 17980
rect 5884 17924 5888 17980
rect 5824 17920 5888 17924
rect 14848 17980 14912 17984
rect 14848 17924 14852 17980
rect 14852 17924 14908 17980
rect 14908 17924 14912 17980
rect 14848 17920 14912 17924
rect 14928 17980 14992 17984
rect 14928 17924 14932 17980
rect 14932 17924 14988 17980
rect 14988 17924 14992 17980
rect 14928 17920 14992 17924
rect 15008 17980 15072 17984
rect 15008 17924 15012 17980
rect 15012 17924 15068 17980
rect 15068 17924 15072 17980
rect 15008 17920 15072 17924
rect 15088 17980 15152 17984
rect 15088 17924 15092 17980
rect 15092 17924 15148 17980
rect 15148 17924 15152 17980
rect 15088 17920 15152 17924
rect 24112 17980 24176 17984
rect 24112 17924 24116 17980
rect 24116 17924 24172 17980
rect 24172 17924 24176 17980
rect 24112 17920 24176 17924
rect 24192 17980 24256 17984
rect 24192 17924 24196 17980
rect 24196 17924 24252 17980
rect 24252 17924 24256 17980
rect 24192 17920 24256 17924
rect 24272 17980 24336 17984
rect 24272 17924 24276 17980
rect 24276 17924 24332 17980
rect 24332 17924 24336 17980
rect 24272 17920 24336 17924
rect 24352 17980 24416 17984
rect 24352 17924 24356 17980
rect 24356 17924 24412 17980
rect 24412 17924 24416 17980
rect 24352 17920 24416 17924
rect 25636 17716 25700 17780
rect 10216 17436 10280 17440
rect 10216 17380 10220 17436
rect 10220 17380 10276 17436
rect 10276 17380 10280 17436
rect 10216 17376 10280 17380
rect 10296 17436 10360 17440
rect 10296 17380 10300 17436
rect 10300 17380 10356 17436
rect 10356 17380 10360 17436
rect 10296 17376 10360 17380
rect 10376 17436 10440 17440
rect 10376 17380 10380 17436
rect 10380 17380 10436 17436
rect 10436 17380 10440 17436
rect 10376 17376 10440 17380
rect 10456 17436 10520 17440
rect 10456 17380 10460 17436
rect 10460 17380 10516 17436
rect 10516 17380 10520 17436
rect 10456 17376 10520 17380
rect 19480 17436 19544 17440
rect 19480 17380 19484 17436
rect 19484 17380 19540 17436
rect 19540 17380 19544 17436
rect 19480 17376 19544 17380
rect 19560 17436 19624 17440
rect 19560 17380 19564 17436
rect 19564 17380 19620 17436
rect 19620 17380 19624 17436
rect 19560 17376 19624 17380
rect 19640 17436 19704 17440
rect 19640 17380 19644 17436
rect 19644 17380 19700 17436
rect 19700 17380 19704 17436
rect 19640 17376 19704 17380
rect 19720 17436 19784 17440
rect 19720 17380 19724 17436
rect 19724 17380 19780 17436
rect 19780 17380 19784 17436
rect 19720 17376 19784 17380
rect 5584 16892 5648 16896
rect 5584 16836 5588 16892
rect 5588 16836 5644 16892
rect 5644 16836 5648 16892
rect 5584 16832 5648 16836
rect 5664 16892 5728 16896
rect 5664 16836 5668 16892
rect 5668 16836 5724 16892
rect 5724 16836 5728 16892
rect 5664 16832 5728 16836
rect 5744 16892 5808 16896
rect 5744 16836 5748 16892
rect 5748 16836 5804 16892
rect 5804 16836 5808 16892
rect 5744 16832 5808 16836
rect 5824 16892 5888 16896
rect 5824 16836 5828 16892
rect 5828 16836 5884 16892
rect 5884 16836 5888 16892
rect 5824 16832 5888 16836
rect 14848 16892 14912 16896
rect 14848 16836 14852 16892
rect 14852 16836 14908 16892
rect 14908 16836 14912 16892
rect 14848 16832 14912 16836
rect 14928 16892 14992 16896
rect 14928 16836 14932 16892
rect 14932 16836 14988 16892
rect 14988 16836 14992 16892
rect 14928 16832 14992 16836
rect 15008 16892 15072 16896
rect 15008 16836 15012 16892
rect 15012 16836 15068 16892
rect 15068 16836 15072 16892
rect 15008 16832 15072 16836
rect 15088 16892 15152 16896
rect 15088 16836 15092 16892
rect 15092 16836 15148 16892
rect 15148 16836 15152 16892
rect 15088 16832 15152 16836
rect 24112 16892 24176 16896
rect 24112 16836 24116 16892
rect 24116 16836 24172 16892
rect 24172 16836 24176 16892
rect 24112 16832 24176 16836
rect 24192 16892 24256 16896
rect 24192 16836 24196 16892
rect 24196 16836 24252 16892
rect 24252 16836 24256 16892
rect 24192 16832 24256 16836
rect 24272 16892 24336 16896
rect 24272 16836 24276 16892
rect 24276 16836 24332 16892
rect 24332 16836 24336 16892
rect 24272 16832 24336 16836
rect 24352 16892 24416 16896
rect 24352 16836 24356 16892
rect 24356 16836 24412 16892
rect 24412 16836 24416 16892
rect 24352 16832 24416 16836
rect 13860 16628 13924 16692
rect 10216 16348 10280 16352
rect 10216 16292 10220 16348
rect 10220 16292 10276 16348
rect 10276 16292 10280 16348
rect 10216 16288 10280 16292
rect 10296 16348 10360 16352
rect 10296 16292 10300 16348
rect 10300 16292 10356 16348
rect 10356 16292 10360 16348
rect 10296 16288 10360 16292
rect 10376 16348 10440 16352
rect 10376 16292 10380 16348
rect 10380 16292 10436 16348
rect 10436 16292 10440 16348
rect 10376 16288 10440 16292
rect 10456 16348 10520 16352
rect 10456 16292 10460 16348
rect 10460 16292 10516 16348
rect 10516 16292 10520 16348
rect 10456 16288 10520 16292
rect 19480 16348 19544 16352
rect 19480 16292 19484 16348
rect 19484 16292 19540 16348
rect 19540 16292 19544 16348
rect 19480 16288 19544 16292
rect 19560 16348 19624 16352
rect 19560 16292 19564 16348
rect 19564 16292 19620 16348
rect 19620 16292 19624 16348
rect 19560 16288 19624 16292
rect 19640 16348 19704 16352
rect 19640 16292 19644 16348
rect 19644 16292 19700 16348
rect 19700 16292 19704 16348
rect 19640 16288 19704 16292
rect 19720 16348 19784 16352
rect 19720 16292 19724 16348
rect 19724 16292 19780 16348
rect 19780 16292 19784 16348
rect 19720 16288 19784 16292
rect 5584 15804 5648 15808
rect 5584 15748 5588 15804
rect 5588 15748 5644 15804
rect 5644 15748 5648 15804
rect 5584 15744 5648 15748
rect 5664 15804 5728 15808
rect 5664 15748 5668 15804
rect 5668 15748 5724 15804
rect 5724 15748 5728 15804
rect 5664 15744 5728 15748
rect 5744 15804 5808 15808
rect 5744 15748 5748 15804
rect 5748 15748 5804 15804
rect 5804 15748 5808 15804
rect 5744 15744 5808 15748
rect 5824 15804 5888 15808
rect 5824 15748 5828 15804
rect 5828 15748 5884 15804
rect 5884 15748 5888 15804
rect 5824 15744 5888 15748
rect 14848 15804 14912 15808
rect 14848 15748 14852 15804
rect 14852 15748 14908 15804
rect 14908 15748 14912 15804
rect 14848 15744 14912 15748
rect 14928 15804 14992 15808
rect 14928 15748 14932 15804
rect 14932 15748 14988 15804
rect 14988 15748 14992 15804
rect 14928 15744 14992 15748
rect 15008 15804 15072 15808
rect 15008 15748 15012 15804
rect 15012 15748 15068 15804
rect 15068 15748 15072 15804
rect 15008 15744 15072 15748
rect 15088 15804 15152 15808
rect 15088 15748 15092 15804
rect 15092 15748 15148 15804
rect 15148 15748 15152 15804
rect 15088 15744 15152 15748
rect 24112 15804 24176 15808
rect 24112 15748 24116 15804
rect 24116 15748 24172 15804
rect 24172 15748 24176 15804
rect 24112 15744 24176 15748
rect 24192 15804 24256 15808
rect 24192 15748 24196 15804
rect 24196 15748 24252 15804
rect 24252 15748 24256 15804
rect 24192 15744 24256 15748
rect 24272 15804 24336 15808
rect 24272 15748 24276 15804
rect 24276 15748 24332 15804
rect 24332 15748 24336 15804
rect 24272 15744 24336 15748
rect 24352 15804 24416 15808
rect 24352 15748 24356 15804
rect 24356 15748 24412 15804
rect 24412 15748 24416 15804
rect 24352 15744 24416 15748
rect 19932 15404 19996 15468
rect 13492 15268 13556 15332
rect 10216 15260 10280 15264
rect 10216 15204 10220 15260
rect 10220 15204 10276 15260
rect 10276 15204 10280 15260
rect 10216 15200 10280 15204
rect 10296 15260 10360 15264
rect 10296 15204 10300 15260
rect 10300 15204 10356 15260
rect 10356 15204 10360 15260
rect 10296 15200 10360 15204
rect 10376 15260 10440 15264
rect 10376 15204 10380 15260
rect 10380 15204 10436 15260
rect 10436 15204 10440 15260
rect 10376 15200 10440 15204
rect 10456 15260 10520 15264
rect 10456 15204 10460 15260
rect 10460 15204 10516 15260
rect 10516 15204 10520 15260
rect 10456 15200 10520 15204
rect 19480 15260 19544 15264
rect 19480 15204 19484 15260
rect 19484 15204 19540 15260
rect 19540 15204 19544 15260
rect 19480 15200 19544 15204
rect 19560 15260 19624 15264
rect 19560 15204 19564 15260
rect 19564 15204 19620 15260
rect 19620 15204 19624 15260
rect 19560 15200 19624 15204
rect 19640 15260 19704 15264
rect 19640 15204 19644 15260
rect 19644 15204 19700 15260
rect 19700 15204 19704 15260
rect 19640 15200 19704 15204
rect 19720 15260 19784 15264
rect 19720 15204 19724 15260
rect 19724 15204 19780 15260
rect 19780 15204 19784 15260
rect 19720 15200 19784 15204
rect 13860 14996 13924 15060
rect 5584 14716 5648 14720
rect 5584 14660 5588 14716
rect 5588 14660 5644 14716
rect 5644 14660 5648 14716
rect 5584 14656 5648 14660
rect 5664 14716 5728 14720
rect 5664 14660 5668 14716
rect 5668 14660 5724 14716
rect 5724 14660 5728 14716
rect 5664 14656 5728 14660
rect 5744 14716 5808 14720
rect 5744 14660 5748 14716
rect 5748 14660 5804 14716
rect 5804 14660 5808 14716
rect 5744 14656 5808 14660
rect 5824 14716 5888 14720
rect 5824 14660 5828 14716
rect 5828 14660 5884 14716
rect 5884 14660 5888 14716
rect 5824 14656 5888 14660
rect 14848 14716 14912 14720
rect 14848 14660 14852 14716
rect 14852 14660 14908 14716
rect 14908 14660 14912 14716
rect 14848 14656 14912 14660
rect 14928 14716 14992 14720
rect 14928 14660 14932 14716
rect 14932 14660 14988 14716
rect 14988 14660 14992 14716
rect 14928 14656 14992 14660
rect 15008 14716 15072 14720
rect 15008 14660 15012 14716
rect 15012 14660 15068 14716
rect 15068 14660 15072 14716
rect 15008 14656 15072 14660
rect 15088 14716 15152 14720
rect 15088 14660 15092 14716
rect 15092 14660 15148 14716
rect 15148 14660 15152 14716
rect 15088 14656 15152 14660
rect 24112 14716 24176 14720
rect 24112 14660 24116 14716
rect 24116 14660 24172 14716
rect 24172 14660 24176 14716
rect 24112 14656 24176 14660
rect 24192 14716 24256 14720
rect 24192 14660 24196 14716
rect 24196 14660 24252 14716
rect 24252 14660 24256 14716
rect 24192 14656 24256 14660
rect 24272 14716 24336 14720
rect 24272 14660 24276 14716
rect 24276 14660 24332 14716
rect 24332 14660 24336 14716
rect 24272 14656 24336 14660
rect 24352 14716 24416 14720
rect 24352 14660 24356 14716
rect 24356 14660 24412 14716
rect 24412 14660 24416 14716
rect 24352 14656 24416 14660
rect 10216 14172 10280 14176
rect 10216 14116 10220 14172
rect 10220 14116 10276 14172
rect 10276 14116 10280 14172
rect 10216 14112 10280 14116
rect 10296 14172 10360 14176
rect 10296 14116 10300 14172
rect 10300 14116 10356 14172
rect 10356 14116 10360 14172
rect 10296 14112 10360 14116
rect 10376 14172 10440 14176
rect 10376 14116 10380 14172
rect 10380 14116 10436 14172
rect 10436 14116 10440 14172
rect 10376 14112 10440 14116
rect 10456 14172 10520 14176
rect 10456 14116 10460 14172
rect 10460 14116 10516 14172
rect 10516 14116 10520 14172
rect 10456 14112 10520 14116
rect 19480 14172 19544 14176
rect 19480 14116 19484 14172
rect 19484 14116 19540 14172
rect 19540 14116 19544 14172
rect 19480 14112 19544 14116
rect 19560 14172 19624 14176
rect 19560 14116 19564 14172
rect 19564 14116 19620 14172
rect 19620 14116 19624 14172
rect 19560 14112 19624 14116
rect 19640 14172 19704 14176
rect 19640 14116 19644 14172
rect 19644 14116 19700 14172
rect 19700 14116 19704 14172
rect 19640 14112 19704 14116
rect 19720 14172 19784 14176
rect 19720 14116 19724 14172
rect 19724 14116 19780 14172
rect 19780 14116 19784 14172
rect 19720 14112 19784 14116
rect 5584 13628 5648 13632
rect 5584 13572 5588 13628
rect 5588 13572 5644 13628
rect 5644 13572 5648 13628
rect 5584 13568 5648 13572
rect 5664 13628 5728 13632
rect 5664 13572 5668 13628
rect 5668 13572 5724 13628
rect 5724 13572 5728 13628
rect 5664 13568 5728 13572
rect 5744 13628 5808 13632
rect 5744 13572 5748 13628
rect 5748 13572 5804 13628
rect 5804 13572 5808 13628
rect 5744 13568 5808 13572
rect 5824 13628 5888 13632
rect 5824 13572 5828 13628
rect 5828 13572 5884 13628
rect 5884 13572 5888 13628
rect 5824 13568 5888 13572
rect 14848 13628 14912 13632
rect 14848 13572 14852 13628
rect 14852 13572 14908 13628
rect 14908 13572 14912 13628
rect 14848 13568 14912 13572
rect 14928 13628 14992 13632
rect 14928 13572 14932 13628
rect 14932 13572 14988 13628
rect 14988 13572 14992 13628
rect 14928 13568 14992 13572
rect 15008 13628 15072 13632
rect 15008 13572 15012 13628
rect 15012 13572 15068 13628
rect 15068 13572 15072 13628
rect 15008 13568 15072 13572
rect 15088 13628 15152 13632
rect 15088 13572 15092 13628
rect 15092 13572 15148 13628
rect 15148 13572 15152 13628
rect 15088 13568 15152 13572
rect 24112 13628 24176 13632
rect 24112 13572 24116 13628
rect 24116 13572 24172 13628
rect 24172 13572 24176 13628
rect 24112 13568 24176 13572
rect 24192 13628 24256 13632
rect 24192 13572 24196 13628
rect 24196 13572 24252 13628
rect 24252 13572 24256 13628
rect 24192 13568 24256 13572
rect 24272 13628 24336 13632
rect 24272 13572 24276 13628
rect 24276 13572 24332 13628
rect 24332 13572 24336 13628
rect 24272 13568 24336 13572
rect 24352 13628 24416 13632
rect 24352 13572 24356 13628
rect 24356 13572 24412 13628
rect 24412 13572 24416 13628
rect 24352 13568 24416 13572
rect 10216 13084 10280 13088
rect 10216 13028 10220 13084
rect 10220 13028 10276 13084
rect 10276 13028 10280 13084
rect 10216 13024 10280 13028
rect 10296 13084 10360 13088
rect 10296 13028 10300 13084
rect 10300 13028 10356 13084
rect 10356 13028 10360 13084
rect 10296 13024 10360 13028
rect 10376 13084 10440 13088
rect 10376 13028 10380 13084
rect 10380 13028 10436 13084
rect 10436 13028 10440 13084
rect 10376 13024 10440 13028
rect 10456 13084 10520 13088
rect 10456 13028 10460 13084
rect 10460 13028 10516 13084
rect 10516 13028 10520 13084
rect 10456 13024 10520 13028
rect 19480 13084 19544 13088
rect 19480 13028 19484 13084
rect 19484 13028 19540 13084
rect 19540 13028 19544 13084
rect 19480 13024 19544 13028
rect 19560 13084 19624 13088
rect 19560 13028 19564 13084
rect 19564 13028 19620 13084
rect 19620 13028 19624 13084
rect 19560 13024 19624 13028
rect 19640 13084 19704 13088
rect 19640 13028 19644 13084
rect 19644 13028 19700 13084
rect 19700 13028 19704 13084
rect 19640 13024 19704 13028
rect 19720 13084 19784 13088
rect 19720 13028 19724 13084
rect 19724 13028 19780 13084
rect 19780 13028 19784 13084
rect 19720 13024 19784 13028
rect 5584 12540 5648 12544
rect 5584 12484 5588 12540
rect 5588 12484 5644 12540
rect 5644 12484 5648 12540
rect 5584 12480 5648 12484
rect 5664 12540 5728 12544
rect 5664 12484 5668 12540
rect 5668 12484 5724 12540
rect 5724 12484 5728 12540
rect 5664 12480 5728 12484
rect 5744 12540 5808 12544
rect 5744 12484 5748 12540
rect 5748 12484 5804 12540
rect 5804 12484 5808 12540
rect 5744 12480 5808 12484
rect 5824 12540 5888 12544
rect 5824 12484 5828 12540
rect 5828 12484 5884 12540
rect 5884 12484 5888 12540
rect 5824 12480 5888 12484
rect 14848 12540 14912 12544
rect 14848 12484 14852 12540
rect 14852 12484 14908 12540
rect 14908 12484 14912 12540
rect 14848 12480 14912 12484
rect 14928 12540 14992 12544
rect 14928 12484 14932 12540
rect 14932 12484 14988 12540
rect 14988 12484 14992 12540
rect 14928 12480 14992 12484
rect 15008 12540 15072 12544
rect 15008 12484 15012 12540
rect 15012 12484 15068 12540
rect 15068 12484 15072 12540
rect 15008 12480 15072 12484
rect 15088 12540 15152 12544
rect 15088 12484 15092 12540
rect 15092 12484 15148 12540
rect 15148 12484 15152 12540
rect 15088 12480 15152 12484
rect 24112 12540 24176 12544
rect 24112 12484 24116 12540
rect 24116 12484 24172 12540
rect 24172 12484 24176 12540
rect 24112 12480 24176 12484
rect 24192 12540 24256 12544
rect 24192 12484 24196 12540
rect 24196 12484 24252 12540
rect 24252 12484 24256 12540
rect 24192 12480 24256 12484
rect 24272 12540 24336 12544
rect 24272 12484 24276 12540
rect 24276 12484 24332 12540
rect 24332 12484 24336 12540
rect 24272 12480 24336 12484
rect 24352 12540 24416 12544
rect 24352 12484 24356 12540
rect 24356 12484 24412 12540
rect 24412 12484 24416 12540
rect 24352 12480 24416 12484
rect 13676 12004 13740 12068
rect 14596 12004 14660 12068
rect 10216 11996 10280 12000
rect 10216 11940 10220 11996
rect 10220 11940 10276 11996
rect 10276 11940 10280 11996
rect 10216 11936 10280 11940
rect 10296 11996 10360 12000
rect 10296 11940 10300 11996
rect 10300 11940 10356 11996
rect 10356 11940 10360 11996
rect 10296 11936 10360 11940
rect 10376 11996 10440 12000
rect 10376 11940 10380 11996
rect 10380 11940 10436 11996
rect 10436 11940 10440 11996
rect 10376 11936 10440 11940
rect 10456 11996 10520 12000
rect 10456 11940 10460 11996
rect 10460 11940 10516 11996
rect 10516 11940 10520 11996
rect 10456 11936 10520 11940
rect 19480 11996 19544 12000
rect 19480 11940 19484 11996
rect 19484 11940 19540 11996
rect 19540 11940 19544 11996
rect 19480 11936 19544 11940
rect 19560 11996 19624 12000
rect 19560 11940 19564 11996
rect 19564 11940 19620 11996
rect 19620 11940 19624 11996
rect 19560 11936 19624 11940
rect 19640 11996 19704 12000
rect 19640 11940 19644 11996
rect 19644 11940 19700 11996
rect 19700 11940 19704 11996
rect 19640 11936 19704 11940
rect 19720 11996 19784 12000
rect 19720 11940 19724 11996
rect 19724 11940 19780 11996
rect 19780 11940 19784 11996
rect 19720 11936 19784 11940
rect 5584 11452 5648 11456
rect 5584 11396 5588 11452
rect 5588 11396 5644 11452
rect 5644 11396 5648 11452
rect 5584 11392 5648 11396
rect 5664 11452 5728 11456
rect 5664 11396 5668 11452
rect 5668 11396 5724 11452
rect 5724 11396 5728 11452
rect 5664 11392 5728 11396
rect 5744 11452 5808 11456
rect 5744 11396 5748 11452
rect 5748 11396 5804 11452
rect 5804 11396 5808 11452
rect 5744 11392 5808 11396
rect 5824 11452 5888 11456
rect 5824 11396 5828 11452
rect 5828 11396 5884 11452
rect 5884 11396 5888 11452
rect 5824 11392 5888 11396
rect 14848 11452 14912 11456
rect 14848 11396 14852 11452
rect 14852 11396 14908 11452
rect 14908 11396 14912 11452
rect 14848 11392 14912 11396
rect 14928 11452 14992 11456
rect 14928 11396 14932 11452
rect 14932 11396 14988 11452
rect 14988 11396 14992 11452
rect 14928 11392 14992 11396
rect 15008 11452 15072 11456
rect 15008 11396 15012 11452
rect 15012 11396 15068 11452
rect 15068 11396 15072 11452
rect 15008 11392 15072 11396
rect 15088 11452 15152 11456
rect 15088 11396 15092 11452
rect 15092 11396 15148 11452
rect 15148 11396 15152 11452
rect 15088 11392 15152 11396
rect 24112 11452 24176 11456
rect 24112 11396 24116 11452
rect 24116 11396 24172 11452
rect 24172 11396 24176 11452
rect 24112 11392 24176 11396
rect 24192 11452 24256 11456
rect 24192 11396 24196 11452
rect 24196 11396 24252 11452
rect 24252 11396 24256 11452
rect 24192 11392 24256 11396
rect 24272 11452 24336 11456
rect 24272 11396 24276 11452
rect 24276 11396 24332 11452
rect 24332 11396 24336 11452
rect 24272 11392 24336 11396
rect 24352 11452 24416 11456
rect 24352 11396 24356 11452
rect 24356 11396 24412 11452
rect 24412 11396 24416 11452
rect 24352 11392 24416 11396
rect 10216 10908 10280 10912
rect 10216 10852 10220 10908
rect 10220 10852 10276 10908
rect 10276 10852 10280 10908
rect 10216 10848 10280 10852
rect 10296 10908 10360 10912
rect 10296 10852 10300 10908
rect 10300 10852 10356 10908
rect 10356 10852 10360 10908
rect 10296 10848 10360 10852
rect 10376 10908 10440 10912
rect 10376 10852 10380 10908
rect 10380 10852 10436 10908
rect 10436 10852 10440 10908
rect 10376 10848 10440 10852
rect 10456 10908 10520 10912
rect 10456 10852 10460 10908
rect 10460 10852 10516 10908
rect 10516 10852 10520 10908
rect 10456 10848 10520 10852
rect 19480 10908 19544 10912
rect 19480 10852 19484 10908
rect 19484 10852 19540 10908
rect 19540 10852 19544 10908
rect 19480 10848 19544 10852
rect 19560 10908 19624 10912
rect 19560 10852 19564 10908
rect 19564 10852 19620 10908
rect 19620 10852 19624 10908
rect 19560 10848 19624 10852
rect 19640 10908 19704 10912
rect 19640 10852 19644 10908
rect 19644 10852 19700 10908
rect 19700 10852 19704 10908
rect 19640 10848 19704 10852
rect 19720 10908 19784 10912
rect 19720 10852 19724 10908
rect 19724 10852 19780 10908
rect 19780 10852 19784 10908
rect 19720 10848 19784 10852
rect 5584 10364 5648 10368
rect 5584 10308 5588 10364
rect 5588 10308 5644 10364
rect 5644 10308 5648 10364
rect 5584 10304 5648 10308
rect 5664 10364 5728 10368
rect 5664 10308 5668 10364
rect 5668 10308 5724 10364
rect 5724 10308 5728 10364
rect 5664 10304 5728 10308
rect 5744 10364 5808 10368
rect 5744 10308 5748 10364
rect 5748 10308 5804 10364
rect 5804 10308 5808 10364
rect 5744 10304 5808 10308
rect 5824 10364 5888 10368
rect 5824 10308 5828 10364
rect 5828 10308 5884 10364
rect 5884 10308 5888 10364
rect 5824 10304 5888 10308
rect 14848 10364 14912 10368
rect 14848 10308 14852 10364
rect 14852 10308 14908 10364
rect 14908 10308 14912 10364
rect 14848 10304 14912 10308
rect 14928 10364 14992 10368
rect 14928 10308 14932 10364
rect 14932 10308 14988 10364
rect 14988 10308 14992 10364
rect 14928 10304 14992 10308
rect 15008 10364 15072 10368
rect 15008 10308 15012 10364
rect 15012 10308 15068 10364
rect 15068 10308 15072 10364
rect 15008 10304 15072 10308
rect 15088 10364 15152 10368
rect 15088 10308 15092 10364
rect 15092 10308 15148 10364
rect 15148 10308 15152 10364
rect 15088 10304 15152 10308
rect 24112 10364 24176 10368
rect 24112 10308 24116 10364
rect 24116 10308 24172 10364
rect 24172 10308 24176 10364
rect 24112 10304 24176 10308
rect 24192 10364 24256 10368
rect 24192 10308 24196 10364
rect 24196 10308 24252 10364
rect 24252 10308 24256 10364
rect 24192 10304 24256 10308
rect 24272 10364 24336 10368
rect 24272 10308 24276 10364
rect 24276 10308 24332 10364
rect 24332 10308 24336 10364
rect 24272 10304 24336 10308
rect 24352 10364 24416 10368
rect 24352 10308 24356 10364
rect 24356 10308 24412 10364
rect 24412 10308 24416 10364
rect 24352 10304 24416 10308
rect 19932 10160 19996 10164
rect 19932 10104 19982 10160
rect 19982 10104 19996 10160
rect 19932 10100 19996 10104
rect 10216 9820 10280 9824
rect 10216 9764 10220 9820
rect 10220 9764 10276 9820
rect 10276 9764 10280 9820
rect 10216 9760 10280 9764
rect 10296 9820 10360 9824
rect 10296 9764 10300 9820
rect 10300 9764 10356 9820
rect 10356 9764 10360 9820
rect 10296 9760 10360 9764
rect 10376 9820 10440 9824
rect 10376 9764 10380 9820
rect 10380 9764 10436 9820
rect 10436 9764 10440 9820
rect 10376 9760 10440 9764
rect 10456 9820 10520 9824
rect 10456 9764 10460 9820
rect 10460 9764 10516 9820
rect 10516 9764 10520 9820
rect 10456 9760 10520 9764
rect 19480 9820 19544 9824
rect 19480 9764 19484 9820
rect 19484 9764 19540 9820
rect 19540 9764 19544 9820
rect 19480 9760 19544 9764
rect 19560 9820 19624 9824
rect 19560 9764 19564 9820
rect 19564 9764 19620 9820
rect 19620 9764 19624 9820
rect 19560 9760 19624 9764
rect 19640 9820 19704 9824
rect 19640 9764 19644 9820
rect 19644 9764 19700 9820
rect 19700 9764 19704 9820
rect 19640 9760 19704 9764
rect 19720 9820 19784 9824
rect 19720 9764 19724 9820
rect 19724 9764 19780 9820
rect 19780 9764 19784 9820
rect 19720 9760 19784 9764
rect 5584 9276 5648 9280
rect 5584 9220 5588 9276
rect 5588 9220 5644 9276
rect 5644 9220 5648 9276
rect 5584 9216 5648 9220
rect 5664 9276 5728 9280
rect 5664 9220 5668 9276
rect 5668 9220 5724 9276
rect 5724 9220 5728 9276
rect 5664 9216 5728 9220
rect 5744 9276 5808 9280
rect 5744 9220 5748 9276
rect 5748 9220 5804 9276
rect 5804 9220 5808 9276
rect 5744 9216 5808 9220
rect 5824 9276 5888 9280
rect 5824 9220 5828 9276
rect 5828 9220 5884 9276
rect 5884 9220 5888 9276
rect 5824 9216 5888 9220
rect 14848 9276 14912 9280
rect 14848 9220 14852 9276
rect 14852 9220 14908 9276
rect 14908 9220 14912 9276
rect 14848 9216 14912 9220
rect 14928 9276 14992 9280
rect 14928 9220 14932 9276
rect 14932 9220 14988 9276
rect 14988 9220 14992 9276
rect 14928 9216 14992 9220
rect 15008 9276 15072 9280
rect 15008 9220 15012 9276
rect 15012 9220 15068 9276
rect 15068 9220 15072 9276
rect 15008 9216 15072 9220
rect 15088 9276 15152 9280
rect 15088 9220 15092 9276
rect 15092 9220 15148 9276
rect 15148 9220 15152 9276
rect 15088 9216 15152 9220
rect 24112 9276 24176 9280
rect 24112 9220 24116 9276
rect 24116 9220 24172 9276
rect 24172 9220 24176 9276
rect 24112 9216 24176 9220
rect 24192 9276 24256 9280
rect 24192 9220 24196 9276
rect 24196 9220 24252 9276
rect 24252 9220 24256 9276
rect 24192 9216 24256 9220
rect 24272 9276 24336 9280
rect 24272 9220 24276 9276
rect 24276 9220 24332 9276
rect 24332 9220 24336 9276
rect 24272 9216 24336 9220
rect 24352 9276 24416 9280
rect 24352 9220 24356 9276
rect 24356 9220 24412 9276
rect 24412 9220 24416 9276
rect 24352 9216 24416 9220
rect 10216 8732 10280 8736
rect 10216 8676 10220 8732
rect 10220 8676 10276 8732
rect 10276 8676 10280 8732
rect 10216 8672 10280 8676
rect 10296 8732 10360 8736
rect 10296 8676 10300 8732
rect 10300 8676 10356 8732
rect 10356 8676 10360 8732
rect 10296 8672 10360 8676
rect 10376 8732 10440 8736
rect 10376 8676 10380 8732
rect 10380 8676 10436 8732
rect 10436 8676 10440 8732
rect 10376 8672 10440 8676
rect 10456 8732 10520 8736
rect 10456 8676 10460 8732
rect 10460 8676 10516 8732
rect 10516 8676 10520 8732
rect 10456 8672 10520 8676
rect 19480 8732 19544 8736
rect 19480 8676 19484 8732
rect 19484 8676 19540 8732
rect 19540 8676 19544 8732
rect 19480 8672 19544 8676
rect 19560 8732 19624 8736
rect 19560 8676 19564 8732
rect 19564 8676 19620 8732
rect 19620 8676 19624 8732
rect 19560 8672 19624 8676
rect 19640 8732 19704 8736
rect 19640 8676 19644 8732
rect 19644 8676 19700 8732
rect 19700 8676 19704 8732
rect 19640 8672 19704 8676
rect 19720 8732 19784 8736
rect 19720 8676 19724 8732
rect 19724 8676 19780 8732
rect 19780 8676 19784 8732
rect 19720 8672 19784 8676
rect 13676 8664 13740 8668
rect 13676 8608 13690 8664
rect 13690 8608 13740 8664
rect 13676 8604 13740 8608
rect 5584 8188 5648 8192
rect 5584 8132 5588 8188
rect 5588 8132 5644 8188
rect 5644 8132 5648 8188
rect 5584 8128 5648 8132
rect 5664 8188 5728 8192
rect 5664 8132 5668 8188
rect 5668 8132 5724 8188
rect 5724 8132 5728 8188
rect 5664 8128 5728 8132
rect 5744 8188 5808 8192
rect 5744 8132 5748 8188
rect 5748 8132 5804 8188
rect 5804 8132 5808 8188
rect 5744 8128 5808 8132
rect 5824 8188 5888 8192
rect 5824 8132 5828 8188
rect 5828 8132 5884 8188
rect 5884 8132 5888 8188
rect 5824 8128 5888 8132
rect 14848 8188 14912 8192
rect 14848 8132 14852 8188
rect 14852 8132 14908 8188
rect 14908 8132 14912 8188
rect 14848 8128 14912 8132
rect 14928 8188 14992 8192
rect 14928 8132 14932 8188
rect 14932 8132 14988 8188
rect 14988 8132 14992 8188
rect 14928 8128 14992 8132
rect 15008 8188 15072 8192
rect 15008 8132 15012 8188
rect 15012 8132 15068 8188
rect 15068 8132 15072 8188
rect 15008 8128 15072 8132
rect 15088 8188 15152 8192
rect 15088 8132 15092 8188
rect 15092 8132 15148 8188
rect 15148 8132 15152 8188
rect 15088 8128 15152 8132
rect 24112 8188 24176 8192
rect 24112 8132 24116 8188
rect 24116 8132 24172 8188
rect 24172 8132 24176 8188
rect 24112 8128 24176 8132
rect 24192 8188 24256 8192
rect 24192 8132 24196 8188
rect 24196 8132 24252 8188
rect 24252 8132 24256 8188
rect 24192 8128 24256 8132
rect 24272 8188 24336 8192
rect 24272 8132 24276 8188
rect 24276 8132 24332 8188
rect 24332 8132 24336 8188
rect 24272 8128 24336 8132
rect 24352 8188 24416 8192
rect 24352 8132 24356 8188
rect 24356 8132 24412 8188
rect 24412 8132 24416 8188
rect 24352 8128 24416 8132
rect 10216 7644 10280 7648
rect 10216 7588 10220 7644
rect 10220 7588 10276 7644
rect 10276 7588 10280 7644
rect 10216 7584 10280 7588
rect 10296 7644 10360 7648
rect 10296 7588 10300 7644
rect 10300 7588 10356 7644
rect 10356 7588 10360 7644
rect 10296 7584 10360 7588
rect 10376 7644 10440 7648
rect 10376 7588 10380 7644
rect 10380 7588 10436 7644
rect 10436 7588 10440 7644
rect 10376 7584 10440 7588
rect 10456 7644 10520 7648
rect 10456 7588 10460 7644
rect 10460 7588 10516 7644
rect 10516 7588 10520 7644
rect 10456 7584 10520 7588
rect 19480 7644 19544 7648
rect 19480 7588 19484 7644
rect 19484 7588 19540 7644
rect 19540 7588 19544 7644
rect 19480 7584 19544 7588
rect 19560 7644 19624 7648
rect 19560 7588 19564 7644
rect 19564 7588 19620 7644
rect 19620 7588 19624 7644
rect 19560 7584 19624 7588
rect 19640 7644 19704 7648
rect 19640 7588 19644 7644
rect 19644 7588 19700 7644
rect 19700 7588 19704 7644
rect 19640 7584 19704 7588
rect 19720 7644 19784 7648
rect 19720 7588 19724 7644
rect 19724 7588 19780 7644
rect 19780 7588 19784 7644
rect 19720 7584 19784 7588
rect 5584 7100 5648 7104
rect 5584 7044 5588 7100
rect 5588 7044 5644 7100
rect 5644 7044 5648 7100
rect 5584 7040 5648 7044
rect 5664 7100 5728 7104
rect 5664 7044 5668 7100
rect 5668 7044 5724 7100
rect 5724 7044 5728 7100
rect 5664 7040 5728 7044
rect 5744 7100 5808 7104
rect 5744 7044 5748 7100
rect 5748 7044 5804 7100
rect 5804 7044 5808 7100
rect 5744 7040 5808 7044
rect 5824 7100 5888 7104
rect 5824 7044 5828 7100
rect 5828 7044 5884 7100
rect 5884 7044 5888 7100
rect 5824 7040 5888 7044
rect 14848 7100 14912 7104
rect 14848 7044 14852 7100
rect 14852 7044 14908 7100
rect 14908 7044 14912 7100
rect 14848 7040 14912 7044
rect 14928 7100 14992 7104
rect 14928 7044 14932 7100
rect 14932 7044 14988 7100
rect 14988 7044 14992 7100
rect 14928 7040 14992 7044
rect 15008 7100 15072 7104
rect 15008 7044 15012 7100
rect 15012 7044 15068 7100
rect 15068 7044 15072 7100
rect 15008 7040 15072 7044
rect 15088 7100 15152 7104
rect 15088 7044 15092 7100
rect 15092 7044 15148 7100
rect 15148 7044 15152 7100
rect 15088 7040 15152 7044
rect 24112 7100 24176 7104
rect 24112 7044 24116 7100
rect 24116 7044 24172 7100
rect 24172 7044 24176 7100
rect 24112 7040 24176 7044
rect 24192 7100 24256 7104
rect 24192 7044 24196 7100
rect 24196 7044 24252 7100
rect 24252 7044 24256 7100
rect 24192 7040 24256 7044
rect 24272 7100 24336 7104
rect 24272 7044 24276 7100
rect 24276 7044 24332 7100
rect 24332 7044 24336 7100
rect 24272 7040 24336 7044
rect 24352 7100 24416 7104
rect 24352 7044 24356 7100
rect 24356 7044 24412 7100
rect 24412 7044 24416 7100
rect 24352 7040 24416 7044
rect 13492 6896 13556 6900
rect 13492 6840 13506 6896
rect 13506 6840 13556 6896
rect 13492 6836 13556 6840
rect 10216 6556 10280 6560
rect 10216 6500 10220 6556
rect 10220 6500 10276 6556
rect 10276 6500 10280 6556
rect 10216 6496 10280 6500
rect 10296 6556 10360 6560
rect 10296 6500 10300 6556
rect 10300 6500 10356 6556
rect 10356 6500 10360 6556
rect 10296 6496 10360 6500
rect 10376 6556 10440 6560
rect 10376 6500 10380 6556
rect 10380 6500 10436 6556
rect 10436 6500 10440 6556
rect 10376 6496 10440 6500
rect 10456 6556 10520 6560
rect 10456 6500 10460 6556
rect 10460 6500 10516 6556
rect 10516 6500 10520 6556
rect 10456 6496 10520 6500
rect 19480 6556 19544 6560
rect 19480 6500 19484 6556
rect 19484 6500 19540 6556
rect 19540 6500 19544 6556
rect 19480 6496 19544 6500
rect 19560 6556 19624 6560
rect 19560 6500 19564 6556
rect 19564 6500 19620 6556
rect 19620 6500 19624 6556
rect 19560 6496 19624 6500
rect 19640 6556 19704 6560
rect 19640 6500 19644 6556
rect 19644 6500 19700 6556
rect 19700 6500 19704 6556
rect 19640 6496 19704 6500
rect 19720 6556 19784 6560
rect 19720 6500 19724 6556
rect 19724 6500 19780 6556
rect 19780 6500 19784 6556
rect 19720 6496 19784 6500
rect 5584 6012 5648 6016
rect 5584 5956 5588 6012
rect 5588 5956 5644 6012
rect 5644 5956 5648 6012
rect 5584 5952 5648 5956
rect 5664 6012 5728 6016
rect 5664 5956 5668 6012
rect 5668 5956 5724 6012
rect 5724 5956 5728 6012
rect 5664 5952 5728 5956
rect 5744 6012 5808 6016
rect 5744 5956 5748 6012
rect 5748 5956 5804 6012
rect 5804 5956 5808 6012
rect 5744 5952 5808 5956
rect 5824 6012 5888 6016
rect 5824 5956 5828 6012
rect 5828 5956 5884 6012
rect 5884 5956 5888 6012
rect 5824 5952 5888 5956
rect 14848 6012 14912 6016
rect 14848 5956 14852 6012
rect 14852 5956 14908 6012
rect 14908 5956 14912 6012
rect 14848 5952 14912 5956
rect 14928 6012 14992 6016
rect 14928 5956 14932 6012
rect 14932 5956 14988 6012
rect 14988 5956 14992 6012
rect 14928 5952 14992 5956
rect 15008 6012 15072 6016
rect 15008 5956 15012 6012
rect 15012 5956 15068 6012
rect 15068 5956 15072 6012
rect 15008 5952 15072 5956
rect 15088 6012 15152 6016
rect 15088 5956 15092 6012
rect 15092 5956 15148 6012
rect 15148 5956 15152 6012
rect 15088 5952 15152 5956
rect 24112 6012 24176 6016
rect 24112 5956 24116 6012
rect 24116 5956 24172 6012
rect 24172 5956 24176 6012
rect 24112 5952 24176 5956
rect 24192 6012 24256 6016
rect 24192 5956 24196 6012
rect 24196 5956 24252 6012
rect 24252 5956 24256 6012
rect 24192 5952 24256 5956
rect 24272 6012 24336 6016
rect 24272 5956 24276 6012
rect 24276 5956 24332 6012
rect 24332 5956 24336 6012
rect 24272 5952 24336 5956
rect 24352 6012 24416 6016
rect 24352 5956 24356 6012
rect 24356 5956 24412 6012
rect 24412 5956 24416 6012
rect 24352 5952 24416 5956
rect 10216 5468 10280 5472
rect 10216 5412 10220 5468
rect 10220 5412 10276 5468
rect 10276 5412 10280 5468
rect 10216 5408 10280 5412
rect 10296 5468 10360 5472
rect 10296 5412 10300 5468
rect 10300 5412 10356 5468
rect 10356 5412 10360 5468
rect 10296 5408 10360 5412
rect 10376 5468 10440 5472
rect 10376 5412 10380 5468
rect 10380 5412 10436 5468
rect 10436 5412 10440 5468
rect 10376 5408 10440 5412
rect 10456 5468 10520 5472
rect 10456 5412 10460 5468
rect 10460 5412 10516 5468
rect 10516 5412 10520 5468
rect 10456 5408 10520 5412
rect 19480 5468 19544 5472
rect 19480 5412 19484 5468
rect 19484 5412 19540 5468
rect 19540 5412 19544 5468
rect 19480 5408 19544 5412
rect 19560 5468 19624 5472
rect 19560 5412 19564 5468
rect 19564 5412 19620 5468
rect 19620 5412 19624 5468
rect 19560 5408 19624 5412
rect 19640 5468 19704 5472
rect 19640 5412 19644 5468
rect 19644 5412 19700 5468
rect 19700 5412 19704 5468
rect 19640 5408 19704 5412
rect 19720 5468 19784 5472
rect 19720 5412 19724 5468
rect 19724 5412 19780 5468
rect 19780 5412 19784 5468
rect 19720 5408 19784 5412
rect 5584 4924 5648 4928
rect 5584 4868 5588 4924
rect 5588 4868 5644 4924
rect 5644 4868 5648 4924
rect 5584 4864 5648 4868
rect 5664 4924 5728 4928
rect 5664 4868 5668 4924
rect 5668 4868 5724 4924
rect 5724 4868 5728 4924
rect 5664 4864 5728 4868
rect 5744 4924 5808 4928
rect 5744 4868 5748 4924
rect 5748 4868 5804 4924
rect 5804 4868 5808 4924
rect 5744 4864 5808 4868
rect 5824 4924 5888 4928
rect 5824 4868 5828 4924
rect 5828 4868 5884 4924
rect 5884 4868 5888 4924
rect 5824 4864 5888 4868
rect 14848 4924 14912 4928
rect 14848 4868 14852 4924
rect 14852 4868 14908 4924
rect 14908 4868 14912 4924
rect 14848 4864 14912 4868
rect 14928 4924 14992 4928
rect 14928 4868 14932 4924
rect 14932 4868 14988 4924
rect 14988 4868 14992 4924
rect 14928 4864 14992 4868
rect 15008 4924 15072 4928
rect 15008 4868 15012 4924
rect 15012 4868 15068 4924
rect 15068 4868 15072 4924
rect 15008 4864 15072 4868
rect 15088 4924 15152 4928
rect 15088 4868 15092 4924
rect 15092 4868 15148 4924
rect 15148 4868 15152 4924
rect 15088 4864 15152 4868
rect 24112 4924 24176 4928
rect 24112 4868 24116 4924
rect 24116 4868 24172 4924
rect 24172 4868 24176 4924
rect 24112 4864 24176 4868
rect 24192 4924 24256 4928
rect 24192 4868 24196 4924
rect 24196 4868 24252 4924
rect 24252 4868 24256 4924
rect 24192 4864 24256 4868
rect 24272 4924 24336 4928
rect 24272 4868 24276 4924
rect 24276 4868 24332 4924
rect 24332 4868 24336 4924
rect 24272 4864 24336 4868
rect 24352 4924 24416 4928
rect 24352 4868 24356 4924
rect 24356 4868 24412 4924
rect 24412 4868 24416 4924
rect 24352 4864 24416 4868
rect 10216 4380 10280 4384
rect 10216 4324 10220 4380
rect 10220 4324 10276 4380
rect 10276 4324 10280 4380
rect 10216 4320 10280 4324
rect 10296 4380 10360 4384
rect 10296 4324 10300 4380
rect 10300 4324 10356 4380
rect 10356 4324 10360 4380
rect 10296 4320 10360 4324
rect 10376 4380 10440 4384
rect 10376 4324 10380 4380
rect 10380 4324 10436 4380
rect 10436 4324 10440 4380
rect 10376 4320 10440 4324
rect 10456 4380 10520 4384
rect 10456 4324 10460 4380
rect 10460 4324 10516 4380
rect 10516 4324 10520 4380
rect 10456 4320 10520 4324
rect 19480 4380 19544 4384
rect 19480 4324 19484 4380
rect 19484 4324 19540 4380
rect 19540 4324 19544 4380
rect 19480 4320 19544 4324
rect 19560 4380 19624 4384
rect 19560 4324 19564 4380
rect 19564 4324 19620 4380
rect 19620 4324 19624 4380
rect 19560 4320 19624 4324
rect 19640 4380 19704 4384
rect 19640 4324 19644 4380
rect 19644 4324 19700 4380
rect 19700 4324 19704 4380
rect 19640 4320 19704 4324
rect 19720 4380 19784 4384
rect 19720 4324 19724 4380
rect 19724 4324 19780 4380
rect 19780 4324 19784 4380
rect 19720 4320 19784 4324
rect 5584 3836 5648 3840
rect 5584 3780 5588 3836
rect 5588 3780 5644 3836
rect 5644 3780 5648 3836
rect 5584 3776 5648 3780
rect 5664 3836 5728 3840
rect 5664 3780 5668 3836
rect 5668 3780 5724 3836
rect 5724 3780 5728 3836
rect 5664 3776 5728 3780
rect 5744 3836 5808 3840
rect 5744 3780 5748 3836
rect 5748 3780 5804 3836
rect 5804 3780 5808 3836
rect 5744 3776 5808 3780
rect 5824 3836 5888 3840
rect 5824 3780 5828 3836
rect 5828 3780 5884 3836
rect 5884 3780 5888 3836
rect 5824 3776 5888 3780
rect 14848 3836 14912 3840
rect 14848 3780 14852 3836
rect 14852 3780 14908 3836
rect 14908 3780 14912 3836
rect 14848 3776 14912 3780
rect 14928 3836 14992 3840
rect 14928 3780 14932 3836
rect 14932 3780 14988 3836
rect 14988 3780 14992 3836
rect 14928 3776 14992 3780
rect 15008 3836 15072 3840
rect 15008 3780 15012 3836
rect 15012 3780 15068 3836
rect 15068 3780 15072 3836
rect 15008 3776 15072 3780
rect 15088 3836 15152 3840
rect 15088 3780 15092 3836
rect 15092 3780 15148 3836
rect 15148 3780 15152 3836
rect 15088 3776 15152 3780
rect 24112 3836 24176 3840
rect 24112 3780 24116 3836
rect 24116 3780 24172 3836
rect 24172 3780 24176 3836
rect 24112 3776 24176 3780
rect 24192 3836 24256 3840
rect 24192 3780 24196 3836
rect 24196 3780 24252 3836
rect 24252 3780 24256 3836
rect 24192 3776 24256 3780
rect 24272 3836 24336 3840
rect 24272 3780 24276 3836
rect 24276 3780 24332 3836
rect 24332 3780 24336 3836
rect 24272 3776 24336 3780
rect 24352 3836 24416 3840
rect 24352 3780 24356 3836
rect 24356 3780 24412 3836
rect 24412 3780 24416 3836
rect 24352 3776 24416 3780
rect 10216 3292 10280 3296
rect 10216 3236 10220 3292
rect 10220 3236 10276 3292
rect 10276 3236 10280 3292
rect 10216 3232 10280 3236
rect 10296 3292 10360 3296
rect 10296 3236 10300 3292
rect 10300 3236 10356 3292
rect 10356 3236 10360 3292
rect 10296 3232 10360 3236
rect 10376 3292 10440 3296
rect 10376 3236 10380 3292
rect 10380 3236 10436 3292
rect 10436 3236 10440 3292
rect 10376 3232 10440 3236
rect 10456 3292 10520 3296
rect 10456 3236 10460 3292
rect 10460 3236 10516 3292
rect 10516 3236 10520 3292
rect 10456 3232 10520 3236
rect 19480 3292 19544 3296
rect 19480 3236 19484 3292
rect 19484 3236 19540 3292
rect 19540 3236 19544 3292
rect 19480 3232 19544 3236
rect 19560 3292 19624 3296
rect 19560 3236 19564 3292
rect 19564 3236 19620 3292
rect 19620 3236 19624 3292
rect 19560 3232 19624 3236
rect 19640 3292 19704 3296
rect 19640 3236 19644 3292
rect 19644 3236 19700 3292
rect 19700 3236 19704 3292
rect 19640 3232 19704 3236
rect 19720 3292 19784 3296
rect 19720 3236 19724 3292
rect 19724 3236 19780 3292
rect 19780 3236 19784 3292
rect 19720 3232 19784 3236
rect 5584 2748 5648 2752
rect 5584 2692 5588 2748
rect 5588 2692 5644 2748
rect 5644 2692 5648 2748
rect 5584 2688 5648 2692
rect 5664 2748 5728 2752
rect 5664 2692 5668 2748
rect 5668 2692 5724 2748
rect 5724 2692 5728 2748
rect 5664 2688 5728 2692
rect 5744 2748 5808 2752
rect 5744 2692 5748 2748
rect 5748 2692 5804 2748
rect 5804 2692 5808 2748
rect 5744 2688 5808 2692
rect 5824 2748 5888 2752
rect 5824 2692 5828 2748
rect 5828 2692 5884 2748
rect 5884 2692 5888 2748
rect 5824 2688 5888 2692
rect 14848 2748 14912 2752
rect 14848 2692 14852 2748
rect 14852 2692 14908 2748
rect 14908 2692 14912 2748
rect 14848 2688 14912 2692
rect 14928 2748 14992 2752
rect 14928 2692 14932 2748
rect 14932 2692 14988 2748
rect 14988 2692 14992 2748
rect 14928 2688 14992 2692
rect 15008 2748 15072 2752
rect 15008 2692 15012 2748
rect 15012 2692 15068 2748
rect 15068 2692 15072 2748
rect 15008 2688 15072 2692
rect 15088 2748 15152 2752
rect 15088 2692 15092 2748
rect 15092 2692 15148 2748
rect 15148 2692 15152 2748
rect 15088 2688 15152 2692
rect 24112 2748 24176 2752
rect 24112 2692 24116 2748
rect 24116 2692 24172 2748
rect 24172 2692 24176 2748
rect 24112 2688 24176 2692
rect 24192 2748 24256 2752
rect 24192 2692 24196 2748
rect 24196 2692 24252 2748
rect 24252 2692 24256 2748
rect 24192 2688 24256 2692
rect 24272 2748 24336 2752
rect 24272 2692 24276 2748
rect 24276 2692 24332 2748
rect 24332 2692 24336 2748
rect 24272 2688 24336 2692
rect 24352 2748 24416 2752
rect 24352 2692 24356 2748
rect 24356 2692 24412 2748
rect 24412 2692 24416 2748
rect 24352 2688 24416 2692
rect 10216 2204 10280 2208
rect 10216 2148 10220 2204
rect 10220 2148 10276 2204
rect 10276 2148 10280 2204
rect 10216 2144 10280 2148
rect 10296 2204 10360 2208
rect 10296 2148 10300 2204
rect 10300 2148 10356 2204
rect 10356 2148 10360 2204
rect 10296 2144 10360 2148
rect 10376 2204 10440 2208
rect 10376 2148 10380 2204
rect 10380 2148 10436 2204
rect 10436 2148 10440 2204
rect 10376 2144 10440 2148
rect 10456 2204 10520 2208
rect 10456 2148 10460 2204
rect 10460 2148 10516 2204
rect 10516 2148 10520 2204
rect 10456 2144 10520 2148
rect 19480 2204 19544 2208
rect 19480 2148 19484 2204
rect 19484 2148 19540 2204
rect 19540 2148 19544 2204
rect 19480 2144 19544 2148
rect 19560 2204 19624 2208
rect 19560 2148 19564 2204
rect 19564 2148 19620 2204
rect 19620 2148 19624 2204
rect 19560 2144 19624 2148
rect 19640 2204 19704 2208
rect 19640 2148 19644 2204
rect 19644 2148 19700 2204
rect 19700 2148 19704 2204
rect 19640 2144 19704 2148
rect 19720 2204 19784 2208
rect 19720 2148 19724 2204
rect 19724 2148 19780 2204
rect 19780 2148 19784 2204
rect 19720 2144 19784 2148
<< metal4 >>
rect 5576 27776 5896 27792
rect 5576 27712 5584 27776
rect 5648 27712 5664 27776
rect 5728 27712 5744 27776
rect 5808 27712 5824 27776
rect 5888 27712 5896 27776
rect 5576 26688 5896 27712
rect 5576 26624 5584 26688
rect 5648 26624 5664 26688
rect 5728 26624 5744 26688
rect 5808 26624 5824 26688
rect 5888 26624 5896 26688
rect 5576 25600 5896 26624
rect 5576 25536 5584 25600
rect 5648 25536 5664 25600
rect 5728 25536 5744 25600
rect 5808 25536 5824 25600
rect 5888 25536 5896 25600
rect 5576 24512 5896 25536
rect 5576 24448 5584 24512
rect 5648 24448 5664 24512
rect 5728 24448 5744 24512
rect 5808 24448 5824 24512
rect 5888 24448 5896 24512
rect 5576 23424 5896 24448
rect 5576 23360 5584 23424
rect 5648 23360 5664 23424
rect 5728 23360 5744 23424
rect 5808 23360 5824 23424
rect 5888 23360 5896 23424
rect 5576 22336 5896 23360
rect 5576 22272 5584 22336
rect 5648 22272 5664 22336
rect 5728 22272 5744 22336
rect 5808 22272 5824 22336
rect 5888 22272 5896 22336
rect 5576 21248 5896 22272
rect 5576 21184 5584 21248
rect 5648 21184 5664 21248
rect 5728 21184 5744 21248
rect 5808 21184 5824 21248
rect 5888 21184 5896 21248
rect 5576 20160 5896 21184
rect 5576 20096 5584 20160
rect 5648 20096 5664 20160
rect 5728 20096 5744 20160
rect 5808 20096 5824 20160
rect 5888 20096 5896 20160
rect 5576 19072 5896 20096
rect 5576 19008 5584 19072
rect 5648 19008 5664 19072
rect 5728 19008 5744 19072
rect 5808 19008 5824 19072
rect 5888 19008 5896 19072
rect 5576 17984 5896 19008
rect 5576 17920 5584 17984
rect 5648 17920 5664 17984
rect 5728 17920 5744 17984
rect 5808 17920 5824 17984
rect 5888 17920 5896 17984
rect 5576 16896 5896 17920
rect 5576 16832 5584 16896
rect 5648 16832 5664 16896
rect 5728 16832 5744 16896
rect 5808 16832 5824 16896
rect 5888 16832 5896 16896
rect 5576 15808 5896 16832
rect 5576 15744 5584 15808
rect 5648 15744 5664 15808
rect 5728 15744 5744 15808
rect 5808 15744 5824 15808
rect 5888 15744 5896 15808
rect 5576 14720 5896 15744
rect 5576 14656 5584 14720
rect 5648 14656 5664 14720
rect 5728 14656 5744 14720
rect 5808 14656 5824 14720
rect 5888 14656 5896 14720
rect 5576 13632 5896 14656
rect 5576 13568 5584 13632
rect 5648 13568 5664 13632
rect 5728 13568 5744 13632
rect 5808 13568 5824 13632
rect 5888 13568 5896 13632
rect 5576 12544 5896 13568
rect 5576 12480 5584 12544
rect 5648 12480 5664 12544
rect 5728 12480 5744 12544
rect 5808 12480 5824 12544
rect 5888 12480 5896 12544
rect 5576 11456 5896 12480
rect 5576 11392 5584 11456
rect 5648 11392 5664 11456
rect 5728 11392 5744 11456
rect 5808 11392 5824 11456
rect 5888 11392 5896 11456
rect 5576 10368 5896 11392
rect 5576 10304 5584 10368
rect 5648 10304 5664 10368
rect 5728 10304 5744 10368
rect 5808 10304 5824 10368
rect 5888 10304 5896 10368
rect 5576 9280 5896 10304
rect 5576 9216 5584 9280
rect 5648 9216 5664 9280
rect 5728 9216 5744 9280
rect 5808 9216 5824 9280
rect 5888 9216 5896 9280
rect 5576 8192 5896 9216
rect 5576 8128 5584 8192
rect 5648 8128 5664 8192
rect 5728 8128 5744 8192
rect 5808 8128 5824 8192
rect 5888 8128 5896 8192
rect 5576 7104 5896 8128
rect 5576 7040 5584 7104
rect 5648 7040 5664 7104
rect 5728 7040 5744 7104
rect 5808 7040 5824 7104
rect 5888 7040 5896 7104
rect 5576 6016 5896 7040
rect 5576 5952 5584 6016
rect 5648 5952 5664 6016
rect 5728 5952 5744 6016
rect 5808 5952 5824 6016
rect 5888 5952 5896 6016
rect 5576 4928 5896 5952
rect 5576 4864 5584 4928
rect 5648 4864 5664 4928
rect 5728 4864 5744 4928
rect 5808 4864 5824 4928
rect 5888 4864 5896 4928
rect 5576 3840 5896 4864
rect 5576 3776 5584 3840
rect 5648 3776 5664 3840
rect 5728 3776 5744 3840
rect 5808 3776 5824 3840
rect 5888 3776 5896 3840
rect 5576 2752 5896 3776
rect 5576 2688 5584 2752
rect 5648 2688 5664 2752
rect 5728 2688 5744 2752
rect 5808 2688 5824 2752
rect 5888 2688 5896 2752
rect 5576 2128 5896 2688
rect 10208 27232 10528 27792
rect 10208 27168 10216 27232
rect 10280 27168 10296 27232
rect 10360 27168 10376 27232
rect 10440 27168 10456 27232
rect 10520 27168 10528 27232
rect 10208 26144 10528 27168
rect 10208 26080 10216 26144
rect 10280 26080 10296 26144
rect 10360 26080 10376 26144
rect 10440 26080 10456 26144
rect 10520 26080 10528 26144
rect 10208 25056 10528 26080
rect 10208 24992 10216 25056
rect 10280 24992 10296 25056
rect 10360 24992 10376 25056
rect 10440 24992 10456 25056
rect 10520 24992 10528 25056
rect 10208 23968 10528 24992
rect 10208 23904 10216 23968
rect 10280 23904 10296 23968
rect 10360 23904 10376 23968
rect 10440 23904 10456 23968
rect 10520 23904 10528 23968
rect 10208 22880 10528 23904
rect 10208 22816 10216 22880
rect 10280 22816 10296 22880
rect 10360 22816 10376 22880
rect 10440 22816 10456 22880
rect 10520 22816 10528 22880
rect 10208 21792 10528 22816
rect 10208 21728 10216 21792
rect 10280 21728 10296 21792
rect 10360 21728 10376 21792
rect 10440 21728 10456 21792
rect 10520 21728 10528 21792
rect 10208 20704 10528 21728
rect 14840 27776 15160 27792
rect 14840 27712 14848 27776
rect 14912 27712 14928 27776
rect 14992 27712 15008 27776
rect 15072 27712 15088 27776
rect 15152 27712 15160 27776
rect 14840 26688 15160 27712
rect 14840 26624 14848 26688
rect 14912 26624 14928 26688
rect 14992 26624 15008 26688
rect 15072 26624 15088 26688
rect 15152 26624 15160 26688
rect 14840 25600 15160 26624
rect 14840 25536 14848 25600
rect 14912 25536 14928 25600
rect 14992 25536 15008 25600
rect 15072 25536 15088 25600
rect 15152 25536 15160 25600
rect 14840 24512 15160 25536
rect 19472 27232 19792 27792
rect 19472 27168 19480 27232
rect 19544 27168 19560 27232
rect 19624 27168 19640 27232
rect 19704 27168 19720 27232
rect 19784 27168 19792 27232
rect 19472 26144 19792 27168
rect 19472 26080 19480 26144
rect 19544 26080 19560 26144
rect 19624 26080 19640 26144
rect 19704 26080 19720 26144
rect 19784 26080 19792 26144
rect 19472 25056 19792 26080
rect 19472 24992 19480 25056
rect 19544 24992 19560 25056
rect 19624 24992 19640 25056
rect 19704 24992 19720 25056
rect 19784 24992 19792 25056
rect 16435 24988 16501 24989
rect 16435 24924 16436 24988
rect 16500 24924 16501 24988
rect 16435 24923 16501 24924
rect 14840 24448 14848 24512
rect 14912 24448 14928 24512
rect 14992 24448 15008 24512
rect 15072 24448 15088 24512
rect 15152 24448 15160 24512
rect 14840 23424 15160 24448
rect 14840 23360 14848 23424
rect 14912 23360 14928 23424
rect 14992 23360 15008 23424
rect 15072 23360 15088 23424
rect 15152 23360 15160 23424
rect 14840 22336 15160 23360
rect 14840 22272 14848 22336
rect 14912 22272 14928 22336
rect 14992 22272 15008 22336
rect 15072 22272 15088 22336
rect 15152 22272 15160 22336
rect 14840 21248 15160 22272
rect 14840 21184 14848 21248
rect 14912 21184 14928 21248
rect 14992 21184 15008 21248
rect 15072 21184 15088 21248
rect 15152 21184 15160 21248
rect 14595 20908 14661 20909
rect 14595 20844 14596 20908
rect 14660 20844 14661 20908
rect 14595 20843 14661 20844
rect 10208 20640 10216 20704
rect 10280 20640 10296 20704
rect 10360 20640 10376 20704
rect 10440 20640 10456 20704
rect 10520 20640 10528 20704
rect 10208 19616 10528 20640
rect 10208 19552 10216 19616
rect 10280 19552 10296 19616
rect 10360 19552 10376 19616
rect 10440 19552 10456 19616
rect 10520 19552 10528 19616
rect 10208 18528 10528 19552
rect 10208 18464 10216 18528
rect 10280 18464 10296 18528
rect 10360 18464 10376 18528
rect 10440 18464 10456 18528
rect 10520 18464 10528 18528
rect 10208 17440 10528 18464
rect 10208 17376 10216 17440
rect 10280 17376 10296 17440
rect 10360 17376 10376 17440
rect 10440 17376 10456 17440
rect 10520 17376 10528 17440
rect 10208 16352 10528 17376
rect 13859 16692 13925 16693
rect 13859 16628 13860 16692
rect 13924 16628 13925 16692
rect 13859 16627 13925 16628
rect 10208 16288 10216 16352
rect 10280 16288 10296 16352
rect 10360 16288 10376 16352
rect 10440 16288 10456 16352
rect 10520 16288 10528 16352
rect 10208 15264 10528 16288
rect 13491 15332 13557 15333
rect 13491 15268 13492 15332
rect 13556 15268 13557 15332
rect 13491 15267 13557 15268
rect 10208 15200 10216 15264
rect 10280 15200 10296 15264
rect 10360 15200 10376 15264
rect 10440 15200 10456 15264
rect 10520 15200 10528 15264
rect 10208 14176 10528 15200
rect 10208 14112 10216 14176
rect 10280 14112 10296 14176
rect 10360 14112 10376 14176
rect 10440 14112 10456 14176
rect 10520 14112 10528 14176
rect 10208 13088 10528 14112
rect 10208 13024 10216 13088
rect 10280 13024 10296 13088
rect 10360 13024 10376 13088
rect 10440 13024 10456 13088
rect 10520 13024 10528 13088
rect 10208 12000 10528 13024
rect 10208 11936 10216 12000
rect 10280 11936 10296 12000
rect 10360 11936 10376 12000
rect 10440 11936 10456 12000
rect 10520 11936 10528 12000
rect 10208 10912 10528 11936
rect 10208 10848 10216 10912
rect 10280 10848 10296 10912
rect 10360 10848 10376 10912
rect 10440 10848 10456 10912
rect 10520 10848 10528 10912
rect 10208 9824 10528 10848
rect 10208 9760 10216 9824
rect 10280 9760 10296 9824
rect 10360 9760 10376 9824
rect 10440 9760 10456 9824
rect 10520 9760 10528 9824
rect 10208 8736 10528 9760
rect 10208 8672 10216 8736
rect 10280 8672 10296 8736
rect 10360 8672 10376 8736
rect 10440 8672 10456 8736
rect 10520 8672 10528 8736
rect 10208 7648 10528 8672
rect 10208 7584 10216 7648
rect 10280 7584 10296 7648
rect 10360 7584 10376 7648
rect 10440 7584 10456 7648
rect 10520 7584 10528 7648
rect 10208 6560 10528 7584
rect 13494 6901 13554 15267
rect 13862 15061 13922 16627
rect 13859 15060 13925 15061
rect 13859 14996 13860 15060
rect 13924 14996 13925 15060
rect 13859 14995 13925 14996
rect 14598 12069 14658 20843
rect 14840 20160 15160 21184
rect 14840 20096 14848 20160
rect 14912 20096 14928 20160
rect 14992 20096 15008 20160
rect 15072 20096 15088 20160
rect 15152 20096 15160 20160
rect 14840 19072 15160 20096
rect 14840 19008 14848 19072
rect 14912 19008 14928 19072
rect 14992 19008 15008 19072
rect 15072 19008 15088 19072
rect 15152 19008 15160 19072
rect 14840 17984 15160 19008
rect 16438 18461 16498 24923
rect 19472 23968 19792 24992
rect 19472 23904 19480 23968
rect 19544 23904 19560 23968
rect 19624 23904 19640 23968
rect 19704 23904 19720 23968
rect 19784 23904 19792 23968
rect 19472 22880 19792 23904
rect 19472 22816 19480 22880
rect 19544 22816 19560 22880
rect 19624 22816 19640 22880
rect 19704 22816 19720 22880
rect 19784 22816 19792 22880
rect 19472 21792 19792 22816
rect 19472 21728 19480 21792
rect 19544 21728 19560 21792
rect 19624 21728 19640 21792
rect 19704 21728 19720 21792
rect 19784 21728 19792 21792
rect 19472 20704 19792 21728
rect 19472 20640 19480 20704
rect 19544 20640 19560 20704
rect 19624 20640 19640 20704
rect 19704 20640 19720 20704
rect 19784 20640 19792 20704
rect 19472 19616 19792 20640
rect 19472 19552 19480 19616
rect 19544 19552 19560 19616
rect 19624 19552 19640 19616
rect 19704 19552 19720 19616
rect 19784 19552 19792 19616
rect 19472 18528 19792 19552
rect 19472 18464 19480 18528
rect 19544 18464 19560 18528
rect 19624 18464 19640 18528
rect 19704 18464 19720 18528
rect 19784 18464 19792 18528
rect 16435 18460 16501 18461
rect 16435 18396 16436 18460
rect 16500 18396 16501 18460
rect 16435 18395 16501 18396
rect 14840 17920 14848 17984
rect 14912 17920 14928 17984
rect 14992 17920 15008 17984
rect 15072 17920 15088 17984
rect 15152 17920 15160 17984
rect 14840 16896 15160 17920
rect 14840 16832 14848 16896
rect 14912 16832 14928 16896
rect 14992 16832 15008 16896
rect 15072 16832 15088 16896
rect 15152 16832 15160 16896
rect 14840 15808 15160 16832
rect 14840 15744 14848 15808
rect 14912 15744 14928 15808
rect 14992 15744 15008 15808
rect 15072 15744 15088 15808
rect 15152 15744 15160 15808
rect 14840 14720 15160 15744
rect 14840 14656 14848 14720
rect 14912 14656 14928 14720
rect 14992 14656 15008 14720
rect 15072 14656 15088 14720
rect 15152 14656 15160 14720
rect 14840 13632 15160 14656
rect 14840 13568 14848 13632
rect 14912 13568 14928 13632
rect 14992 13568 15008 13632
rect 15072 13568 15088 13632
rect 15152 13568 15160 13632
rect 14840 12544 15160 13568
rect 14840 12480 14848 12544
rect 14912 12480 14928 12544
rect 14992 12480 15008 12544
rect 15072 12480 15088 12544
rect 15152 12480 15160 12544
rect 13675 12068 13741 12069
rect 13675 12004 13676 12068
rect 13740 12004 13741 12068
rect 13675 12003 13741 12004
rect 14595 12068 14661 12069
rect 14595 12004 14596 12068
rect 14660 12004 14661 12068
rect 14595 12003 14661 12004
rect 13678 8669 13738 12003
rect 14840 11456 15160 12480
rect 14840 11392 14848 11456
rect 14912 11392 14928 11456
rect 14992 11392 15008 11456
rect 15072 11392 15088 11456
rect 15152 11392 15160 11456
rect 14840 10368 15160 11392
rect 14840 10304 14848 10368
rect 14912 10304 14928 10368
rect 14992 10304 15008 10368
rect 15072 10304 15088 10368
rect 15152 10304 15160 10368
rect 14840 9280 15160 10304
rect 14840 9216 14848 9280
rect 14912 9216 14928 9280
rect 14992 9216 15008 9280
rect 15072 9216 15088 9280
rect 15152 9216 15160 9280
rect 13675 8668 13741 8669
rect 13675 8604 13676 8668
rect 13740 8604 13741 8668
rect 13675 8603 13741 8604
rect 14840 8192 15160 9216
rect 14840 8128 14848 8192
rect 14912 8128 14928 8192
rect 14992 8128 15008 8192
rect 15072 8128 15088 8192
rect 15152 8128 15160 8192
rect 14840 7104 15160 8128
rect 14840 7040 14848 7104
rect 14912 7040 14928 7104
rect 14992 7040 15008 7104
rect 15072 7040 15088 7104
rect 15152 7040 15160 7104
rect 13491 6900 13557 6901
rect 13491 6836 13492 6900
rect 13556 6836 13557 6900
rect 13491 6835 13557 6836
rect 10208 6496 10216 6560
rect 10280 6496 10296 6560
rect 10360 6496 10376 6560
rect 10440 6496 10456 6560
rect 10520 6496 10528 6560
rect 10208 5472 10528 6496
rect 10208 5408 10216 5472
rect 10280 5408 10296 5472
rect 10360 5408 10376 5472
rect 10440 5408 10456 5472
rect 10520 5408 10528 5472
rect 10208 4384 10528 5408
rect 10208 4320 10216 4384
rect 10280 4320 10296 4384
rect 10360 4320 10376 4384
rect 10440 4320 10456 4384
rect 10520 4320 10528 4384
rect 10208 3296 10528 4320
rect 10208 3232 10216 3296
rect 10280 3232 10296 3296
rect 10360 3232 10376 3296
rect 10440 3232 10456 3296
rect 10520 3232 10528 3296
rect 10208 2208 10528 3232
rect 10208 2144 10216 2208
rect 10280 2144 10296 2208
rect 10360 2144 10376 2208
rect 10440 2144 10456 2208
rect 10520 2144 10528 2208
rect 10208 2128 10528 2144
rect 14840 6016 15160 7040
rect 14840 5952 14848 6016
rect 14912 5952 14928 6016
rect 14992 5952 15008 6016
rect 15072 5952 15088 6016
rect 15152 5952 15160 6016
rect 14840 4928 15160 5952
rect 14840 4864 14848 4928
rect 14912 4864 14928 4928
rect 14992 4864 15008 4928
rect 15072 4864 15088 4928
rect 15152 4864 15160 4928
rect 14840 3840 15160 4864
rect 14840 3776 14848 3840
rect 14912 3776 14928 3840
rect 14992 3776 15008 3840
rect 15072 3776 15088 3840
rect 15152 3776 15160 3840
rect 14840 2752 15160 3776
rect 14840 2688 14848 2752
rect 14912 2688 14928 2752
rect 14992 2688 15008 2752
rect 15072 2688 15088 2752
rect 15152 2688 15160 2752
rect 14840 2128 15160 2688
rect 19472 17440 19792 18464
rect 19472 17376 19480 17440
rect 19544 17376 19560 17440
rect 19624 17376 19640 17440
rect 19704 17376 19720 17440
rect 19784 17376 19792 17440
rect 19472 16352 19792 17376
rect 19472 16288 19480 16352
rect 19544 16288 19560 16352
rect 19624 16288 19640 16352
rect 19704 16288 19720 16352
rect 19784 16288 19792 16352
rect 19472 15264 19792 16288
rect 24104 27776 24424 27792
rect 24104 27712 24112 27776
rect 24176 27712 24192 27776
rect 24256 27712 24272 27776
rect 24336 27712 24352 27776
rect 24416 27712 24424 27776
rect 24104 26688 24424 27712
rect 24104 26624 24112 26688
rect 24176 26624 24192 26688
rect 24256 26624 24272 26688
rect 24336 26624 24352 26688
rect 24416 26624 24424 26688
rect 24104 25600 24424 26624
rect 25635 26348 25701 26349
rect 25635 26284 25636 26348
rect 25700 26284 25701 26348
rect 25635 26283 25701 26284
rect 24104 25536 24112 25600
rect 24176 25536 24192 25600
rect 24256 25536 24272 25600
rect 24336 25536 24352 25600
rect 24416 25536 24424 25600
rect 24104 24512 24424 25536
rect 24104 24448 24112 24512
rect 24176 24448 24192 24512
rect 24256 24448 24272 24512
rect 24336 24448 24352 24512
rect 24416 24448 24424 24512
rect 24104 23424 24424 24448
rect 24104 23360 24112 23424
rect 24176 23360 24192 23424
rect 24256 23360 24272 23424
rect 24336 23360 24352 23424
rect 24416 23360 24424 23424
rect 24104 22336 24424 23360
rect 24104 22272 24112 22336
rect 24176 22272 24192 22336
rect 24256 22272 24272 22336
rect 24336 22272 24352 22336
rect 24416 22272 24424 22336
rect 24104 21248 24424 22272
rect 24104 21184 24112 21248
rect 24176 21184 24192 21248
rect 24256 21184 24272 21248
rect 24336 21184 24352 21248
rect 24416 21184 24424 21248
rect 24104 20160 24424 21184
rect 24104 20096 24112 20160
rect 24176 20096 24192 20160
rect 24256 20096 24272 20160
rect 24336 20096 24352 20160
rect 24416 20096 24424 20160
rect 24104 19072 24424 20096
rect 24104 19008 24112 19072
rect 24176 19008 24192 19072
rect 24256 19008 24272 19072
rect 24336 19008 24352 19072
rect 24416 19008 24424 19072
rect 24104 17984 24424 19008
rect 24104 17920 24112 17984
rect 24176 17920 24192 17984
rect 24256 17920 24272 17984
rect 24336 17920 24352 17984
rect 24416 17920 24424 17984
rect 24104 16896 24424 17920
rect 25638 17781 25698 26283
rect 25635 17780 25701 17781
rect 25635 17716 25636 17780
rect 25700 17716 25701 17780
rect 25635 17715 25701 17716
rect 24104 16832 24112 16896
rect 24176 16832 24192 16896
rect 24256 16832 24272 16896
rect 24336 16832 24352 16896
rect 24416 16832 24424 16896
rect 24104 15808 24424 16832
rect 24104 15744 24112 15808
rect 24176 15744 24192 15808
rect 24256 15744 24272 15808
rect 24336 15744 24352 15808
rect 24416 15744 24424 15808
rect 19931 15468 19997 15469
rect 19931 15404 19932 15468
rect 19996 15404 19997 15468
rect 19931 15403 19997 15404
rect 19472 15200 19480 15264
rect 19544 15200 19560 15264
rect 19624 15200 19640 15264
rect 19704 15200 19720 15264
rect 19784 15200 19792 15264
rect 19472 14176 19792 15200
rect 19472 14112 19480 14176
rect 19544 14112 19560 14176
rect 19624 14112 19640 14176
rect 19704 14112 19720 14176
rect 19784 14112 19792 14176
rect 19472 13088 19792 14112
rect 19472 13024 19480 13088
rect 19544 13024 19560 13088
rect 19624 13024 19640 13088
rect 19704 13024 19720 13088
rect 19784 13024 19792 13088
rect 19472 12000 19792 13024
rect 19472 11936 19480 12000
rect 19544 11936 19560 12000
rect 19624 11936 19640 12000
rect 19704 11936 19720 12000
rect 19784 11936 19792 12000
rect 19472 10912 19792 11936
rect 19472 10848 19480 10912
rect 19544 10848 19560 10912
rect 19624 10848 19640 10912
rect 19704 10848 19720 10912
rect 19784 10848 19792 10912
rect 19472 9824 19792 10848
rect 19934 10165 19994 15403
rect 24104 14720 24424 15744
rect 24104 14656 24112 14720
rect 24176 14656 24192 14720
rect 24256 14656 24272 14720
rect 24336 14656 24352 14720
rect 24416 14656 24424 14720
rect 24104 13632 24424 14656
rect 24104 13568 24112 13632
rect 24176 13568 24192 13632
rect 24256 13568 24272 13632
rect 24336 13568 24352 13632
rect 24416 13568 24424 13632
rect 24104 12544 24424 13568
rect 24104 12480 24112 12544
rect 24176 12480 24192 12544
rect 24256 12480 24272 12544
rect 24336 12480 24352 12544
rect 24416 12480 24424 12544
rect 24104 11456 24424 12480
rect 24104 11392 24112 11456
rect 24176 11392 24192 11456
rect 24256 11392 24272 11456
rect 24336 11392 24352 11456
rect 24416 11392 24424 11456
rect 24104 10368 24424 11392
rect 24104 10304 24112 10368
rect 24176 10304 24192 10368
rect 24256 10304 24272 10368
rect 24336 10304 24352 10368
rect 24416 10304 24424 10368
rect 19931 10164 19997 10165
rect 19931 10100 19932 10164
rect 19996 10100 19997 10164
rect 19931 10099 19997 10100
rect 19472 9760 19480 9824
rect 19544 9760 19560 9824
rect 19624 9760 19640 9824
rect 19704 9760 19720 9824
rect 19784 9760 19792 9824
rect 19472 8736 19792 9760
rect 19472 8672 19480 8736
rect 19544 8672 19560 8736
rect 19624 8672 19640 8736
rect 19704 8672 19720 8736
rect 19784 8672 19792 8736
rect 19472 7648 19792 8672
rect 19472 7584 19480 7648
rect 19544 7584 19560 7648
rect 19624 7584 19640 7648
rect 19704 7584 19720 7648
rect 19784 7584 19792 7648
rect 19472 6560 19792 7584
rect 19472 6496 19480 6560
rect 19544 6496 19560 6560
rect 19624 6496 19640 6560
rect 19704 6496 19720 6560
rect 19784 6496 19792 6560
rect 19472 5472 19792 6496
rect 19472 5408 19480 5472
rect 19544 5408 19560 5472
rect 19624 5408 19640 5472
rect 19704 5408 19720 5472
rect 19784 5408 19792 5472
rect 19472 4384 19792 5408
rect 19472 4320 19480 4384
rect 19544 4320 19560 4384
rect 19624 4320 19640 4384
rect 19704 4320 19720 4384
rect 19784 4320 19792 4384
rect 19472 3296 19792 4320
rect 19472 3232 19480 3296
rect 19544 3232 19560 3296
rect 19624 3232 19640 3296
rect 19704 3232 19720 3296
rect 19784 3232 19792 3296
rect 19472 2208 19792 3232
rect 19472 2144 19480 2208
rect 19544 2144 19560 2208
rect 19624 2144 19640 2208
rect 19704 2144 19720 2208
rect 19784 2144 19792 2208
rect 19472 2128 19792 2144
rect 24104 9280 24424 10304
rect 24104 9216 24112 9280
rect 24176 9216 24192 9280
rect 24256 9216 24272 9280
rect 24336 9216 24352 9280
rect 24416 9216 24424 9280
rect 24104 8192 24424 9216
rect 24104 8128 24112 8192
rect 24176 8128 24192 8192
rect 24256 8128 24272 8192
rect 24336 8128 24352 8192
rect 24416 8128 24424 8192
rect 24104 7104 24424 8128
rect 24104 7040 24112 7104
rect 24176 7040 24192 7104
rect 24256 7040 24272 7104
rect 24336 7040 24352 7104
rect 24416 7040 24424 7104
rect 24104 6016 24424 7040
rect 24104 5952 24112 6016
rect 24176 5952 24192 6016
rect 24256 5952 24272 6016
rect 24336 5952 24352 6016
rect 24416 5952 24424 6016
rect 24104 4928 24424 5952
rect 24104 4864 24112 4928
rect 24176 4864 24192 4928
rect 24256 4864 24272 4928
rect 24336 4864 24352 4928
rect 24416 4864 24424 4928
rect 24104 3840 24424 4864
rect 24104 3776 24112 3840
rect 24176 3776 24192 3840
rect 24256 3776 24272 3840
rect 24336 3776 24352 3840
rect 24416 3776 24424 3840
rect 24104 2752 24424 3776
rect 24104 2688 24112 2752
rect 24176 2688 24192 2752
rect 24256 2688 24272 2752
rect 24336 2688 24352 2752
rect 24416 2688 24424 2752
rect 24104 2128 24424 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__C
timestamp 1644511149
transform -1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__A_N
timestamp 1644511149
transform 1 0 18308 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__B
timestamp 1644511149
transform 1 0 18676 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__C
timestamp 1644511149
transform -1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A
timestamp 1644511149
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__B
timestamp 1644511149
transform -1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__A0
timestamp 1644511149
transform 1 0 25392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__A0
timestamp 1644511149
transform -1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A0
timestamp 1644511149
transform 1 0 17480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__A0
timestamp 1644511149
transform 1 0 21528 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A0
timestamp 1644511149
transform 1 0 15916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A0
timestamp 1644511149
transform 1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__A0
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A0
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A
timestamp 1644511149
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__B
timestamp 1644511149
transform -1 0 21252 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A
timestamp 1644511149
transform 1 0 20700 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__B
timestamp 1644511149
transform -1 0 18492 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A1
timestamp 1644511149
transform 1 0 12696 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A1
timestamp 1644511149
transform 1 0 13156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A1
timestamp 1644511149
transform 1 0 10764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A1
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A1
timestamp 1644511149
transform -1 0 10580 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A1
timestamp 1644511149
transform 1 0 12696 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A1
timestamp 1644511149
transform -1 0 11960 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A1
timestamp 1644511149
transform 1 0 14720 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A
timestamp 1644511149
transform 1 0 17848 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__C_N
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A0
timestamp 1644511149
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A0
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A0
timestamp 1644511149
transform 1 0 12144 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A0
timestamp 1644511149
transform -1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A0
timestamp 1644511149
transform 1 0 14536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A0
timestamp 1644511149
transform 1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A0
timestamp 1644511149
transform 1 0 19596 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A0
timestamp 1644511149
transform 1 0 14904 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A0
timestamp 1644511149
transform 1 0 12512 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A0
timestamp 1644511149
transform 1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A0
timestamp 1644511149
transform 1 0 14628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A0
timestamp 1644511149
transform -1 0 16836 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A0
timestamp 1644511149
transform -1 0 13524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A0
timestamp 1644511149
transform -1 0 14260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A_N
timestamp 1644511149
transform -1 0 20240 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B
timestamp 1644511149
transform 1 0 13248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__C
timestamp 1644511149
transform 1 0 23184 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A0
timestamp 1644511149
transform -1 0 18860 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A0
timestamp 1644511149
transform 1 0 18216 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A0
timestamp 1644511149
transform -1 0 18768 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A0
timestamp 1644511149
transform -1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A0
timestamp 1644511149
transform -1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B1
timestamp 1644511149
transform -1 0 18216 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1
timestamp 1644511149
transform 1 0 18676 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A0
timestamp 1644511149
transform 1 0 17112 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A0
timestamp 1644511149
transform 1 0 16376 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A
timestamp 1644511149
transform -1 0 20424 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__C1
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__C1
timestamp 1644511149
transform 1 0 25668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__C1
timestamp 1644511149
transform -1 0 27600 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A
timestamp 1644511149
transform 1 0 25852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A_N
timestamp 1644511149
transform -1 0 22448 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B
timestamp 1644511149
transform 1 0 10488 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1644511149
transform -1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__C1
timestamp 1644511149
transform -1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__C1
timestamp 1644511149
transform 1 0 16744 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B
timestamp 1644511149
transform 1 0 20976 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__C1
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__C1
timestamp 1644511149
transform -1 0 15640 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__C1
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__C1
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__C1
timestamp 1644511149
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1644511149
transform -1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1644511149
transform 1 0 7360 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1644511149
transform -1 0 5336 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A0
timestamp 1644511149
transform -1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__C1
timestamp 1644511149
transform 1 0 19964 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__C1
timestamp 1644511149
transform 1 0 21252 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A0
timestamp 1644511149
transform -1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__C1
timestamp 1644511149
transform -1 0 10856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A0
timestamp 1644511149
transform -1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__D
timestamp 1644511149
transform 1 0 25024 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__D
timestamp 1644511149
transform 1 0 26772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clock_A
timestamp 1644511149
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clock_A
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clock_A
timestamp 1644511149
transform -1 0 10488 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clock_A
timestamp 1644511149
transform -1 0 8096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clock_A
timestamp 1644511149
transform -1 0 12420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clock_A
timestamp 1644511149
transform 1 0 23828 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clock_A
timestamp 1644511149
transform -1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clock_A
timestamp 1644511149
transform 1 0 20976 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clock_A
timestamp 1644511149
transform 1 0 23644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 27876 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 27876 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 27876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 25208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 27968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 27968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 18768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 2024 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 27876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform 1 0 26496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 27876 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 16284 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 25024 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 24196 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform 1 0 3312 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 2300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 2300 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1644511149
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62
timestamp 1644511149
transform 1 0 6808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70
timestamp 1644511149
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1644511149
transform 1 0 8096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1644511149
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_188
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1644511149
transform 1 0 24840 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_262
timestamp 1644511149
transform 1 0 25208 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_268
timestamp 1644511149
transform 1 0 25760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_286
timestamp 1644511149
transform 1 0 27416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_297
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_19
timestamp 1644511149
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_31
timestamp 1644511149
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_43
timestamp 1644511149
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 1644511149
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1644511149
transform 1 0 18032 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1644511149
transform 1 0 19136 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297
timestamp 1644511149
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp 1644511149
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_6
timestamp 1644511149
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_18
timestamp 1644511149
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1644511149
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_292
timestamp 1644511149
transform 1 0 27968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp 1644511149
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_177
timestamp 1644511149
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_180
timestamp 1644511149
transform 1 0 17664 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_192
timestamp 1644511149
transform 1 0 18768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1644511149
transform 1 0 20424 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1644511149
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_234
timestamp 1644511149
transform 1 0 22632 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_246
timestamp 1644511149
transform 1 0 23736 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_258
timestamp 1644511149
transform 1 0 24840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_270
timestamp 1644511149
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1644511149
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1644511149
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_159
timestamp 1644511149
transform 1 0 15732 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_176
timestamp 1644511149
transform 1 0 17296 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1644511149
transform 1 0 20148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_227
timestamp 1644511149
transform 1 0 21988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp 1644511149
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_124
timestamp 1644511149
transform 1 0 12512 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_136
timestamp 1644511149
transform 1 0 13616 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_144
timestamp 1644511149
transform 1 0 14352 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_155
timestamp 1644511149
transform 1 0 15364 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_159
timestamp 1644511149
transform 1 0 15732 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1644511149
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_171
timestamp 1644511149
transform 1 0 16836 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_176
timestamp 1644511149
transform 1 0 17296 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_194
timestamp 1644511149
transform 1 0 18952 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_198
timestamp 1644511149
transform 1 0 19320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1644511149
transform 1 0 20240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1644511149
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_238
timestamp 1644511149
transform 1 0 23000 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_243
timestamp 1644511149
transform 1 0 23460 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_248
timestamp 1644511149
transform 1 0 23920 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_266
timestamp 1644511149
transform 1 0 25576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1644511149
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1644511149
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_157
timestamp 1644511149
transform 1 0 15548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1644511149
transform 1 0 16100 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_174
timestamp 1644511149
transform 1 0 17112 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_185
timestamp 1644511149
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_200
timestamp 1644511149
transform 1 0 19504 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_212
timestamp 1644511149
transform 1 0 20608 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_225
timestamp 1644511149
transform 1 0 21804 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_238
timestamp 1644511149
transform 1 0 23000 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1644511149
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_262
timestamp 1644511149
transform 1 0 25208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_266
timestamp 1644511149
transform 1 0 25576 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_278
timestamp 1644511149
transform 1 0 26680 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_290
timestamp 1644511149
transform 1 0 27784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1644511149
transform 1 0 28520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_102
timestamp 1644511149
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1644511149
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp 1644511149
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1644511149
transform 1 0 13616 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_147
timestamp 1644511149
transform 1 0 14628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_151
timestamp 1644511149
transform 1 0 14996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1644511149
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_173
timestamp 1644511149
transform 1 0 17020 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1644511149
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_188
timestamp 1644511149
transform 1 0 18400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_229
timestamp 1644511149
transform 1 0 22172 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_240
timestamp 1644511149
transform 1 0 23184 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_252
timestamp 1644511149
transform 1 0 24288 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_258
timestamp 1644511149
transform 1 0 24840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_268
timestamp 1644511149
transform 1 0 25760 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_291
timestamp 1644511149
transform 1 0 27876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_297
timestamp 1644511149
transform 1 0 28428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_96
timestamp 1644511149
transform 1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1644511149
transform 1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_123
timestamp 1644511149
transform 1 0 12420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_131
timestamp 1644511149
transform 1 0 13156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1644511149
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_143
timestamp 1644511149
transform 1 0 14260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_150
timestamp 1644511149
transform 1 0 14904 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_168
timestamp 1644511149
transform 1 0 16560 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_188
timestamp 1644511149
transform 1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1644511149
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_207
timestamp 1644511149
transform 1 0 20148 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_225
timestamp 1644511149
transform 1 0 21804 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1644511149
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_272
timestamp 1644511149
transform 1 0 26128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp 1644511149
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_19
timestamp 1644511149
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_31
timestamp 1644511149
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_43
timestamp 1644511149
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp 1644511149
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_95
timestamp 1644511149
transform 1 0 9844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_99
timestamp 1644511149
transform 1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1644511149
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_130
timestamp 1644511149
transform 1 0 13064 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_141
timestamp 1644511149
transform 1 0 14076 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_151
timestamp 1644511149
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_157
timestamp 1644511149
transform 1 0 15548 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1644511149
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 1644511149
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_191
timestamp 1644511149
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_197
timestamp 1644511149
transform 1 0 19228 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_208
timestamp 1644511149
transform 1 0 20240 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_213
timestamp 1644511149
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_228
timestamp 1644511149
transform 1 0 22080 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_234
timestamp 1644511149
transform 1 0 22632 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_239
timestamp 1644511149
transform 1 0 23092 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_245
timestamp 1644511149
transform 1 0 23644 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_250
timestamp 1644511149
transform 1 0 24104 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_267
timestamp 1644511149
transform 1 0 25668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_289
timestamp 1644511149
transform 1 0 27692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_292
timestamp 1644511149
transform 1 0 27968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_297
timestamp 1644511149
transform 1 0 28428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1644511149
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1644511149
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_112
timestamp 1644511149
transform 1 0 11408 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1644511149
transform 1 0 11776 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1644511149
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1644511149
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_148
timestamp 1644511149
transform 1 0 14720 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 1644511149
transform 1 0 16468 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_174
timestamp 1644511149
transform 1 0 17112 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1644511149
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_199
timestamp 1644511149
transform 1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1644511149
transform 1 0 20424 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_217
timestamp 1644511149
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_235
timestamp 1644511149
transform 1 0 22724 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1644511149
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_257
timestamp 1644511149
transform 1 0 24748 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_272
timestamp 1644511149
transform 1 0 26128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_279
timestamp 1644511149
transform 1 0 26772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_291
timestamp 1644511149
transform 1 0 27876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_84
timestamp 1644511149
transform 1 0 8832 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1644511149
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_95
timestamp 1644511149
transform 1 0 9844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1644511149
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1644511149
transform 1 0 11960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_122
timestamp 1644511149
transform 1 0 12328 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_126
timestamp 1644511149
transform 1 0 12696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_144
timestamp 1644511149
transform 1 0 14352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_148
timestamp 1644511149
transform 1 0 14720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_159
timestamp 1644511149
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1644511149
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_171
timestamp 1644511149
transform 1 0 16836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1644511149
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_179
timestamp 1644511149
transform 1 0 17572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_186
timestamp 1644511149
transform 1 0 18216 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1644511149
transform 1 0 19872 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1644511149
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_259
timestamp 1644511149
transform 1 0 24932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1644511149
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_291
timestamp 1644511149
transform 1 0 27876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 1644511149
transform 1 0 28428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_9
timestamp 1644511149
transform 1 0 1932 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_13
timestamp 1644511149
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1644511149
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp 1644511149
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_105
timestamp 1644511149
transform 1 0 10764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_125
timestamp 1644511149
transform 1 0 12604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1644511149
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1644511149
transform 1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_158
timestamp 1644511149
transform 1 0 15640 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_178
timestamp 1644511149
transform 1 0 17480 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1644511149
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_199
timestamp 1644511149
transform 1 0 19412 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_210
timestamp 1644511149
transform 1 0 20424 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_215
timestamp 1644511149
transform 1 0 20884 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_220
timestamp 1644511149
transform 1 0 21344 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_224
timestamp 1644511149
transform 1 0 21712 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_237
timestamp 1644511149
transform 1 0 22908 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_243
timestamp 1644511149
transform 1 0 23460 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1644511149
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_259
timestamp 1644511149
transform 1 0 24932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_266
timestamp 1644511149
transform 1 0 25576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_295
timestamp 1644511149
transform 1 0 28244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_89
timestamp 1644511149
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_97
timestamp 1644511149
transform 1 0 10028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_102
timestamp 1644511149
transform 1 0 10488 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1644511149
transform 1 0 10856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1644511149
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_116
timestamp 1644511149
transform 1 0 11776 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_122
timestamp 1644511149
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_127
timestamp 1644511149
transform 1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_134
timestamp 1644511149
transform 1 0 13432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1644511149
transform 1 0 14444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_152
timestamp 1644511149
transform 1 0 15088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1644511149
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_172
timestamp 1644511149
transform 1 0 16928 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_199
timestamp 1644511149
transform 1 0 19412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1644511149
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 1644511149
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_242
timestamp 1644511149
transform 1 0 23368 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_248
timestamp 1644511149
transform 1 0 23920 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_265
timestamp 1644511149
transform 1 0 25484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_269
timestamp 1644511149
transform 1 0 25852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1644511149
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_287
timestamp 1644511149
transform 1 0 27508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_292
timestamp 1644511149
transform 1 0 27968 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_298
timestamp 1644511149
transform 1 0 28520 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_6
timestamp 1644511149
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1644511149
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1644511149
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_72
timestamp 1644511149
transform 1 0 7728 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_87
timestamp 1644511149
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_92
timestamp 1644511149
transform 1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_99
timestamp 1644511149
transform 1 0 10212 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_111
timestamp 1644511149
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_123
timestamp 1644511149
transform 1 0 12420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_131
timestamp 1644511149
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1644511149
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_150
timestamp 1644511149
transform 1 0 14904 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_162
timestamp 1644511149
transform 1 0 16008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1644511149
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1644511149
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_174
timestamp 1644511149
transform 1 0 17112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_180
timestamp 1644511149
transform 1 0 17664 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_184
timestamp 1644511149
transform 1 0 18032 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1644511149
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_199
timestamp 1644511149
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_207
timestamp 1644511149
transform 1 0 20148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_211
timestamp 1644511149
transform 1 0 20516 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_228
timestamp 1644511149
transform 1 0 22080 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_232
timestamp 1644511149
transform 1 0 22448 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_237
timestamp 1644511149
transform 1 0 22908 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_246
timestamp 1644511149
transform 1 0 23736 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1644511149
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_259
timestamp 1644511149
transform 1 0 24932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_269
timestamp 1644511149
transform 1 0 25852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_286
timestamp 1644511149
transform 1 0 27416 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1644511149
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1644511149
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_63
timestamp 1644511149
transform 1 0 6900 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_68
timestamp 1644511149
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_75
timestamp 1644511149
transform 1 0 8004 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_86
timestamp 1644511149
transform 1 0 9016 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 1644511149
transform 1 0 9568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1644511149
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1644511149
transform 1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_133
timestamp 1644511149
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_141
timestamp 1644511149
transform 1 0 14076 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1644511149
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1644511149
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1644511149
transform 1 0 17204 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_187
timestamp 1644511149
transform 1 0 18308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_194
timestamp 1644511149
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1644511149
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1644511149
transform 1 0 20056 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1644511149
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_229
timestamp 1644511149
transform 1 0 22172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1644511149
transform 1 0 23092 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1644511149
transform 1 0 23460 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_256
timestamp 1644511149
transform 1 0 24656 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_262
timestamp 1644511149
transform 1 0 25208 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_270
timestamp 1644511149
transform 1 0 25944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1644511149
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1644511149
transform 1 0 6624 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_71
timestamp 1644511149
transform 1 0 7636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1644511149
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_94
timestamp 1644511149
transform 1 0 9752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_100
timestamp 1644511149
transform 1 0 10304 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_104
timestamp 1644511149
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_110
timestamp 1644511149
transform 1 0 11224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_114
timestamp 1644511149
transform 1 0 11592 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_132
timestamp 1644511149
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1644511149
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1644511149
transform 1 0 14536 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1644511149
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_161
timestamp 1644511149
transform 1 0 15916 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1644511149
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_182
timestamp 1644511149
transform 1 0 17848 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1644511149
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1644511149
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_213
timestamp 1644511149
transform 1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_220
timestamp 1644511149
transform 1 0 21344 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_230
timestamp 1644511149
transform 1 0 22264 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_240
timestamp 1644511149
transform 1 0 23184 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1644511149
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_257
timestamp 1644511149
transform 1 0 24748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_263
timestamp 1644511149
transform 1 0 25300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_271
timestamp 1644511149
transform 1 0 26036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_275
timestamp 1644511149
transform 1 0 26404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_281
timestamp 1644511149
transform 1 0 26956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_285
timestamp 1644511149
transform 1 0 27324 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_293
timestamp 1644511149
transform 1 0 28060 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1644511149
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_45
timestamp 1644511149
transform 1 0 5244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1644511149
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1644511149
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_70
timestamp 1644511149
transform 1 0 7544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_89
timestamp 1644511149
transform 1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1644511149
transform 1 0 9752 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1644511149
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_119
timestamp 1644511149
transform 1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_130
timestamp 1644511149
transform 1 0 13064 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_134
timestamp 1644511149
transform 1 0 13432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1644511149
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_154
timestamp 1644511149
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1644511149
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_179
timestamp 1644511149
transform 1 0 17572 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_187
timestamp 1644511149
transform 1 0 18308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_192
timestamp 1644511149
transform 1 0 18768 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1644511149
transform 1 0 19412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_213
timestamp 1644511149
transform 1 0 20700 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_218
timestamp 1644511149
transform 1 0 21160 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1644511149
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_228
timestamp 1644511149
transform 1 0 22080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_235
timestamp 1644511149
transform 1 0 22724 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_247
timestamp 1644511149
transform 1 0 23828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_267
timestamp 1644511149
transform 1 0 25668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_271
timestamp 1644511149
transform 1 0 26036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_297
timestamp 1644511149
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_61
timestamp 1644511149
transform 1 0 6716 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_69
timestamp 1644511149
transform 1 0 7452 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_91
timestamp 1644511149
transform 1 0 9476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_127
timestamp 1644511149
transform 1 0 12788 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1644511149
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_151
timestamp 1644511149
transform 1 0 14996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_155
timestamp 1644511149
transform 1 0 15364 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1644511149
transform 1 0 16376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_170
timestamp 1644511149
transform 1 0 16744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_185
timestamp 1644511149
transform 1 0 18124 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1644511149
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_207
timestamp 1644511149
transform 1 0 20148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_225
timestamp 1644511149
transform 1 0 21804 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1644511149
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_244
timestamp 1644511149
transform 1 0 23552 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1644511149
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_258
timestamp 1644511149
transform 1 0 24840 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_264
timestamp 1644511149
transform 1 0 25392 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_269
timestamp 1644511149
transform 1 0 25852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_276
timestamp 1644511149
transform 1 0 26496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_280
timestamp 1644511149
transform 1 0 26864 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1644511149
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_46
timestamp 1644511149
transform 1 0 5336 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1644511149
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_66
timestamp 1644511149
transform 1 0 7176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_86
timestamp 1644511149
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_97
timestamp 1644511149
transform 1 0 10028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_104
timestamp 1644511149
transform 1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1644511149
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_115
timestamp 1644511149
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_127
timestamp 1644511149
transform 1 0 12788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_153
timestamp 1644511149
transform 1 0 15180 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_178
timestamp 1644511149
transform 1 0 17480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_183
timestamp 1644511149
transform 1 0 17940 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_189
timestamp 1644511149
transform 1 0 18492 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_207
timestamp 1644511149
transform 1 0 20148 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1644511149
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_231
timestamp 1644511149
transform 1 0 22356 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_238
timestamp 1644511149
transform 1 0 23000 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_242
timestamp 1644511149
transform 1 0 23368 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_255
timestamp 1644511149
transform 1 0 24564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_263
timestamp 1644511149
transform 1 0 25300 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_269
timestamp 1644511149
transform 1 0 25852 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1644511149
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_284
timestamp 1644511149
transform 1 0 27232 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_288
timestamp 1644511149
transform 1 0 27600 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_292
timestamp 1644511149
transform 1 0 27968 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1644511149
transform 1 0 28428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_55
timestamp 1644511149
transform 1 0 6164 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_67
timestamp 1644511149
transform 1 0 7268 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_73
timestamp 1644511149
transform 1 0 7820 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1644511149
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1644511149
transform 1 0 11684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_119
timestamp 1644511149
transform 1 0 12052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_130
timestamp 1644511149
transform 1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1644511149
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1644511149
transform 1 0 14996 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1644511149
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_169
timestamp 1644511149
transform 1 0 16652 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_181
timestamp 1644511149
transform 1 0 17756 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_187
timestamp 1644511149
transform 1 0 18308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1644511149
transform 1 0 19780 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_211
timestamp 1644511149
transform 1 0 20516 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1644511149
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_219
timestamp 1644511149
transform 1 0 21252 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_230
timestamp 1644511149
transform 1 0 22264 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_237
timestamp 1644511149
transform 1 0 22908 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_246
timestamp 1644511149
transform 1 0 23736 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1644511149
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1644511149
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_267
timestamp 1644511149
transform 1 0 25668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_275
timestamp 1644511149
transform 1 0 26404 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_287
timestamp 1644511149
transform 1 0 27508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_294
timestamp 1644511149
transform 1 0 28152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_298
timestamp 1644511149
transform 1 0 28520 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_43
timestamp 1644511149
transform 1 0 5060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_46
timestamp 1644511149
transform 1 0 5336 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1644511149
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_66
timestamp 1644511149
transform 1 0 7176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_79
timestamp 1644511149
transform 1 0 8372 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_87
timestamp 1644511149
transform 1 0 9108 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_99
timestamp 1644511149
transform 1 0 10212 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_104
timestamp 1644511149
transform 1 0 10672 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1644511149
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1644511149
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp 1644511149
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1644511149
transform 1 0 13156 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_141
timestamp 1644511149
transform 1 0 14076 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1644511149
transform 1 0 14996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1644511149
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_171
timestamp 1644511149
transform 1 0 16836 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_182
timestamp 1644511149
transform 1 0 17848 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_186
timestamp 1644511149
transform 1 0 18216 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_204
timestamp 1644511149
transform 1 0 19872 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_211
timestamp 1644511149
transform 1 0 20516 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1644511149
transform 1 0 20884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1644511149
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_230
timestamp 1644511149
transform 1 0 22264 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_235
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1644511149
transform 1 0 24472 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_297
timestamp 1644511149
transform 1 0 28428 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_60
timestamp 1644511149
transform 1 0 6624 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1644511149
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1644511149
transform 1 0 9200 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_92
timestamp 1644511149
transform 1 0 9568 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_116
timestamp 1644511149
transform 1 0 11776 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_126
timestamp 1644511149
transform 1 0 12696 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1644511149
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1644511149
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1644511149
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_172
timestamp 1644511149
transform 1 0 16928 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_188
timestamp 1644511149
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1644511149
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_201
timestamp 1644511149
transform 1 0 19596 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_230
timestamp 1644511149
transform 1 0 22264 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_242
timestamp 1644511149
transform 1 0 23368 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1644511149
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_260
timestamp 1644511149
transform 1 0 25024 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_264
timestamp 1644511149
transform 1 0 25392 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_270
timestamp 1644511149
transform 1 0 25944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_281
timestamp 1644511149
transform 1 0 26956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_287
timestamp 1644511149
transform 1 0 27508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1644511149
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_6
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_18
timestamp 1644511149
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_30
timestamp 1644511149
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_42
timestamp 1644511149
transform 1 0 4968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_46
timestamp 1644511149
transform 1 0 5336 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1644511149
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_65
timestamp 1644511149
transform 1 0 7084 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_73
timestamp 1644511149
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_80
timestamp 1644511149
transform 1 0 8464 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_89
timestamp 1644511149
transform 1 0 9292 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_100
timestamp 1644511149
transform 1 0 10304 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_106
timestamp 1644511149
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1644511149
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_129
timestamp 1644511149
transform 1 0 12972 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1644511149
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1644511149
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_178
timestamp 1644511149
transform 1 0 17480 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_185
timestamp 1644511149
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_191
timestamp 1644511149
transform 1 0 18676 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_196
timestamp 1644511149
transform 1 0 19136 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1644511149
transform 1 0 19872 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_208
timestamp 1644511149
transform 1 0 20240 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_216
timestamp 1644511149
transform 1 0 20976 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1644511149
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_241
timestamp 1644511149
transform 1 0 23276 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_247
timestamp 1644511149
transform 1 0 23828 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_265
timestamp 1644511149
transform 1 0 25484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1644511149
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_297
timestamp 1644511149
transform 1 0 28428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1644511149
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_49
timestamp 1644511149
transform 1 0 5612 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_66
timestamp 1644511149
transform 1 0 7176 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_72
timestamp 1644511149
transform 1 0 7728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1644511149
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_88
timestamp 1644511149
transform 1 0 9200 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_112
timestamp 1644511149
transform 1 0 11408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_122
timestamp 1644511149
transform 1 0 12328 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_128
timestamp 1644511149
transform 1 0 12880 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1644511149
transform 1 0 14812 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_171
timestamp 1644511149
transform 1 0 16836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1644511149
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_201
timestamp 1644511149
transform 1 0 19596 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_210
timestamp 1644511149
transform 1 0 20424 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_222
timestamp 1644511149
transform 1 0 21528 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_228
timestamp 1644511149
transform 1 0 22080 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_240
timestamp 1644511149
transform 1 0 23184 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_256
timestamp 1644511149
transform 1 0 24656 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_269
timestamp 1644511149
transform 1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_276
timestamp 1644511149
transform 1 0 26496 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_296
timestamp 1644511149
transform 1 0 28336 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1644511149
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1644511149
transform 1 0 6808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_73
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_95
timestamp 1644511149
transform 1 0 9844 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_103
timestamp 1644511149
transform 1 0 10580 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1644511149
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_126
timestamp 1644511149
transform 1 0 12696 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_134
timestamp 1644511149
transform 1 0 13432 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1644511149
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_148
timestamp 1644511149
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_158
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1644511149
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_178
timestamp 1644511149
transform 1 0 17480 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_185
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_189
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_201
timestamp 1644511149
transform 1 0 19596 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1644511149
transform 1 0 20516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1644511149
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_235
timestamp 1644511149
transform 1 0 22724 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_244
timestamp 1644511149
transform 1 0 23552 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_252
timestamp 1644511149
transform 1 0 24288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_267
timestamp 1644511149
transform 1 0 25668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1644511149
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_287
timestamp 1644511149
transform 1 0 27508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_291
timestamp 1644511149
transform 1 0 27876 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1644511149
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_6
timestamp 1644511149
transform 1 0 1656 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp 1644511149
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1644511149
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_61
timestamp 1644511149
transform 1 0 6716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1644511149
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_76
timestamp 1644511149
transform 1 0 8096 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1644511149
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_101
timestamp 1644511149
transform 1 0 10396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_107
timestamp 1644511149
transform 1 0 10948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_119
timestamp 1644511149
transform 1 0 12052 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_131
timestamp 1644511149
transform 1 0 13156 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1644511149
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_149
timestamp 1644511149
transform 1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_158
timestamp 1644511149
transform 1 0 15640 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_166
timestamp 1644511149
transform 1 0 16376 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_172
timestamp 1644511149
transform 1 0 16928 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1644511149
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1644511149
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_207
timestamp 1644511149
transform 1 0 20148 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_216
timestamp 1644511149
transform 1 0 20976 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_225
timestamp 1644511149
transform 1 0 21804 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_230
timestamp 1644511149
transform 1 0 22264 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_241
timestamp 1644511149
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1644511149
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_260
timestamp 1644511149
transform 1 0 25024 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_266
timestamp 1644511149
transform 1 0 25576 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_272
timestamp 1644511149
transform 1 0 26128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1644511149
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_19
timestamp 1644511149
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 1644511149
transform 1 0 8096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_87
timestamp 1644511149
transform 1 0 9108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_92
timestamp 1644511149
transform 1 0 9568 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1644511149
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_121
timestamp 1644511149
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_131
timestamp 1644511149
transform 1 0 13156 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_139
timestamp 1644511149
transform 1 0 13892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1644511149
transform 1 0 15732 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1644511149
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_173
timestamp 1644511149
transform 1 0 17020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1644511149
transform 1 0 18032 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_188
timestamp 1644511149
transform 1 0 18400 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_192
timestamp 1644511149
transform 1 0 18768 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_196
timestamp 1644511149
transform 1 0 19136 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_204
timestamp 1644511149
transform 1 0 19872 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_214
timestamp 1644511149
transform 1 0 20792 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_238
timestamp 1644511149
transform 1 0 23000 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_244
timestamp 1644511149
transform 1 0 23552 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_258
timestamp 1644511149
transform 1 0 24840 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1644511149
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_284
timestamp 1644511149
transform 1 0 27232 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_292
timestamp 1644511149
transform 1 0 27968 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_297
timestamp 1644511149
transform 1 0 28428 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_61
timestamp 1644511149
transform 1 0 6716 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_66
timestamp 1644511149
transform 1 0 7176 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_72
timestamp 1644511149
transform 1 0 7728 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_101
timestamp 1644511149
transform 1 0 10396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_118
timestamp 1644511149
transform 1 0 11960 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1644511149
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_147
timestamp 1644511149
transform 1 0 14628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_154
timestamp 1644511149
transform 1 0 15272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_160
timestamp 1644511149
transform 1 0 15824 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_171
timestamp 1644511149
transform 1 0 16836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1644511149
transform 1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1644511149
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_203
timestamp 1644511149
transform 1 0 19780 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_216
timestamp 1644511149
transform 1 0 20976 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_224
timestamp 1644511149
transform 1 0 21712 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_232
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1644511149
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_271
timestamp 1644511149
transform 1 0 26036 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_282
timestamp 1644511149
transform 1 0 27048 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_288
timestamp 1644511149
transform 1 0 27600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_295
timestamp 1644511149
transform 1 0 28244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_73
timestamp 1644511149
transform 1 0 7820 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_76
timestamp 1644511149
transform 1 0 8096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_82
timestamp 1644511149
transform 1 0 8648 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_89
timestamp 1644511149
transform 1 0 9292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_102
timestamp 1644511149
transform 1 0 10488 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1644511149
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1644511149
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_122
timestamp 1644511149
transform 1 0 12328 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_128
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_133
timestamp 1644511149
transform 1 0 13340 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_140
timestamp 1644511149
transform 1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_147
timestamp 1644511149
transform 1 0 14628 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1644511149
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1644511149
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_172
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1644511149
transform 1 0 17572 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_183
timestamp 1644511149
transform 1 0 17940 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_188
timestamp 1644511149
transform 1 0 18400 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1644511149
transform 1 0 19044 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1644511149
transform 1 0 19780 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1644511149
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1644511149
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_228
timestamp 1644511149
transform 1 0 22080 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_241
timestamp 1644511149
transform 1 0 23276 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_245
timestamp 1644511149
transform 1 0 23644 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_252
timestamp 1644511149
transform 1 0 24288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_258
timestamp 1644511149
transform 1 0 24840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_267
timestamp 1644511149
transform 1 0 25668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_271
timestamp 1644511149
transform 1 0 26036 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1644511149
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_297
timestamp 1644511149
transform 1 0 28428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1644511149
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_101
timestamp 1644511149
transform 1 0 10396 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_114
timestamp 1644511149
transform 1 0 11592 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_124
timestamp 1644511149
transform 1 0 12512 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_128
timestamp 1644511149
transform 1 0 12880 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1644511149
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1644511149
transform 1 0 14996 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_161
timestamp 1644511149
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_182
timestamp 1644511149
transform 1 0 17848 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_186
timestamp 1644511149
transform 1 0 18216 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1644511149
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_214
timestamp 1644511149
transform 1 0 20792 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1644511149
transform 1 0 21160 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_225
timestamp 1644511149
transform 1 0 21804 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_232
timestamp 1644511149
transform 1 0 22448 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_236
timestamp 1644511149
transform 1 0 22816 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_244
timestamp 1644511149
transform 1 0 23552 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1644511149
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_261
timestamp 1644511149
transform 1 0 25116 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_266
timestamp 1644511149
transform 1 0 25576 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_274
timestamp 1644511149
transform 1 0 26312 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_280
timestamp 1644511149
transform 1 0 26864 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_292
timestamp 1644511149
transform 1 0 27968 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1644511149
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_92
timestamp 1644511149
transform 1 0 9568 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_104
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_129
timestamp 1644511149
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_136
timestamp 1644511149
transform 1 0 13616 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_154
timestamp 1644511149
transform 1 0 15272 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1644511149
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1644511149
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_182
timestamp 1644511149
transform 1 0 17848 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_189
timestamp 1644511149
transform 1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_198
timestamp 1644511149
transform 1 0 19320 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1644511149
transform 1 0 19872 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1644511149
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_243
timestamp 1644511149
transform 1 0 23460 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_247
timestamp 1644511149
transform 1 0 23828 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_259
timestamp 1644511149
transform 1 0 24932 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1644511149
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_271
timestamp 1644511149
transform 1 0 26036 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1644511149
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 1644511149
transform 1 0 28428 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_115
timestamp 1644511149
transform 1 0 11684 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_118
timestamp 1644511149
transform 1 0 11960 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_128
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_156
timestamp 1644511149
transform 1 0 15456 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_164
timestamp 1644511149
transform 1 0 16192 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_168
timestamp 1644511149
transform 1 0 16560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_172
timestamp 1644511149
transform 1 0 16928 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_176
timestamp 1644511149
transform 1 0 17296 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1644511149
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_203
timestamp 1644511149
transform 1 0 19780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_207
timestamp 1644511149
transform 1 0 20148 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_217
timestamp 1644511149
transform 1 0 21068 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_231
timestamp 1644511149
transform 1 0 22356 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_237
timestamp 1644511149
transform 1 0 22908 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_243
timestamp 1644511149
transform 1 0 23460 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1644511149
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_259
timestamp 1644511149
transform 1 0 24932 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1644511149
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_273
timestamp 1644511149
transform 1 0 26220 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_279
timestamp 1644511149
transform 1 0 26772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp 1644511149
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_146
timestamp 1644511149
transform 1 0 14536 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1644511149
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_177
timestamp 1644511149
transform 1 0 17388 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1644511149
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1644511149
transform 1 0 19872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_208
timestamp 1644511149
transform 1 0 20240 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_241
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_250
timestamp 1644511149
transform 1 0 24104 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_257
timestamp 1644511149
transform 1 0 24748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_262
timestamp 1644511149
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_268
timestamp 1644511149
transform 1 0 25760 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_272
timestamp 1644511149
transform 1 0 26128 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_297
timestamp 1644511149
transform 1 0 28428 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_6
timestamp 1644511149
transform 1 0 1656 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_18
timestamp 1644511149
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1644511149
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_129
timestamp 1644511149
transform 1 0 12972 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1644511149
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_146
timestamp 1644511149
transform 1 0 14536 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_150
timestamp 1644511149
transform 1 0 14904 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_161
timestamp 1644511149
transform 1 0 15916 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_176
timestamp 1644511149
transform 1 0 17296 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_185
timestamp 1644511149
transform 1 0 18124 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1644511149
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_208
timestamp 1644511149
transform 1 0 20240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_238
timestamp 1644511149
transform 1 0 23000 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1644511149
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_261
timestamp 1644511149
transform 1 0 25116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_267
timestamp 1644511149
transform 1 0 25668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_285
timestamp 1644511149
transform 1 0 27324 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_293
timestamp 1644511149
transform 1 0 28060 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp 1644511149
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_123
timestamp 1644511149
transform 1 0 12420 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_147
timestamp 1644511149
transform 1 0 14628 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1644511149
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_179
timestamp 1644511149
transform 1 0 17572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_191
timestamp 1644511149
transform 1 0 18676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_204
timestamp 1644511149
transform 1 0 19872 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_212
timestamp 1644511149
transform 1 0 20608 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_242
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_254
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1644511149
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_263
timestamp 1644511149
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_268
timestamp 1644511149
transform 1 0 25760 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 1644511149
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_297
timestamp 1644511149
transform 1 0 28428 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_127
timestamp 1644511149
transform 1 0 12788 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1644511149
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_38_150
timestamp 1644511149
transform 1 0 14904 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_156
timestamp 1644511149
transform 1 0 15456 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_174
timestamp 1644511149
transform 1 0 17112 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_182
timestamp 1644511149
transform 1 0 17848 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_190
timestamp 1644511149
transform 1 0 18584 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1644511149
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_208
timestamp 1644511149
transform 1 0 20240 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_214
timestamp 1644511149
transform 1 0 20792 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_218
timestamp 1644511149
transform 1 0 21160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_222
timestamp 1644511149
transform 1 0 21528 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_227
timestamp 1644511149
transform 1 0 21988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_232
timestamp 1644511149
transform 1 0 22448 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_240
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1644511149
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_257
timestamp 1644511149
transform 1 0 24748 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_262
timestamp 1644511149
transform 1 0 25208 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_272
timestamp 1644511149
transform 1 0 26128 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp 1644511149
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_6
timestamp 1644511149
transform 1 0 1656 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_18
timestamp 1644511149
transform 1 0 2760 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_30
timestamp 1644511149
transform 1 0 3864 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_42
timestamp 1644511149
transform 1 0 4968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1644511149
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_153
timestamp 1644511149
transform 1 0 15180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_163
timestamp 1644511149
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1644511149
transform 1 0 17572 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_183
timestamp 1644511149
transform 1 0 17940 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_201
timestamp 1644511149
transform 1 0 19596 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_206
timestamp 1644511149
transform 1 0 20056 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_212
timestamp 1644511149
transform 1 0 20608 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1644511149
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_235
timestamp 1644511149
transform 1 0 22724 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_243
timestamp 1644511149
transform 1 0 23460 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_252
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_259
timestamp 1644511149
transform 1 0 24932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1644511149
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_291
timestamp 1644511149
transform 1 0 27876 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_297
timestamp 1644511149
transform 1 0 28428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1644511149
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_147
timestamp 1644511149
transform 1 0 14628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_154
timestamp 1644511149
transform 1 0 15272 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_158
timestamp 1644511149
transform 1 0 15640 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_186
timestamp 1644511149
transform 1 0 18216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1644511149
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_220
timestamp 1644511149
transform 1 0 21344 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_224
timestamp 1644511149
transform 1 0 21712 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1644511149
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1644511149
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_260
timestamp 1644511149
transform 1 0 25024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_269
timestamp 1644511149
transform 1 0 25852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_274
timestamp 1644511149
transform 1 0 26312 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_286
timestamp 1644511149
transform 1 0 27416 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_298
timestamp 1644511149
transform 1 0 28520 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_155
timestamp 1644511149
transform 1 0 15364 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_159
timestamp 1644511149
transform 1 0 15732 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_165
timestamp 1644511149
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_176
timestamp 1644511149
transform 1 0 17296 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_180
timestamp 1644511149
transform 1 0 17664 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_191
timestamp 1644511149
transform 1 0 18676 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_197
timestamp 1644511149
transform 1 0 19228 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_207
timestamp 1644511149
transform 1 0 20148 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_213
timestamp 1644511149
transform 1 0 20700 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1644511149
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_230
timestamp 1644511149
transform 1 0 22264 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_235
timestamp 1644511149
transform 1 0 22724 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1644511149
transform 1 0 23092 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1644511149
transform 1 0 23460 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_247
timestamp 1644511149
transform 1 0 23828 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_266
timestamp 1644511149
transform 1 0 25576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1644511149
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_291
timestamp 1644511149
transform 1 0 27876 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_297
timestamp 1644511149
transform 1 0 28428 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_171
timestamp 1644511149
transform 1 0 16836 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_179
timestamp 1644511149
transform 1 0 17572 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1644511149
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_203
timestamp 1644511149
transform 1 0 19780 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_207
timestamp 1644511149
transform 1 0 20148 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_215
timestamp 1644511149
transform 1 0 20884 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_225
timestamp 1644511149
transform 1 0 21804 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_243
timestamp 1644511149
transform 1 0 23460 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1644511149
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_262
timestamp 1644511149
transform 1 0 25208 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_284
timestamp 1644511149
transform 1 0 27232 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_296
timestamp 1644511149
transform 1 0 28336 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_153
timestamp 1644511149
transform 1 0 15180 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_157
timestamp 1644511149
transform 1 0 15548 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_163
timestamp 1644511149
transform 1 0 16100 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1644511149
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_177
timestamp 1644511149
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_182
timestamp 1644511149
transform 1 0 17848 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_186
timestamp 1644511149
transform 1 0 18216 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_194
timestamp 1644511149
transform 1 0 18952 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_202
timestamp 1644511149
transform 1 0 19688 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_208
timestamp 1644511149
transform 1 0 20240 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_231
timestamp 1644511149
transform 1 0 22356 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_236
timestamp 1644511149
transform 1 0 22816 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_242
timestamp 1644511149
transform 1 0 23368 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_259
timestamp 1644511149
transform 1 0 24932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_263
timestamp 1644511149
transform 1 0 25300 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_271
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_9
timestamp 1644511149
transform 1 0 1932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_13
timestamp 1644511149
transform 1 0 2300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1644511149
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_161
timestamp 1644511149
transform 1 0 15916 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_179
timestamp 1644511149
transform 1 0 17572 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_183
timestamp 1644511149
transform 1 0 17940 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_204
timestamp 1644511149
transform 1 0 19872 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_211
timestamp 1644511149
transform 1 0 20516 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_215
timestamp 1644511149
transform 1 0 20884 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_222
timestamp 1644511149
transform 1 0 21528 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_229
timestamp 1644511149
transform 1 0 22172 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_241
timestamp 1644511149
transform 1 0 23276 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1644511149
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_259
timestamp 1644511149
transform 1 0 24932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_262
timestamp 1644511149
transform 1 0 25208 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_274
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_278
timestamp 1644511149
transform 1 0 26680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_281
timestamp 1644511149
transform 1 0 26956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp 1644511149
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_6
timestamp 1644511149
transform 1 0 1656 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_10
timestamp 1644511149
transform 1 0 2024 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_22
timestamp 1644511149
transform 1 0 3128 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_34
timestamp 1644511149
transform 1 0 4232 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_46
timestamp 1644511149
transform 1 0 5336 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1644511149
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_131
timestamp 1644511149
transform 1 0 13156 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_148
timestamp 1644511149
transform 1 0 14720 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1644511149
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_177
timestamp 1644511149
transform 1 0 17388 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_194
timestamp 1644511149
transform 1 0 18952 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_212
timestamp 1644511149
transform 1 0 20608 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1644511149
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_241
timestamp 1644511149
transform 1 0 23276 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_251
timestamp 1644511149
transform 1 0 24196 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_259
timestamp 1644511149
transform 1 0 24932 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1644511149
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_297
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_7
timestamp 1644511149
transform 1 0 1748 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_13
timestamp 1644511149
transform 1 0 2300 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_21
timestamp 1644511149
transform 1 0 3036 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1644511149
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_37
timestamp 1644511149
transform 1 0 4508 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_49
timestamp 1644511149
transform 1 0 5612 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_55
timestamp 1644511149
transform 1 0 6164 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_60
timestamp 1644511149
transform 1 0 6624 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_72
timestamp 1644511149
transform 1 0 7728 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_113
timestamp 1644511149
transform 1 0 11500 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_125
timestamp 1644511149
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1644511149
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_145
timestamp 1644511149
transform 1 0 14444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_149
timestamp 1644511149
transform 1 0 14812 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_154
timestamp 1644511149
transform 1 0 15272 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_166
timestamp 1644511149
transform 1 0 16376 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_173
timestamp 1644511149
transform 1 0 17020 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_181
timestamp 1644511149
transform 1 0 17756 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1644511149
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1644511149
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_200
timestamp 1644511149
transform 1 0 19504 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_207
timestamp 1644511149
transform 1 0 20148 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_212
timestamp 1644511149
transform 1 0 20608 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_228
timestamp 1644511149
transform 1 0 22080 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_240
timestamp 1644511149
transform 1 0 23184 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_257
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_260
timestamp 1644511149
transform 1 0 25024 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_268
timestamp 1644511149
transform 1 0 25760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_278
timestamp 1644511149
transform 1 0 26680 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_281
timestamp 1644511149
transform 1 0 26956 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0522_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0523_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 14996 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0524_
timestamp 1644511149
transform 1 0 14168 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0525_
timestamp 1644511149
transform 1 0 15272 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_1  _0526_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24656 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0527_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22908 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0528_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0529_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0530_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0531_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28152 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0532_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0533_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24656 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0534_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25024 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0535_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23644 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0536_
timestamp 1644511149
transform -1 0 27508 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0537_
timestamp 1644511149
transform -1 0 25668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0538_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0539_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0540_
timestamp 1644511149
transform 1 0 24932 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0541_
timestamp 1644511149
transform -1 0 25116 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0542_
timestamp 1644511149
transform 1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0543_
timestamp 1644511149
transform -1 0 23092 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0544_
timestamp 1644511149
transform 1 0 22356 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0545_
timestamp 1644511149
transform -1 0 23644 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0546_
timestamp 1644511149
transform 1 0 22172 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0547_
timestamp 1644511149
transform -1 0 22172 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0548_
timestamp 1644511149
transform 1 0 22172 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0549_
timestamp 1644511149
transform -1 0 22632 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0550_
timestamp 1644511149
transform -1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0551_
timestamp 1644511149
transform 1 0 20976 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0552_
timestamp 1644511149
transform 1 0 20424 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1644511149
transform -1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0554_
timestamp 1644511149
transform 1 0 19412 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0555_
timestamp 1644511149
transform 1 0 19320 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0556_
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0557_
timestamp 1644511149
transform -1 0 20148 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0558_
timestamp 1644511149
transform 1 0 19412 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 1644511149
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0560_
timestamp 1644511149
transform -1 0 22908 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0561_
timestamp 1644511149
transform 1 0 22080 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0562_
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0563_
timestamp 1644511149
transform 1 0 23276 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0564_
timestamp 1644511149
transform 1 0 23552 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0565_
timestamp 1644511149
transform -1 0 24104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21528 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0567_
timestamp 1644511149
transform 1 0 22080 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0568_
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0569_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23736 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1644511149
transform -1 0 17940 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0571_
timestamp 1644511149
transform -1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0572_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0573_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20976 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0574_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0575_
timestamp 1644511149
transform 1 0 12144 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0576_
timestamp 1644511149
transform 1 0 22356 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0577_
timestamp 1644511149
transform -1 0 23184 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0578_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22264 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0579_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20884 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1644511149
transform 1 0 20792 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0581_
timestamp 1644511149
transform -1 0 18492 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0582_
timestamp 1644511149
transform 1 0 23552 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0583_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0584_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0585_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0586_
timestamp 1644511149
transform -1 0 25852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0587_
timestamp 1644511149
transform -1 0 25484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0588_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0589_
timestamp 1644511149
transform 1 0 17572 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0590_
timestamp 1644511149
transform 1 0 17388 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _0591_
timestamp 1644511149
transform 1 0 18032 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _0592_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0593_
timestamp 1644511149
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0594_
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0595_
timestamp 1644511149
transform 1 0 17848 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0596_
timestamp 1644511149
transform 1 0 18216 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0597_
timestamp 1644511149
transform -1 0 19228 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0598_
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0599_
timestamp 1644511149
transform 1 0 23552 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1644511149
transform -1 0 23920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0601_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0602_
timestamp 1644511149
transform -1 0 20424 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0603_
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0604_
timestamp 1644511149
transform 1 0 20424 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 1644511149
transform 1 0 17664 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0606_
timestamp 1644511149
transform -1 0 18124 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0607_
timestamp 1644511149
transform -1 0 17296 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0608_
timestamp 1644511149
transform 1 0 19596 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0609_
timestamp 1644511149
transform 1 0 19688 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0610_
timestamp 1644511149
transform 1 0 20608 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0611_
timestamp 1644511149
transform -1 0 12788 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0612_
timestamp 1644511149
transform 1 0 9936 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0614_
timestamp 1644511149
transform -1 0 16376 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1644511149
transform -1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0616_
timestamp 1644511149
transform 1 0 17204 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0617_
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1644511149
transform -1 0 17020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0619_
timestamp 1644511149
transform 1 0 19044 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0620_
timestamp 1644511149
transform -1 0 18860 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1644511149
transform -1 0 21344 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1644511149
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0623_
timestamp 1644511149
transform 1 0 16652 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1644511149
transform -1 0 17572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0625_
timestamp 1644511149
transform -1 0 11224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1644511149
transform 1 0 8188 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1644511149
transform 1 0 8004 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0628_
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0629_
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0630_
timestamp 1644511149
transform -1 0 8372 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 1644511149
transform -1 0 8004 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0632_
timestamp 1644511149
transform -1 0 10028 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0633_
timestamp 1644511149
transform -1 0 10672 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1644511149
transform 1 0 7636 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0635_
timestamp 1644511149
transform 1 0 7360 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1644511149
transform 1 0 8004 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0637_
timestamp 1644511149
transform 1 0 9200 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0638_
timestamp 1644511149
transform 1 0 9200 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1644511149
transform -1 0 10212 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0640_
timestamp 1644511149
transform 1 0 7544 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0641_
timestamp 1644511149
transform 1 0 7360 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0643_
timestamp 1644511149
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0644_
timestamp 1644511149
transform 1 0 8004 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0646_
timestamp 1644511149
transform 1 0 9476 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0647_
timestamp 1644511149
transform 1 0 8832 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1644511149
transform 1 0 10396 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0649_
timestamp 1644511149
transform 1 0 9476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0650_
timestamp 1644511149
transform 1 0 9936 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0651_
timestamp 1644511149
transform 1 0 9016 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0652_
timestamp 1644511149
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1644511149
transform -1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0654_
timestamp 1644511149
transform -1 0 17664 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0655_
timestamp 1644511149
transform -1 0 18768 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0656_
timestamp 1644511149
transform -1 0 16928 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0657_
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0658_
timestamp 1644511149
transform 1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0659_
timestamp 1644511149
transform -1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0660_
timestamp 1644511149
transform -1 0 17388 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0661_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16100 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1644511149
transform 1 0 12420 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0663_
timestamp 1644511149
transform 1 0 13616 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0664_
timestamp 1644511149
transform -1 0 12236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0665_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11960 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0666_
timestamp 1644511149
transform 1 0 12420 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0667_
timestamp 1644511149
transform -1 0 13156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0668_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0669_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0670_
timestamp 1644511149
transform 1 0 11316 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0671_
timestamp 1644511149
transform 1 0 11592 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0672_
timestamp 1644511149
transform -1 0 11224 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0673_
timestamp 1644511149
transform -1 0 12052 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0674_
timestamp 1644511149
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0675_
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0676_
timestamp 1644511149
transform -1 0 13616 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0677_
timestamp 1644511149
transform 1 0 11776 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0678_
timestamp 1644511149
transform -1 0 12972 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0679_
timestamp 1644511149
transform 1 0 12144 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0680_
timestamp 1644511149
transform -1 0 15456 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0681_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0682_
timestamp 1644511149
transform 1 0 18032 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 1644511149
transform 1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0684_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17388 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _0685_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_2  _0686_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0687_
timestamp 1644511149
transform -1 0 14536 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0688_
timestamp 1644511149
transform -1 0 13156 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0689_
timestamp 1644511149
transform 1 0 10028 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1644511149
transform -1 0 10028 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 1644511149
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1644511149
transform 1 0 10488 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0693_
timestamp 1644511149
transform -1 0 10212 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0694_
timestamp 1644511149
transform -1 0 9568 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0695_
timestamp 1644511149
transform 1 0 10580 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0696_
timestamp 1644511149
transform -1 0 9844 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1644511149
transform -1 0 8648 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 1644511149
transform 1 0 10396 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0699_
timestamp 1644511149
transform -1 0 10488 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 1644511149
transform -1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0701_
timestamp 1644511149
transform -1 0 12420 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 1644511149
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0703_
timestamp 1644511149
transform -1 0 11960 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0704_
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1644511149
transform 1 0 12420 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0706_
timestamp 1644511149
transform 1 0 11776 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1644511149
transform 1 0 12512 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0708_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18492 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 1644511149
transform 1 0 17664 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0710_
timestamp 1644511149
transform -1 0 17756 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0711_
timestamp 1644511149
transform -1 0 18952 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0712_
timestamp 1644511149
transform 1 0 15180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0713_
timestamp 1644511149
transform 1 0 15272 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0714_
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0715_
timestamp 1644511149
transform -1 0 16928 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0716_
timestamp 1644511149
transform -1 0 15732 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1644511149
transform -1 0 16376 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0718_
timestamp 1644511149
transform -1 0 13800 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 1644511149
transform 1 0 13616 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0720_
timestamp 1644511149
transform 1 0 12972 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0721_
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0722_
timestamp 1644511149
transform 1 0 10856 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 1644511149
transform 1 0 13800 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0724_
timestamp 1644511149
transform 1 0 13156 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0725_
timestamp 1644511149
transform -1 0 13800 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0726_
timestamp 1644511149
transform 1 0 15088 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0727_
timestamp 1644511149
transform 1 0 14444 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0728_
timestamp 1644511149
transform -1 0 16376 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0729_
timestamp 1644511149
transform 1 0 12512 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0730_
timestamp 1644511149
transform -1 0 12420 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0731_
timestamp 1644511149
transform 1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1644511149
transform 1 0 13248 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0733_
timestamp 1644511149
transform 1 0 12144 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0734_
timestamp 1644511149
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0735_
timestamp 1644511149
transform 1 0 19412 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0736_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17480 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _0737_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17020 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0738_
timestamp 1644511149
transform 1 0 18308 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0739_
timestamp 1644511149
transform -1 0 17480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0740_
timestamp 1644511149
transform 1 0 17664 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0741_
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0742_
timestamp 1644511149
transform -1 0 15824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0743_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0745_
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0746_
timestamp 1644511149
transform -1 0 17296 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0747_
timestamp 1644511149
transform 1 0 19412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1644511149
transform 1 0 17204 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0749_
timestamp 1644511149
transform -1 0 17572 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0750_
timestamp 1644511149
transform -1 0 16928 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0751_
timestamp 1644511149
transform 1 0 17572 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0752_
timestamp 1644511149
transform 1 0 17848 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 1644511149
transform 1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0754_
timestamp 1644511149
transform -1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0755_
timestamp 1644511149
transform 1 0 16008 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0756_
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0757_
timestamp 1644511149
transform 1 0 17020 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1644511149
transform -1 0 19320 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0759_
timestamp 1644511149
transform -1 0 19044 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0760_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18952 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0761_
timestamp 1644511149
transform 1 0 19412 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0762_
timestamp 1644511149
transform -1 0 17848 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0763_
timestamp 1644511149
transform -1 0 18492 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0764_
timestamp 1644511149
transform 1 0 17572 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0765_
timestamp 1644511149
transform -1 0 16376 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0766_
timestamp 1644511149
transform -1 0 16192 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0767_
timestamp 1644511149
transform 1 0 15640 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0768_
timestamp 1644511149
transform 1 0 18952 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0769_
timestamp 1644511149
transform -1 0 27324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp 1644511149
transform 1 0 25760 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0771_
timestamp 1644511149
transform 1 0 25944 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0772_
timestamp 1644511149
transform 1 0 27692 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0773_
timestamp 1644511149
transform -1 0 25668 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0774_
timestamp 1644511149
transform 1 0 24288 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0775_
timestamp 1644511149
transform -1 0 28244 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0776_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24932 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0777_
timestamp 1644511149
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _0778_
timestamp 1644511149
transform -1 0 25024 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0779_
timestamp 1644511149
transform -1 0 21528 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0780_
timestamp 1644511149
transform -1 0 22264 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0781_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0782_
timestamp 1644511149
transform 1 0 16928 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0783_
timestamp 1644511149
transform 1 0 17940 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0784_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20240 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1644511149
transform 1 0 19780 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0786_
timestamp 1644511149
transform 1 0 16652 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0787_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19044 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0788_
timestamp 1644511149
transform 1 0 17480 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _0789_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18216 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0790_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0791_
timestamp 1644511149
transform -1 0 25760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0792_
timestamp 1644511149
transform -1 0 23460 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0793_
timestamp 1644511149
transform -1 0 21068 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0794_
timestamp 1644511149
transform -1 0 22080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1644511149
transform -1 0 22724 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0796_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21068 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0797_
timestamp 1644511149
transform 1 0 20332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0798_
timestamp 1644511149
transform 1 0 19964 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0799_
timestamp 1644511149
transform 1 0 20700 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0800_
timestamp 1644511149
transform 1 0 19412 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0801_
timestamp 1644511149
transform 1 0 20056 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0802_
timestamp 1644511149
transform -1 0 23000 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0803_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21528 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0804_
timestamp 1644511149
transform -1 0 19596 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0805_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0806_
timestamp 1644511149
transform -1 0 21528 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0807_
timestamp 1644511149
transform 1 0 19780 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0808_
timestamp 1644511149
transform -1 0 22264 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0809_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0810_
timestamp 1644511149
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0811_
timestamp 1644511149
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0812_
timestamp 1644511149
transform 1 0 19228 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0813_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19044 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0814_
timestamp 1644511149
transform 1 0 20516 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0815_
timestamp 1644511149
transform 1 0 21620 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0816_
timestamp 1644511149
transform -1 0 22080 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0817_
timestamp 1644511149
transform 1 0 23736 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0818_
timestamp 1644511149
transform -1 0 24012 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0819_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0820_
timestamp 1644511149
transform -1 0 21528 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0821_
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0822_
timestamp 1644511149
transform 1 0 25300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0823_
timestamp 1644511149
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1644511149
transform 1 0 21988 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0825_
timestamp 1644511149
transform 1 0 21160 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0826_
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0827_
timestamp 1644511149
transform 1 0 24748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0828_
timestamp 1644511149
transform 1 0 25300 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a221oi_1  _0829_
timestamp 1644511149
transform -1 0 23736 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0830_
timestamp 1644511149
transform -1 0 25484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0831_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 20976 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0832_
timestamp 1644511149
transform 1 0 20148 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0833_
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0834_
timestamp 1644511149
transform -1 0 25024 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0835_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0836_
timestamp 1644511149
transform -1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0837_
timestamp 1644511149
transform 1 0 22080 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0838_
timestamp 1644511149
transform 1 0 27140 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0839_
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _0840_
timestamp 1644511149
transform -1 0 26312 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0841_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22816 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0842_
timestamp 1644511149
transform 1 0 26312 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0843_
timestamp 1644511149
transform -1 0 19596 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0844_
timestamp 1644511149
transform -1 0 27508 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0845_
timestamp 1644511149
transform -1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0846_
timestamp 1644511149
transform 1 0 25852 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0847_
timestamp 1644511149
transform -1 0 26588 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0848_
timestamp 1644511149
transform 1 0 26036 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 1644511149
transform -1 0 27232 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0850_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17204 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0851_
timestamp 1644511149
transform 1 0 16100 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0852_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16928 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0853_
timestamp 1644511149
transform -1 0 16100 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0854_
timestamp 1644511149
transform -1 0 17572 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0855_
timestamp 1644511149
transform -1 0 16376 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0856_
timestamp 1644511149
transform -1 0 16192 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0857_
timestamp 1644511149
transform 1 0 13616 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _0858_
timestamp 1644511149
transform 1 0 15916 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0859_
timestamp 1644511149
transform -1 0 14996 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0860_
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0861_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15456 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0862_
timestamp 1644511149
transform -1 0 14996 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0863_
timestamp 1644511149
transform -1 0 13800 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0864_
timestamp 1644511149
transform 1 0 13064 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0865_
timestamp 1644511149
transform -1 0 14812 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0866_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0867_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _0868_
timestamp 1644511149
transform 1 0 12972 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0869_
timestamp 1644511149
transform -1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0870_
timestamp 1644511149
transform 1 0 14812 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1644511149
transform -1 0 15640 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0872_
timestamp 1644511149
transform 1 0 14536 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0873_
timestamp 1644511149
transform 1 0 15824 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1644511149
transform 1 0 14168 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0875_
timestamp 1644511149
transform -1 0 15548 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0876_
timestamp 1644511149
transform 1 0 13340 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0877_
timestamp 1644511149
transform -1 0 15088 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0878_
timestamp 1644511149
transform -1 0 14720 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0879_
timestamp 1644511149
transform 1 0 13156 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0880_
timestamp 1644511149
transform 1 0 12420 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0881_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0882_
timestamp 1644511149
transform -1 0 18124 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0883_
timestamp 1644511149
transform 1 0 12880 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0884_
timestamp 1644511149
transform 1 0 14260 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0885_
timestamp 1644511149
transform 1 0 14076 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0886_
timestamp 1644511149
transform 1 0 13064 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0887_
timestamp 1644511149
transform -1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0888_
timestamp 1644511149
transform 1 0 13340 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0889_
timestamp 1644511149
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0890_
timestamp 1644511149
transform -1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0892_
timestamp 1644511149
transform 1 0 13984 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0893_
timestamp 1644511149
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0894_
timestamp 1644511149
transform 1 0 15824 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 1644511149
transform 1 0 14168 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0896_
timestamp 1644511149
transform -1 0 15916 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0897_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0898_
timestamp 1644511149
transform -1 0 20608 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _0899_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0900_
timestamp 1644511149
transform 1 0 20424 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0901_
timestamp 1644511149
transform -1 0 20240 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0903_
timestamp 1644511149
transform -1 0 16100 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0904_
timestamp 1644511149
transform 1 0 16468 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform -1 0 21068 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0906_
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 1644511149
transform 1 0 14720 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0908_
timestamp 1644511149
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0909_
timestamp 1644511149
transform -1 0 15180 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0910_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0911_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0912_
timestamp 1644511149
transform -1 0 21528 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0913_
timestamp 1644511149
transform 1 0 15824 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0914_
timestamp 1644511149
transform 1 0 17756 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0915_
timestamp 1644511149
transform -1 0 16836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0916_
timestamp 1644511149
transform -1 0 16284 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0917_
timestamp 1644511149
transform 1 0 15272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0918_
timestamp 1644511149
transform 1 0 17572 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0919_
timestamp 1644511149
transform -1 0 18676 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0920_
timestamp 1644511149
transform 1 0 17572 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _0921_
timestamp 1644511149
transform -1 0 17572 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0922_
timestamp 1644511149
transform -1 0 19504 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0923_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0924_
timestamp 1644511149
transform 1 0 19412 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0926_
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _0927_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18952 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0928_
timestamp 1644511149
transform 1 0 18308 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0929_
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0930_
timestamp 1644511149
transform -1 0 20700 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0931_
timestamp 1644511149
transform -1 0 18492 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0932_
timestamp 1644511149
transform 1 0 17940 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0933_
timestamp 1644511149
transform 1 0 19320 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0934_
timestamp 1644511149
transform 1 0 19504 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0935_
timestamp 1644511149
transform -1 0 20148 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0936_
timestamp 1644511149
transform 1 0 20056 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1644511149
transform -1 0 21528 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0939_
timestamp 1644511149
transform -1 0 22356 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0940_
timestamp 1644511149
transform -1 0 22816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0941_
timestamp 1644511149
transform -1 0 22172 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0942_
timestamp 1644511149
transform -1 0 21528 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0943_
timestamp 1644511149
transform 1 0 22448 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0944_
timestamp 1644511149
transform -1 0 20884 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0945_
timestamp 1644511149
transform -1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _0946_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1644511149
transform -1 0 22264 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0948_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 22448 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0949_
timestamp 1644511149
transform -1 0 8096 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 1644511149
transform 1 0 6808 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0951_
timestamp 1644511149
transform 1 0 6440 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0952_
timestamp 1644511149
transform -1 0 7360 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0953_
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0954_
timestamp 1644511149
transform -1 0 5888 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 1644511149
transform -1 0 5244 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0957_
timestamp 1644511149
transform -1 0 5980 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0958_
timestamp 1644511149
transform -1 0 5336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0959_
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0960_
timestamp 1644511149
transform -1 0 5980 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 1644511149
transform 1 0 5428 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0962_
timestamp 1644511149
transform 1 0 6992 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0963_
timestamp 1644511149
transform -1 0 6808 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0965_
timestamp 1644511149
transform 1 0 8280 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0966_
timestamp 1644511149
transform -1 0 7360 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0967_
timestamp 1644511149
transform 1 0 6900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0968_
timestamp 1644511149
transform 1 0 9200 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0969_
timestamp 1644511149
transform 1 0 8832 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0970_
timestamp 1644511149
transform 1 0 9292 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0971_
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0972_
timestamp 1644511149
transform -1 0 9568 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0973_
timestamp 1644511149
transform -1 0 8648 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0974_
timestamp 1644511149
transform 1 0 22356 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0975_
timestamp 1644511149
transform -1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0976_
timestamp 1644511149
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0977_
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0978_
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0979_
timestamp 1644511149
transform 1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0980_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1644511149
transform 1 0 25300 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0982_
timestamp 1644511149
transform -1 0 25668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _0983_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24288 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0984_
timestamp 1644511149
transform 1 0 23736 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform -1 0 26496 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0986_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0987_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25208 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0988_
timestamp 1644511149
transform -1 0 25760 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0989_
timestamp 1644511149
transform -1 0 26312 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0990_
timestamp 1644511149
transform -1 0 26864 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 1644511149
transform 1 0 21344 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0992_
timestamp 1644511149
transform -1 0 24932 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0993_
timestamp 1644511149
transform -1 0 23552 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform -1 0 25392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0995_
timestamp 1644511149
transform -1 0 26220 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0996_
timestamp 1644511149
transform -1 0 26772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0997_
timestamp 1644511149
transform 1 0 24656 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0998_
timestamp 1644511149
transform -1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0999_
timestamp 1644511149
transform 1 0 26128 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1000_
timestamp 1644511149
transform 1 0 26036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1001_
timestamp 1644511149
transform -1 0 27324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1002_
timestamp 1644511149
transform -1 0 24104 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1003_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24472 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1004_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1005_
timestamp 1644511149
transform 1 0 23368 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1006_
timestamp 1644511149
transform 1 0 21804 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1007_
timestamp 1644511149
transform -1 0 24104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1008_
timestamp 1644511149
transform -1 0 24104 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1009_
timestamp 1644511149
transform 1 0 24932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1010_
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1011_
timestamp 1644511149
transform -1 0 22356 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1012_
timestamp 1644511149
transform -1 0 27508 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1013_
timestamp 1644511149
transform -1 0 26588 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1014_
timestamp 1644511149
transform -1 0 26680 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1015_
timestamp 1644511149
transform -1 0 25116 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1016_
timestamp 1644511149
transform -1 0 26496 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1644511149
transform -1 0 27600 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1018_
timestamp 1644511149
transform -1 0 26036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _1019_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1020_
timestamp 1644511149
transform -1 0 26680 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1644511149
transform -1 0 27232 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1022_
timestamp 1644511149
transform 1 0 25944 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1023_
timestamp 1644511149
transform -1 0 25576 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1024_
timestamp 1644511149
transform -1 0 26128 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1025_
timestamp 1644511149
transform 1 0 26036 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1026_
timestamp 1644511149
transform -1 0 22448 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1027_
timestamp 1644511149
transform 1 0 24932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1644511149
transform 1 0 23828 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1644511149
transform -1 0 24932 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1031_
timestamp 1644511149
transform -1 0 23828 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1644511149
transform 1 0 26312 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1033_
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _1034_
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1035_
timestamp 1644511149
transform 1 0 24932 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1036_
timestamp 1644511149
transform 1 0 25392 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1037_
timestamp 1644511149
transform 1 0 25300 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1038_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25392 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1039_
timestamp 1644511149
transform 1 0 14720 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1040_
timestamp 1644511149
transform 1 0 13524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1041_
timestamp 1644511149
transform -1 0 14904 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1042_
timestamp 1644511149
transform 1 0 12236 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1043_
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1044_
timestamp 1644511149
transform 1 0 20792 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1045_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21896 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1644511149
transform 1 0 20608 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1644511149
transform -1 0 27416 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1644511149
transform 1 0 24104 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1644511149
transform 1 0 17480 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1644511149
transform 1 0 15824 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1644511149
transform 1 0 16928 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1644511149
transform -1 0 21528 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1644511149
transform 1 0 17296 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1644511149
transform 1 0 7820 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1644511149
transform 1 0 7820 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1644511149
transform 1 0 7544 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1644511149
transform 1 0 10212 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1644511149
transform -1 0 8648 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1644511149
transform 1 0 8372 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1644511149
transform 1 0 9660 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1644511149
transform 1 0 9660 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1644511149
transform 1 0 12328 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1644511149
transform 1 0 10488 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1644511149
transform 1 0 9936 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1644511149
transform 1 0 9752 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1644511149
transform 1 0 12236 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1644511149
transform 1 0 13800 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1644511149
transform 1 0 9292 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1644511149
transform 1 0 9752 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1644511149
transform 1 0 10120 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1644511149
transform 1 0 11868 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1644511149
transform -1 0 19412 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1644511149
transform -1 0 17480 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1644511149
transform 1 0 14996 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1644511149
transform 1 0 12880 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1644511149
transform -1 0 16560 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1644511149
transform 1 0 11592 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1644511149
transform 1 0 11868 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1644511149
transform 1 0 17480 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1644511149
transform 1 0 17480 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1091_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18308 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1644511149
transform 1 0 16376 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1093_
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1644511149
transform 1 0 17480 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1095_
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1644511149
transform 1 0 26956 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1644511149
transform 1 0 26772 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1644511149
transform -1 0 26128 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1644511149
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1644511149
transform -1 0 23644 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1644511149
transform 1 0 20516 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1644511149
transform 1 0 18952 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1644511149
transform 1 0 18492 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1644511149
transform 1 0 21252 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1644511149
transform -1 0 24932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1644511149
transform 1 0 20424 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1644511149
transform 1 0 18676 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1644511149
transform 1 0 19964 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1644511149
transform -1 0 23276 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1644511149
transform 1 0 24196 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1644511149
transform 1 0 23000 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1644511149
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1644511149
transform 1 0 25208 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1644511149
transform -1 0 13800 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1644511149
transform -1 0 2852 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1644511149
transform -1 0 2852 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1644511149
transform 1 0 13248 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1126_
timestamp 1644511149
transform 1 0 15640 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1127_
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1644511149
transform 1 0 14812 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1644511149
transform 1 0 16100 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1644511149
transform 1 0 18124 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1644511149
transform 1 0 17480 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1644511149
transform -1 0 20608 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1644511149
transform -1 0 23276 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1644511149
transform -1 0 23460 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1644511149
transform -1 0 7728 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1644511149
transform 1 0 5152 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1644511149
transform 1 0 5244 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1644511149
transform 1 0 5152 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1644511149
transform 1 0 5704 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1644511149
transform 1 0 6624 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1644511149
transform 1 0 20056 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1644511149
transform 1 0 22632 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 1644511149
transform 1 0 26956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1644511149
transform 1 0 21896 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1644511149
transform 1 0 26864 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1644511149
transform 1 0 26956 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1644511149
transform 1 0 23460 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1644511149
transform 1 0 22632 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1644511149
transform -1 0 27232 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1644511149
transform 1 0 25208 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1644511149
transform 1 0 14260 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1644511149
transform 1 0 11316 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1644511149
transform -1 0 14628 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1160__33 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1161__34
timestamp 1644511149
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1162__35
timestamp 1644511149
transform -1 0 12604 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1163__36
timestamp 1644511149
transform 1 0 28152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1164__37
timestamp 1644511149
transform -1 0 2300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1165__38
timestamp 1644511149
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1166__39
timestamp 1644511149
transform -1 0 1656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1167__40
timestamp 1644511149
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1168__41
timestamp 1644511149
transform 1 0 28152 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1169__42
timestamp 1644511149
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1170__43
timestamp 1644511149
transform 1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1171__44
timestamp 1644511149
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1172__45
timestamp 1644511149
transform -1 0 1656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1173__46
timestamp 1644511149
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1174__47
timestamp 1644511149
transform -1 0 20608 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1175__48
timestamp 1644511149
transform -1 0 26128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1176__49
timestamp 1644511149
transform -1 0 27416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1177__50
timestamp 1644511149
transform -1 0 19504 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1178__51
timestamp 1644511149
transform 1 0 28152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1179__52
timestamp 1644511149
transform -1 0 6624 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1180__53
timestamp 1644511149
transform -1 0 1656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1181__54
timestamp 1644511149
transform 1 0 28152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1182__55
timestamp 1644511149
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1183__56
timestamp 1644511149
transform -1 0 22080 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clock pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14996 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_clock
timestamp 1644511149
transform -1 0 9568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_clock
timestamp 1644511149
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_clock
timestamp 1644511149
transform -1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_clock
timestamp 1644511149
transform 1 0 11868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_clock
timestamp 1644511149
transform -1 0 20056 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_clock
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_clock
timestamp 1644511149
transform 1 0 19504 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_clock
timestamp 1644511149
transform 1 0 23092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_clock
timestamp 1644511149
transform -1 0 8556 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_clock
timestamp 1644511149
transform -1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_clock
timestamp 1644511149
transform -1 0 13156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_clock
timestamp 1644511149
transform 1 0 13432 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_clock
timestamp 1644511149
transform -1 0 7728 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_clock
timestamp 1644511149
transform -1 0 8648 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_clock
timestamp 1644511149
transform 1 0 13248 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_clock
timestamp 1644511149
transform -1 0 13248 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_clock
timestamp 1644511149
transform -1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_clock
timestamp 1644511149
transform -1 0 19964 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_clock
timestamp 1644511149
transform -1 0 24748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_clock
timestamp 1644511149
transform 1 0 24932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_clock
timestamp 1644511149
transform -1 0 18400 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_clock
timestamp 1644511149
transform 1 0 20424 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_clock
timestamp 1644511149
transform 1 0 24472 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_clock
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform -1 0 28428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1644511149
transform -1 0 28428 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1644511149
transform -1 0 28428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 28152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 28152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1644511149
transform -1 0 28428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input12 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27140 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input13
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1644511149
transform -1 0 28428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform -1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input16
timestamp 1644511149
transform 1 0 25208 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1644511149
transform 1 0 24380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1644511149
transform 1 0 3956 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1644511149
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1644511149
transform 1 0 1564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform -1 0 28428 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1644511149
transform 1 0 28060 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1644511149
transform -1 0 28428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1644511149
transform 1 0 27876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1644511149
transform 1 0 16652 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1644511149
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1644511149
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1644511149
transform 1 0 14904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1644511149
transform -1 0 28428 0 1 26112
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 14968 800 15088 6 clock
port 0 nsew signal input
rlabel metal3 s 29200 24488 30000 24608 6 io_rxd
port 1 nsew signal input
rlabel metal3 s 29200 5448 30000 5568 6 io_txd
port 2 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 io_uartInt
port 3 nsew signal tristate
rlabel metal3 s 29200 23128 30000 23248 6 io_uart_select
port 4 nsew signal input
rlabel metal3 s 29200 17688 30000 17808 6 io_wbs_ack_o
port 5 nsew signal tristate
rlabel metal2 s 13542 29200 13598 30000 6 io_wbs_data_o[0]
port 6 nsew signal tristate
rlabel metal2 s 12254 29200 12310 30000 6 io_wbs_data_o[10]
port 7 nsew signal tristate
rlabel metal3 s 29200 10888 30000 11008 6 io_wbs_data_o[11]
port 8 nsew signal tristate
rlabel metal2 s 1950 29200 2006 30000 6 io_wbs_data_o[12]
port 9 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 io_wbs_data_o[13]
port 10 nsew signal tristate
rlabel metal3 s 0 27208 800 27328 6 io_wbs_data_o[14]
port 11 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 io_wbs_data_o[15]
port 12 nsew signal tristate
rlabel metal3 s 29200 21768 30000 21888 6 io_wbs_data_o[16]
port 13 nsew signal tristate
rlabel metal3 s 0 21768 800 21888 6 io_wbs_data_o[17]
port 14 nsew signal tristate
rlabel metal3 s 29200 19048 30000 19168 6 io_wbs_data_o[18]
port 15 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 io_wbs_data_o[19]
port 16 nsew signal tristate
rlabel metal2 s 27710 29200 27766 30000 6 io_wbs_data_o[1]
port 17 nsew signal tristate
rlabel metal3 s 0 23128 800 23248 6 io_wbs_data_o[20]
port 18 nsew signal tristate
rlabel metal3 s 0 10888 800 11008 6 io_wbs_data_o[21]
port 19 nsew signal tristate
rlabel metal2 s 19982 29200 20038 30000 6 io_wbs_data_o[22]
port 20 nsew signal tristate
rlabel metal2 s 25778 0 25834 800 6 io_wbs_data_o[23]
port 21 nsew signal tristate
rlabel metal2 s 27066 0 27122 800 6 io_wbs_data_o[24]
port 22 nsew signal tristate
rlabel metal2 s 18694 29200 18750 30000 6 io_wbs_data_o[25]
port 23 nsew signal tristate
rlabel metal3 s 29200 20408 30000 20528 6 io_wbs_data_o[26]
port 24 nsew signal tristate
rlabel metal2 s 5814 29200 5870 30000 6 io_wbs_data_o[27]
port 25 nsew signal tristate
rlabel metal3 s 0 17688 800 17808 6 io_wbs_data_o[28]
port 26 nsew signal tristate
rlabel metal3 s 29200 12248 30000 12368 6 io_wbs_data_o[29]
port 27 nsew signal tristate
rlabel metal2 s 16118 29200 16174 30000 6 io_wbs_data_o[2]
port 28 nsew signal tristate
rlabel metal3 s 29200 2728 30000 2848 6 io_wbs_data_o[30]
port 29 nsew signal tristate
rlabel metal2 s 21270 29200 21326 30000 6 io_wbs_data_o[31]
port 30 nsew signal tristate
rlabel metal3 s 0 2728 800 2848 6 io_wbs_data_o[3]
port 31 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 io_wbs_data_o[4]
port 32 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 io_wbs_data_o[5]
port 33 nsew signal tristate
rlabel metal2 s 14830 29200 14886 30000 6 io_wbs_data_o[6]
port 34 nsew signal tristate
rlabel metal3 s 29200 28568 30000 28688 6 io_wbs_data_o[7]
port 35 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 io_wbs_data_o[8]
port 36 nsew signal tristate
rlabel metal3 s 29200 8 30000 128 6 io_wbs_data_o[9]
port 37 nsew signal tristate
rlabel metal3 s 29200 9528 30000 9648 6 io_wbs_m2s_addr[0]
port 38 nsew signal input
rlabel metal2 s 18 29200 74 30000 6 io_wbs_m2s_addr[10]
port 39 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 io_wbs_m2s_addr[11]
port 40 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 io_wbs_m2s_addr[12]
port 41 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 io_wbs_m2s_addr[13]
port 42 nsew signal input
rlabel metal3 s 29200 25848 30000 25968 6 io_wbs_m2s_addr[14]
port 43 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 io_wbs_m2s_addr[15]
port 44 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 io_wbs_m2s_addr[1]
port 45 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 io_wbs_m2s_addr[2]
port 46 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 io_wbs_m2s_addr[3]
port 47 nsew signal input
rlabel metal3 s 29200 8168 30000 8288 6 io_wbs_m2s_addr[4]
port 48 nsew signal input
rlabel metal3 s 29200 4088 30000 4208 6 io_wbs_m2s_addr[5]
port 49 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 io_wbs_m2s_addr[6]
port 50 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 io_wbs_m2s_addr[7]
port 51 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 io_wbs_m2s_addr[8]
port 52 nsew signal input
rlabel metal2 s 8390 29200 8446 30000 6 io_wbs_m2s_addr[9]
port 53 nsew signal input
rlabel metal3 s 29200 6808 30000 6928 6 io_wbs_m2s_data[0]
port 54 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_wbs_m2s_data[10]
port 55 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_wbs_m2s_data[11]
port 56 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 io_wbs_m2s_data[12]
port 57 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_wbs_m2s_data[13]
port 58 nsew signal input
rlabel metal2 s 10966 29200 11022 30000 6 io_wbs_m2s_data[14]
port 59 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_wbs_m2s_data[15]
port 60 nsew signal input
rlabel metal2 s 18 0 74 800 6 io_wbs_m2s_data[16]
port 61 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_wbs_m2s_data[17]
port 62 nsew signal input
rlabel metal2 s 9678 29200 9734 30000 6 io_wbs_m2s_data[18]
port 63 nsew signal input
rlabel metal2 s 17406 29200 17462 30000 6 io_wbs_m2s_data[19]
port 64 nsew signal input
rlabel metal2 s 26422 29200 26478 30000 6 io_wbs_m2s_data[1]
port 65 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_wbs_m2s_data[20]
port 66 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 io_wbs_m2s_data[21]
port 67 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 io_wbs_m2s_data[22]
port 68 nsew signal input
rlabel metal2 s 28998 29200 29054 30000 6 io_wbs_m2s_data[23]
port 69 nsew signal input
rlabel metal2 s 22558 29200 22614 30000 6 io_wbs_m2s_data[24]
port 70 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 io_wbs_m2s_data[25]
port 71 nsew signal input
rlabel metal3 s 29200 27208 30000 27328 6 io_wbs_m2s_data[26]
port 72 nsew signal input
rlabel metal3 s 29200 1368 30000 1488 6 io_wbs_m2s_data[27]
port 73 nsew signal input
rlabel metal2 s 4526 29200 4582 30000 6 io_wbs_m2s_data[28]
port 74 nsew signal input
rlabel metal3 s 29200 14968 30000 15088 6 io_wbs_m2s_data[29]
port 75 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 io_wbs_m2s_data[2]
port 76 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 io_wbs_m2s_data[30]
port 77 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 io_wbs_m2s_data[31]
port 78 nsew signal input
rlabel metal3 s 29200 16328 30000 16448 6 io_wbs_m2s_data[3]
port 79 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 io_wbs_m2s_data[4]
port 80 nsew signal input
rlabel metal2 s 25134 29200 25190 30000 6 io_wbs_m2s_data[5]
port 81 nsew signal input
rlabel metal2 s 23846 29200 23902 30000 6 io_wbs_m2s_data[6]
port 82 nsew signal input
rlabel metal2 s 3238 29200 3294 30000 6 io_wbs_m2s_data[7]
port 83 nsew signal input
rlabel metal2 s 7102 29200 7158 30000 6 io_wbs_m2s_data[8]
port 84 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_wbs_m2s_data[9]
port 85 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 io_wbs_m2s_stb
port 86 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 io_wbs_m2s_we
port 87 nsew signal input
rlabel metal3 s 29200 13608 30000 13728 6 reset
port 88 nsew signal input
rlabel metal4 s 5576 2128 5896 27792 6 vccd1
port 89 nsew power input
rlabel metal4 s 14840 2128 15160 27792 6 vccd1
port 89 nsew power input
rlabel metal4 s 24104 2128 24424 27792 6 vccd1
port 89 nsew power input
rlabel metal4 s 10208 2128 10528 27792 6 vssd1
port 90 nsew ground input
rlabel metal4 s 19472 2128 19792 27792 6 vssd1
port 90 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
