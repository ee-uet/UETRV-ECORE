VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO WB_InterConnect
  CLASS BLOCK ;
  FOREIGN WB_InterConnect ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 1100.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END clock
  PIN io_dbus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END io_dbus_addr[0]
  PIN io_dbus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END io_dbus_addr[10]
  PIN io_dbus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END io_dbus_addr[11]
  PIN io_dbus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END io_dbus_addr[12]
  PIN io_dbus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END io_dbus_addr[13]
  PIN io_dbus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END io_dbus_addr[14]
  PIN io_dbus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END io_dbus_addr[15]
  PIN io_dbus_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END io_dbus_addr[16]
  PIN io_dbus_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END io_dbus_addr[17]
  PIN io_dbus_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END io_dbus_addr[18]
  PIN io_dbus_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END io_dbus_addr[19]
  PIN io_dbus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END io_dbus_addr[1]
  PIN io_dbus_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END io_dbus_addr[20]
  PIN io_dbus_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END io_dbus_addr[21]
  PIN io_dbus_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END io_dbus_addr[22]
  PIN io_dbus_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END io_dbus_addr[23]
  PIN io_dbus_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END io_dbus_addr[24]
  PIN io_dbus_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END io_dbus_addr[25]
  PIN io_dbus_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END io_dbus_addr[26]
  PIN io_dbus_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END io_dbus_addr[27]
  PIN io_dbus_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END io_dbus_addr[28]
  PIN io_dbus_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END io_dbus_addr[29]
  PIN io_dbus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END io_dbus_addr[2]
  PIN io_dbus_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END io_dbus_addr[30]
  PIN io_dbus_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END io_dbus_addr[31]
  PIN io_dbus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END io_dbus_addr[3]
  PIN io_dbus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_dbus_addr[4]
  PIN io_dbus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END io_dbus_addr[5]
  PIN io_dbus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END io_dbus_addr[6]
  PIN io_dbus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END io_dbus_addr[7]
  PIN io_dbus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END io_dbus_addr[8]
  PIN io_dbus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END io_dbus_addr[9]
  PIN io_dbus_ld_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END io_dbus_ld_type[0]
  PIN io_dbus_ld_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END io_dbus_ld_type[1]
  PIN io_dbus_ld_type[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END io_dbus_ld_type[2]
  PIN io_dbus_rd_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END io_dbus_rd_en
  PIN io_dbus_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END io_dbus_rdata[0]
  PIN io_dbus_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END io_dbus_rdata[10]
  PIN io_dbus_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END io_dbus_rdata[11]
  PIN io_dbus_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END io_dbus_rdata[12]
  PIN io_dbus_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END io_dbus_rdata[13]
  PIN io_dbus_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END io_dbus_rdata[14]
  PIN io_dbus_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END io_dbus_rdata[15]
  PIN io_dbus_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END io_dbus_rdata[16]
  PIN io_dbus_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END io_dbus_rdata[17]
  PIN io_dbus_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END io_dbus_rdata[18]
  PIN io_dbus_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END io_dbus_rdata[19]
  PIN io_dbus_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END io_dbus_rdata[1]
  PIN io_dbus_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END io_dbus_rdata[20]
  PIN io_dbus_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END io_dbus_rdata[21]
  PIN io_dbus_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END io_dbus_rdata[22]
  PIN io_dbus_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END io_dbus_rdata[23]
  PIN io_dbus_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END io_dbus_rdata[24]
  PIN io_dbus_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END io_dbus_rdata[25]
  PIN io_dbus_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END io_dbus_rdata[26]
  PIN io_dbus_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 475.360 4.000 475.960 ;
    END
  END io_dbus_rdata[27]
  PIN io_dbus_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END io_dbus_rdata[28]
  PIN io_dbus_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END io_dbus_rdata[29]
  PIN io_dbus_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END io_dbus_rdata[2]
  PIN io_dbus_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.960 4.000 523.560 ;
    END
  END io_dbus_rdata[30]
  PIN io_dbus_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END io_dbus_rdata[31]
  PIN io_dbus_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END io_dbus_rdata[3]
  PIN io_dbus_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END io_dbus_rdata[4]
  PIN io_dbus_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END io_dbus_rdata[5]
  PIN io_dbus_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END io_dbus_rdata[6]
  PIN io_dbus_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_dbus_rdata[7]
  PIN io_dbus_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END io_dbus_rdata[8]
  PIN io_dbus_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END io_dbus_rdata[9]
  PIN io_dbus_st_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END io_dbus_st_type[0]
  PIN io_dbus_st_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END io_dbus_st_type[1]
  PIN io_dbus_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_dbus_valid
  PIN io_dbus_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END io_dbus_wdata[0]
  PIN io_dbus_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END io_dbus_wdata[10]
  PIN io_dbus_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END io_dbus_wdata[11]
  PIN io_dbus_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END io_dbus_wdata[12]
  PIN io_dbus_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END io_dbus_wdata[13]
  PIN io_dbus_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END io_dbus_wdata[14]
  PIN io_dbus_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END io_dbus_wdata[15]
  PIN io_dbus_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END io_dbus_wdata[16]
  PIN io_dbus_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END io_dbus_wdata[17]
  PIN io_dbus_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END io_dbus_wdata[18]
  PIN io_dbus_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END io_dbus_wdata[19]
  PIN io_dbus_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_dbus_wdata[1]
  PIN io_dbus_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END io_dbus_wdata[20]
  PIN io_dbus_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END io_dbus_wdata[21]
  PIN io_dbus_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END io_dbus_wdata[22]
  PIN io_dbus_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END io_dbus_wdata[23]
  PIN io_dbus_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END io_dbus_wdata[24]
  PIN io_dbus_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END io_dbus_wdata[25]
  PIN io_dbus_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END io_dbus_wdata[26]
  PIN io_dbus_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END io_dbus_wdata[27]
  PIN io_dbus_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END io_dbus_wdata[28]
  PIN io_dbus_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.080 4.000 512.680 ;
    END
  END io_dbus_wdata[29]
  PIN io_dbus_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END io_dbus_wdata[2]
  PIN io_dbus_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 528.400 4.000 529.000 ;
    END
  END io_dbus_wdata[30]
  PIN io_dbus_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END io_dbus_wdata[31]
  PIN io_dbus_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_dbus_wdata[3]
  PIN io_dbus_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END io_dbus_wdata[4]
  PIN io_dbus_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END io_dbus_wdata[5]
  PIN io_dbus_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END io_dbus_wdata[6]
  PIN io_dbus_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END io_dbus_wdata[7]
  PIN io_dbus_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END io_dbus_wdata[8]
  PIN io_dbus_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END io_dbus_wdata[9]
  PIN io_dbus_wr_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END io_dbus_wr_en
  PIN io_dmem_io_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 1096.000 21.530 1100.000 ;
    END
  END io_dmem_io_addr[0]
  PIN io_dmem_io_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 1096.000 56.490 1100.000 ;
    END
  END io_dmem_io_addr[1]
  PIN io_dmem_io_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 1096.000 91.450 1100.000 ;
    END
  END io_dmem_io_addr[2]
  PIN io_dmem_io_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 1096.000 126.410 1100.000 ;
    END
  END io_dmem_io_addr[3]
  PIN io_dmem_io_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 1096.000 161.370 1100.000 ;
    END
  END io_dmem_io_addr[4]
  PIN io_dmem_io_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 1096.000 187.590 1100.000 ;
    END
  END io_dmem_io_addr[5]
  PIN io_dmem_io_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 1096.000 213.810 1100.000 ;
    END
  END io_dmem_io_addr[6]
  PIN io_dmem_io_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 1096.000 240.030 1100.000 ;
    END
  END io_dmem_io_addr[7]
  PIN io_dmem_io_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 1096.000 266.250 1100.000 ;
    END
  END io_dmem_io_addr[8]
  PIN io_dmem_io_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 1096.000 4.510 1100.000 ;
    END
  END io_dmem_io_cs
  PIN io_dmem_io_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 1096.000 30.270 1100.000 ;
    END
  END io_dmem_io_rdata[0]
  PIN io_dmem_io_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 1096.000 309.950 1100.000 ;
    END
  END io_dmem_io_rdata[10]
  PIN io_dmem_io_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 1096.000 327.430 1100.000 ;
    END
  END io_dmem_io_rdata[11]
  PIN io_dmem_io_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 1096.000 344.910 1100.000 ;
    END
  END io_dmem_io_rdata[12]
  PIN io_dmem_io_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 1096.000 362.390 1100.000 ;
    END
  END io_dmem_io_rdata[13]
  PIN io_dmem_io_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 1096.000 379.410 1100.000 ;
    END
  END io_dmem_io_rdata[14]
  PIN io_dmem_io_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 1096.000 396.890 1100.000 ;
    END
  END io_dmem_io_rdata[15]
  PIN io_dmem_io_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 1096.000 414.370 1100.000 ;
    END
  END io_dmem_io_rdata[16]
  PIN io_dmem_io_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 1096.000 431.850 1100.000 ;
    END
  END io_dmem_io_rdata[17]
  PIN io_dmem_io_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 1096.000 449.330 1100.000 ;
    END
  END io_dmem_io_rdata[18]
  PIN io_dmem_io_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 1096.000 466.810 1100.000 ;
    END
  END io_dmem_io_rdata[19]
  PIN io_dmem_io_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 1096.000 65.230 1100.000 ;
    END
  END io_dmem_io_rdata[1]
  PIN io_dmem_io_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 1096.000 484.290 1100.000 ;
    END
  END io_dmem_io_rdata[20]
  PIN io_dmem_io_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 1096.000 501.770 1100.000 ;
    END
  END io_dmem_io_rdata[21]
  PIN io_dmem_io_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 1096.000 519.250 1100.000 ;
    END
  END io_dmem_io_rdata[22]
  PIN io_dmem_io_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 1096.000 536.730 1100.000 ;
    END
  END io_dmem_io_rdata[23]
  PIN io_dmem_io_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 1096.000 554.210 1100.000 ;
    END
  END io_dmem_io_rdata[24]
  PIN io_dmem_io_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 1096.000 571.690 1100.000 ;
    END
  END io_dmem_io_rdata[25]
  PIN io_dmem_io_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 1096.000 589.170 1100.000 ;
    END
  END io_dmem_io_rdata[26]
  PIN io_dmem_io_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 1096.000 606.650 1100.000 ;
    END
  END io_dmem_io_rdata[27]
  PIN io_dmem_io_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 1096.000 624.130 1100.000 ;
    END
  END io_dmem_io_rdata[28]
  PIN io_dmem_io_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 1096.000 641.610 1100.000 ;
    END
  END io_dmem_io_rdata[29]
  PIN io_dmem_io_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1096.000 100.190 1100.000 ;
    END
  END io_dmem_io_rdata[2]
  PIN io_dmem_io_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 1096.000 659.090 1100.000 ;
    END
  END io_dmem_io_rdata[30]
  PIN io_dmem_io_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 1096.000 676.570 1100.000 ;
    END
  END io_dmem_io_rdata[31]
  PIN io_dmem_io_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 1096.000 135.150 1100.000 ;
    END
  END io_dmem_io_rdata[3]
  PIN io_dmem_io_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 1096.000 170.110 1100.000 ;
    END
  END io_dmem_io_rdata[4]
  PIN io_dmem_io_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 1096.000 196.330 1100.000 ;
    END
  END io_dmem_io_rdata[5]
  PIN io_dmem_io_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 1096.000 222.550 1100.000 ;
    END
  END io_dmem_io_rdata[6]
  PIN io_dmem_io_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 1096.000 248.770 1100.000 ;
    END
  END io_dmem_io_rdata[7]
  PIN io_dmem_io_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 1096.000 274.990 1100.000 ;
    END
  END io_dmem_io_rdata[8]
  PIN io_dmem_io_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 1096.000 292.470 1100.000 ;
    END
  END io_dmem_io_rdata[9]
  PIN io_dmem_io_st_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1096.000 39.010 1100.000 ;
    END
  END io_dmem_io_st_type[0]
  PIN io_dmem_io_st_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 1096.000 73.970 1100.000 ;
    END
  END io_dmem_io_st_type[1]
  PIN io_dmem_io_st_type[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 1096.000 108.930 1100.000 ;
    END
  END io_dmem_io_st_type[2]
  PIN io_dmem_io_st_type[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 1096.000 143.890 1100.000 ;
    END
  END io_dmem_io_st_type[3]
  PIN io_dmem_io_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 1096.000 47.750 1100.000 ;
    END
  END io_dmem_io_wdata[0]
  PIN io_dmem_io_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 1096.000 318.690 1100.000 ;
    END
  END io_dmem_io_wdata[10]
  PIN io_dmem_io_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 1096.000 336.170 1100.000 ;
    END
  END io_dmem_io_wdata[11]
  PIN io_dmem_io_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 1096.000 353.650 1100.000 ;
    END
  END io_dmem_io_wdata[12]
  PIN io_dmem_io_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 1096.000 371.130 1100.000 ;
    END
  END io_dmem_io_wdata[13]
  PIN io_dmem_io_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 1096.000 388.150 1100.000 ;
    END
  END io_dmem_io_wdata[14]
  PIN io_dmem_io_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 1096.000 405.630 1100.000 ;
    END
  END io_dmem_io_wdata[15]
  PIN io_dmem_io_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 1096.000 423.110 1100.000 ;
    END
  END io_dmem_io_wdata[16]
  PIN io_dmem_io_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 1096.000 440.590 1100.000 ;
    END
  END io_dmem_io_wdata[17]
  PIN io_dmem_io_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 1096.000 458.070 1100.000 ;
    END
  END io_dmem_io_wdata[18]
  PIN io_dmem_io_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 1096.000 475.550 1100.000 ;
    END
  END io_dmem_io_wdata[19]
  PIN io_dmem_io_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 1096.000 82.710 1100.000 ;
    END
  END io_dmem_io_wdata[1]
  PIN io_dmem_io_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 1096.000 493.030 1100.000 ;
    END
  END io_dmem_io_wdata[20]
  PIN io_dmem_io_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 1096.000 510.510 1100.000 ;
    END
  END io_dmem_io_wdata[21]
  PIN io_dmem_io_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 1096.000 527.990 1100.000 ;
    END
  END io_dmem_io_wdata[22]
  PIN io_dmem_io_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 1096.000 545.470 1100.000 ;
    END
  END io_dmem_io_wdata[23]
  PIN io_dmem_io_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 1096.000 562.950 1100.000 ;
    END
  END io_dmem_io_wdata[24]
  PIN io_dmem_io_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 1096.000 580.430 1100.000 ;
    END
  END io_dmem_io_wdata[25]
  PIN io_dmem_io_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 1096.000 597.910 1100.000 ;
    END
  END io_dmem_io_wdata[26]
  PIN io_dmem_io_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 1096.000 615.390 1100.000 ;
    END
  END io_dmem_io_wdata[27]
  PIN io_dmem_io_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 1096.000 632.870 1100.000 ;
    END
  END io_dmem_io_wdata[28]
  PIN io_dmem_io_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 1096.000 650.350 1100.000 ;
    END
  END io_dmem_io_wdata[29]
  PIN io_dmem_io_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 1096.000 117.670 1100.000 ;
    END
  END io_dmem_io_wdata[2]
  PIN io_dmem_io_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 1096.000 667.830 1100.000 ;
    END
  END io_dmem_io_wdata[30]
  PIN io_dmem_io_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 1096.000 685.310 1100.000 ;
    END
  END io_dmem_io_wdata[31]
  PIN io_dmem_io_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 1096.000 152.630 1100.000 ;
    END
  END io_dmem_io_wdata[3]
  PIN io_dmem_io_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 1096.000 178.850 1100.000 ;
    END
  END io_dmem_io_wdata[4]
  PIN io_dmem_io_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 1096.000 205.070 1100.000 ;
    END
  END io_dmem_io_wdata[5]
  PIN io_dmem_io_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 1096.000 231.290 1100.000 ;
    END
  END io_dmem_io_wdata[6]
  PIN io_dmem_io_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 1096.000 257.510 1100.000 ;
    END
  END io_dmem_io_wdata[7]
  PIN io_dmem_io_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1096.000 283.730 1100.000 ;
    END
  END io_dmem_io_wdata[8]
  PIN io_dmem_io_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 1096.000 301.210 1100.000 ;
    END
  END io_dmem_io_wdata[9]
  PIN io_dmem_io_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 1096.000 12.790 1100.000 ;
    END
  END io_dmem_io_wr_en
  PIN io_ibus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END io_ibus_addr[0]
  PIN io_ibus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END io_ibus_addr[10]
  PIN io_ibus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END io_ibus_addr[11]
  PIN io_ibus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END io_ibus_addr[12]
  PIN io_ibus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END io_ibus_addr[13]
  PIN io_ibus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END io_ibus_addr[14]
  PIN io_ibus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END io_ibus_addr[15]
  PIN io_ibus_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END io_ibus_addr[16]
  PIN io_ibus_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.760 4.000 734.360 ;
    END
  END io_ibus_addr[17]
  PIN io_ibus_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END io_ibus_addr[18]
  PIN io_ibus_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END io_ibus_addr[19]
  PIN io_ibus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.120 4.000 565.720 ;
    END
  END io_ibus_addr[1]
  PIN io_ibus_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END io_ibus_addr[20]
  PIN io_ibus_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.920 4.000 776.520 ;
    END
  END io_ibus_addr[21]
  PIN io_ibus_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END io_ibus_addr[22]
  PIN io_ibus_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 796.320 4.000 796.920 ;
    END
  END io_ibus_addr[23]
  PIN io_ibus_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.200 4.000 807.800 ;
    END
  END io_ibus_addr[24]
  PIN io_ibus_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END io_ibus_addr[25]
  PIN io_ibus_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END io_ibus_addr[26]
  PIN io_ibus_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 838.480 4.000 839.080 ;
    END
  END io_ibus_addr[27]
  PIN io_ibus_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 849.360 4.000 849.960 ;
    END
  END io_ibus_addr[28]
  PIN io_ibus_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 4.000 860.160 ;
    END
  END io_ibus_addr[29]
  PIN io_ibus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END io_ibus_addr[2]
  PIN io_ibus_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END io_ibus_addr[30]
  PIN io_ibus_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END io_ibus_addr[31]
  PIN io_ibus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END io_ibus_addr[3]
  PIN io_ibus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 596.400 4.000 597.000 ;
    END
  END io_ibus_addr[4]
  PIN io_ibus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.280 4.000 607.880 ;
    END
  END io_ibus_addr[5]
  PIN io_ibus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END io_ibus_addr[6]
  PIN io_ibus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END io_ibus_addr[7]
  PIN io_ibus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END io_ibus_addr[8]
  PIN io_ibus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END io_ibus_addr[9]
  PIN io_ibus_inst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END io_ibus_inst[0]
  PIN io_ibus_inst[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END io_ibus_inst[10]
  PIN io_ibus_inst[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.280 4.000 675.880 ;
    END
  END io_ibus_inst[11]
  PIN io_ibus_inst[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.160 4.000 686.760 ;
    END
  END io_ibus_inst[12]
  PIN io_ibus_inst[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END io_ibus_inst[13]
  PIN io_ibus_inst[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END io_ibus_inst[14]
  PIN io_ibus_inst[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END io_ibus_inst[15]
  PIN io_ibus_inst[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 728.320 4.000 728.920 ;
    END
  END io_ibus_inst[16]
  PIN io_ibus_inst[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END io_ibus_inst[17]
  PIN io_ibus_inst[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END io_ibus_inst[18]
  PIN io_ibus_inst[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 759.600 4.000 760.200 ;
    END
  END io_ibus_inst[19]
  PIN io_ibus_inst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END io_ibus_inst[1]
  PIN io_ibus_inst[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 770.480 4.000 771.080 ;
    END
  END io_ibus_inst[20]
  PIN io_ibus_inst[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END io_ibus_inst[21]
  PIN io_ibus_inst[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 791.560 4.000 792.160 ;
    END
  END io_ibus_inst[22]
  PIN io_ibus_inst[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.760 4.000 802.360 ;
    END
  END io_ibus_inst[23]
  PIN io_ibus_inst[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END io_ibus_inst[24]
  PIN io_ibus_inst[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END io_ibus_inst[25]
  PIN io_ibus_inst[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.720 4.000 834.320 ;
    END
  END io_ibus_inst[26]
  PIN io_ibus_inst[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.920 4.000 844.520 ;
    END
  END io_ibus_inst[27]
  PIN io_ibus_inst[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.800 4.000 855.400 ;
    END
  END io_ibus_inst[28]
  PIN io_ibus_inst[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END io_ibus_inst[29]
  PIN io_ibus_inst[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END io_ibus_inst[2]
  PIN io_ibus_inst[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END io_ibus_inst[30]
  PIN io_ibus_inst[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.080 4.000 886.680 ;
    END
  END io_ibus_inst[31]
  PIN io_ibus_inst[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END io_ibus_inst[3]
  PIN io_ibus_inst[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END io_ibus_inst[4]
  PIN io_ibus_inst[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 4.000 613.320 ;
    END
  END io_ibus_inst[5]
  PIN io_ibus_inst[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END io_ibus_inst[6]
  PIN io_ibus_inst[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.120 4.000 633.720 ;
    END
  END io_ibus_inst[7]
  PIN io_ibus_inst[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.000 4.000 644.600 ;
    END
  END io_ibus_inst[8]
  PIN io_ibus_inst[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END io_ibus_inst[9]
  PIN io_ibus_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END io_ibus_valid
  PIN io_imem_io_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END io_imem_io_addr[0]
  PIN io_imem_io_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 662.360 1100.000 662.960 ;
    END
  END io_imem_io_addr[1]
  PIN io_imem_io_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 1096.000 746.030 1100.000 ;
    END
  END io_imem_io_addr[2]
  PIN io_imem_io_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 1096.000 754.770 1100.000 ;
    END
  END io_imem_io_addr[3]
  PIN io_imem_io_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END io_imem_io_addr[4]
  PIN io_imem_io_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END io_imem_io_addr[5]
  PIN io_imem_io_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END io_imem_io_addr[6]
  PIN io_imem_io_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END io_imem_io_addr[7]
  PIN io_imem_io_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 775.920 1100.000 776.520 ;
    END
  END io_imem_io_addr[8]
  PIN io_imem_io_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 601.160 1100.000 601.760 ;
    END
  END io_imem_io_cs
  PIN io_imem_io_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 1096.000 702.790 1100.000 ;
    END
  END io_imem_io_rdata[0]
  PIN io_imem_io_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 816.720 1100.000 817.320 ;
    END
  END io_imem_io_rdata[10]
  PIN io_imem_io_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.960 4.000 965.560 ;
    END
  END io_imem_io_rdata[11]
  PIN io_imem_io_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 847.320 1100.000 847.920 ;
    END
  END io_imem_io_rdata[12]
  PIN io_imem_io_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 868.400 1100.000 869.000 ;
    END
  END io_imem_io_rdata[13]
  PIN io_imem_io_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END io_imem_io_rdata[14]
  PIN io_imem_io_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END io_imem_io_rdata[15]
  PIN io_imem_io_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END io_imem_io_rdata[16]
  PIN io_imem_io_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.120 4.000 1007.720 ;
    END
  END io_imem_io_rdata[17]
  PIN io_imem_io_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.000 4.000 1018.600 ;
    END
  END io_imem_io_rdata[18]
  PIN io_imem_io_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.250 1096.000 964.530 1100.000 ;
    END
  END io_imem_io_rdata[19]
  PIN io_imem_io_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 1096.000 729.010 1100.000 ;
    END
  END io_imem_io_rdata[1]
  PIN io_imem_io_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END io_imem_io_rdata[20]
  PIN io_imem_io_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END io_imem_io_rdata[21]
  PIN io_imem_io_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.210 1096.000 999.490 1100.000 ;
    END
  END io_imem_io_rdata[22]
  PIN io_imem_io_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.280 4.000 1049.880 ;
    END
  END io_imem_io_rdata[23]
  PIN io_imem_io_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.160 4.000 1060.760 ;
    END
  END io_imem_io_rdata[24]
  PIN io_imem_io_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 991.480 1100.000 992.080 ;
    END
  END io_imem_io_rdata[25]
  PIN io_imem_io_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.430 1096.000 1025.710 1100.000 ;
    END
  END io_imem_io_rdata[26]
  PIN io_imem_io_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 1096.000 1034.450 1100.000 ;
    END
  END io_imem_io_rdata[27]
  PIN io_imem_io_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END io_imem_io_rdata[28]
  PIN io_imem_io_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 1096.000 1069.410 1100.000 ;
    END
  END io_imem_io_rdata[29]
  PIN io_imem_io_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END io_imem_io_rdata[2]
  PIN io_imem_io_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1063.560 1100.000 1064.160 ;
    END
  END io_imem_io_rdata[30]
  PIN io_imem_io_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1073.760 1100.000 1074.360 ;
    END
  END io_imem_io_rdata[31]
  PIN io_imem_io_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END io_imem_io_rdata[3]
  PIN io_imem_io_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.120 4.000 939.720 ;
    END
  END io_imem_io_rdata[4]
  PIN io_imem_io_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.880 4.000 944.480 ;
    END
  END io_imem_io_rdata[5]
  PIN io_imem_io_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 734.440 1100.000 735.040 ;
    END
  END io_imem_io_rdata[6]
  PIN io_imem_io_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 754.840 1100.000 755.440 ;
    END
  END io_imem_io_rdata[7]
  PIN io_imem_io_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 1096.000 842.170 1100.000 ;
    END
  END io_imem_io_rdata[8]
  PIN io_imem_io_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 954.760 4.000 955.360 ;
    END
  END io_imem_io_rdata[9]
  PIN io_imem_io_st_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 641.960 1100.000 642.560 ;
    END
  END io_imem_io_st_type[0]
  PIN io_imem_io_st_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 1096.000 737.750 1100.000 ;
    END
  END io_imem_io_st_type[1]
  PIN io_imem_io_st_type[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END io_imem_io_st_type[2]
  PIN io_imem_io_st_type[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1096.000 763.510 1100.000 ;
    END
  END io_imem_io_st_type[3]
  PIN io_imem_io_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 1096.000 711.530 1100.000 ;
    END
  END io_imem_io_wdata[0]
  PIN io_imem_io_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 826.920 1100.000 827.520 ;
    END
  END io_imem_io_wdata[10]
  PIN io_imem_io_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END io_imem_io_wdata[11]
  PIN io_imem_io_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.840 4.000 976.440 ;
    END
  END io_imem_io_wdata[12]
  PIN io_imem_io_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 878.600 1100.000 879.200 ;
    END
  END io_imem_io_wdata[13]
  PIN io_imem_io_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 0.000 629.650 4.000 ;
    END
  END io_imem_io_wdata[14]
  PIN io_imem_io_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 0.000 669.670 4.000 ;
    END
  END io_imem_io_wdata[15]
  PIN io_imem_io_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END io_imem_io_wdata[16]
  PIN io_imem_io_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 1096.000 947.050 1100.000 ;
    END
  END io_imem_io_wdata[17]
  PIN io_imem_io_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END io_imem_io_wdata[18]
  PIN io_imem_io_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.990 1096.000 973.270 1100.000 ;
    END
  END io_imem_io_wdata[19]
  PIN io_imem_io_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END io_imem_io_wdata[1]
  PIN io_imem_io_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 0.000 809.510 4.000 ;
    END
  END io_imem_io_wdata[20]
  PIN io_imem_io_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 929.600 1100.000 930.200 ;
    END
  END io_imem_io_wdata[21]
  PIN io_imem_io_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 940.480 1100.000 941.080 ;
    END
  END io_imem_io_wdata[22]
  PIN io_imem_io_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 971.080 1100.000 971.680 ;
    END
  END io_imem_io_wdata[23]
  PIN io_imem_io_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 981.280 1100.000 981.880 ;
    END
  END io_imem_io_wdata[24]
  PIN io_imem_io_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1001.680 1100.000 1002.280 ;
    END
  END io_imem_io_wdata[25]
  PIN io_imem_io_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END io_imem_io_wdata[26]
  PIN io_imem_io_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.530 0.000 949.810 4.000 ;
    END
  END io_imem_io_wdata[27]
  PIN io_imem_io_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 0.000 989.830 4.000 ;
    END
  END io_imem_io_wdata[28]
  PIN io_imem_io_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END io_imem_io_wdata[29]
  PIN io_imem_io_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END io_imem_io_wdata[2]
  PIN io_imem_io_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 1096.000 1095.630 1100.000 ;
    END
  END io_imem_io_wdata[30]
  PIN io_imem_io_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 0.000 1069.870 4.000 ;
    END
  END io_imem_io_wdata[31]
  PIN io_imem_io_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 1096.000 772.250 1100.000 ;
    END
  END io_imem_io_wdata[3]
  PIN io_imem_io_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END io_imem_io_wdata[4]
  PIN io_imem_io_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END io_imem_io_wdata[5]
  PIN io_imem_io_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END io_imem_io_wdata[6]
  PIN io_imem_io_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 1096.000 833.430 1100.000 ;
    END
  END io_imem_io_wdata[7]
  PIN io_imem_io_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 786.120 1100.000 786.720 ;
    END
  END io_imem_io_wdata[8]
  PIN io_imem_io_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 1096.000 850.910 1100.000 ;
    END
  END io_imem_io_wdata[9]
  PIN io_imem_io_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 611.360 1100.000 611.960 ;
    END
  END io_imem_io_wr_en
  PIN io_m1_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 621.560 1100.000 622.160 ;
    END
  END io_m1_ack_i
  PIN io_m1_addr_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END io_m1_addr_sel
  PIN io_m1_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.800 4.000 923.400 ;
    END
  END io_m1_data_i[0]
  PIN io_m1_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END io_m1_data_i[10]
  PIN io_m1_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 970.400 4.000 971.000 ;
    END
  END io_m1_data_i[11]
  PIN io_m1_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 1096.000 885.870 1100.000 ;
    END
  END io_m1_data_i[12]
  PIN io_m1_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END io_m1_data_i[13]
  PIN io_m1_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 1096.000 912.090 1100.000 ;
    END
  END io_m1_data_i[14]
  PIN io_m1_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 991.480 4.000 992.080 ;
    END
  END io_m1_data_i[15]
  PIN io_m1_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 1096.000 938.310 1100.000 ;
    END
  END io_m1_data_i[16]
  PIN io_m1_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1012.560 4.000 1013.160 ;
    END
  END io_m1_data_i[17]
  PIN io_m1_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 0.000 769.490 4.000 ;
    END
  END io_m1_data_i[18]
  PIN io_m1_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.730 1096.000 982.010 1100.000 ;
    END
  END io_m1_data_i[19]
  PIN io_m1_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END io_m1_data_i[1]
  PIN io_m1_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1039.080 4.000 1039.680 ;
    END
  END io_m1_data_i[20]
  PIN io_m1_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.250 0.000 849.530 4.000 ;
    END
  END io_m1_data_i[21]
  PIN io_m1_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 950.680 1100.000 951.280 ;
    END
  END io_m1_data_i[22]
  PIN io_m1_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END io_m1_data_i[23]
  PIN io_m1_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 0.000 889.550 4.000 ;
    END
  END io_m1_data_i[24]
  PIN io_m1_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1070.360 4.000 1070.960 ;
    END
  END io_m1_data_i[25]
  PIN io_m1_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1086.000 4.000 1086.600 ;
    END
  END io_m1_data_i[26]
  PIN io_m1_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.910 1096.000 1043.190 1100.000 ;
    END
  END io_m1_data_i[27]
  PIN io_m1_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.390 1096.000 1060.670 1100.000 ;
    END
  END io_m1_data_i[28]
  PIN io_m1_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.870 1096.000 1078.150 1100.000 ;
    END
  END io_m1_data_i[29]
  PIN io_m1_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 683.440 1100.000 684.040 ;
    END
  END io_m1_data_i[2]
  PIN io_m1_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.880 4.000 1097.480 ;
    END
  END io_m1_data_i[30]
  PIN io_m1_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1083.960 1100.000 1084.560 ;
    END
  END io_m1_data_i[31]
  PIN io_m1_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 1096.000 780.990 1100.000 ;
    END
  END io_m1_data_i[3]
  PIN io_m1_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 714.040 1100.000 714.640 ;
    END
  END io_m1_data_i[4]
  PIN io_m1_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.930 1096.000 807.210 1100.000 ;
    END
  END io_m1_data_i[5]
  PIN io_m1_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1096.000 824.690 1100.000 ;
    END
  END io_m1_data_i[6]
  PIN io_m1_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 765.040 1100.000 765.640 ;
    END
  END io_m1_data_i[7]
  PIN io_m1_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 949.320 4.000 949.920 ;
    END
  END io_m1_data_i[8]
  PIN io_m1_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 959.520 4.000 960.120 ;
    END
  END io_m1_data_i[9]
  PIN io_m2_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_m2_ack_i
  PIN io_m2_addr_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END io_m2_addr_sel
  PIN io_m2_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 1096.000 720.270 1100.000 ;
    END
  END io_m2_data_i[0]
  PIN io_m2_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END io_m2_data_i[10]
  PIN io_m2_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 1096.000 868.390 1100.000 ;
    END
  END io_m2_data_i[11]
  PIN io_m2_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 1096.000 894.610 1100.000 ;
    END
  END io_m2_data_i[12]
  PIN io_m2_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.070 1096.000 903.350 1100.000 ;
    END
  END io_m2_data_i[13]
  PIN io_m2_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END io_m2_data_i[14]
  PIN io_m2_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.920 4.000 997.520 ;
    END
  END io_m2_data_i[15]
  PIN io_m2_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END io_m2_data_i[16]
  PIN io_m2_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 888.800 1100.000 889.400 ;
    END
  END io_m2_data_i[17]
  PIN io_m2_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.510 1096.000 955.790 1100.000 ;
    END
  END io_m2_data_i[18]
  PIN io_m2_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1022.760 4.000 1023.360 ;
    END
  END io_m2_data_i[19]
  PIN io_m2_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 672.560 1100.000 673.160 ;
    END
  END io_m2_data_i[1]
  PIN io_m2_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 909.200 1100.000 909.800 ;
    END
  END io_m2_data_i[20]
  PIN io_m2_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END io_m2_data_i[21]
  PIN io_m2_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 1096.000 1008.230 1100.000 ;
    END
  END io_m2_data_i[22]
  PIN io_m2_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.720 4.000 1055.320 ;
    END
  END io_m2_data_i[23]
  PIN io_m2_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END io_m2_data_i[24]
  PIN io_m2_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.800 4.000 1076.400 ;
    END
  END io_m2_data_i[25]
  PIN io_m2_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1011.880 1100.000 1012.480 ;
    END
  END io_m2_data_i[26]
  PIN io_m2_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1032.960 1100.000 1033.560 ;
    END
  END io_m2_data_i[27]
  PIN io_m2_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1043.160 1100.000 1043.760 ;
    END
  END io_m2_data_i[28]
  PIN io_m2_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 0.000 1009.610 4.000 ;
    END
  END io_m2_data_i[29]
  PIN io_m2_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 693.640 1100.000 694.240 ;
    END
  END io_m2_data_i[2]
  PIN io_m2_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.570 0.000 1029.850 4.000 ;
    END
  END io_m2_data_i[30]
  PIN io_m2_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 0.000 1089.650 4.000 ;
    END
  END io_m2_data_i[31]
  PIN io_m2_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 1096.000 789.730 1100.000 ;
    END
  END io_m2_data_i[3]
  PIN io_m2_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 724.240 1100.000 724.840 ;
    END
  END io_m2_data_i[4]
  PIN io_m2_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END io_m2_data_i[5]
  PIN io_m2_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 744.640 1100.000 745.240 ;
    END
  END io_m2_data_i[6]
  PIN io_m2_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END io_m2_data_i[7]
  PIN io_m2_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 796.320 1100.000 796.920 ;
    END
  END io_m2_data_i[8]
  PIN io_m2_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 806.520 1100.000 807.120 ;
    END
  END io_m2_data_i[9]
  PIN io_m3_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.720 4.000 902.320 ;
    END
  END io_m3_ack_i
  PIN io_m3_addr_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.160 4.000 907.760 ;
    END
  END io_m3_addr_sel
  PIN io_m3_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 652.160 1100.000 652.760 ;
    END
  END io_m3_data_i[0]
  PIN io_m3_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 837.120 1100.000 837.720 ;
    END
  END io_m3_data_i[10]
  PIN io_m3_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850 1096.000 877.130 1100.000 ;
    END
  END io_m3_data_i[11]
  PIN io_m3_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 858.200 1100.000 858.800 ;
    END
  END io_m3_data_i[12]
  PIN io_m3_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END io_m3_data_i[13]
  PIN io_m3_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 1096.000 920.830 1100.000 ;
    END
  END io_m3_data_i[14]
  PIN io_m3_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 1096.000 929.570 1100.000 ;
    END
  END io_m3_data_i[15]
  PIN io_m3_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.680 4.000 1002.280 ;
    END
  END io_m3_data_i[16]
  PIN io_m3_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 899.000 1100.000 899.600 ;
    END
  END io_m3_data_i[17]
  PIN io_m3_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END io_m3_data_i[18]
  PIN io_m3_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1028.200 4.000 1028.800 ;
    END
  END io_m3_data_i[19]
  PIN io_m3_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.680 4.000 934.280 ;
    END
  END io_m3_data_i[1]
  PIN io_m3_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 919.400 1100.000 920.000 ;
    END
  END io_m3_data_i[20]
  PIN io_m3_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 1096.000 990.750 1100.000 ;
    END
  END io_m3_data_i[21]
  PIN io_m3_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 960.880 1100.000 961.480 ;
    END
  END io_m3_data_i[22]
  PIN io_m3_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 1096.000 1016.970 1100.000 ;
    END
  END io_m3_data_i[23]
  PIN io_m3_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.920 4.000 1065.520 ;
    END
  END io_m3_data_i[24]
  PIN io_m3_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END io_m3_data_i[25]
  PIN io_m3_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1022.760 1100.000 1023.360 ;
    END
  END io_m3_data_i[26]
  PIN io_m3_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 1096.000 1051.930 1100.000 ;
    END
  END io_m3_data_i[27]
  PIN io_m3_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1053.360 1100.000 1053.960 ;
    END
  END io_m3_data_i[28]
  PIN io_m3_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.610 1096.000 1086.890 1100.000 ;
    END
  END io_m3_data_i[29]
  PIN io_m3_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 703.840 1100.000 704.440 ;
    END
  END io_m3_data_i[2]
  PIN io_m3_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.350 0.000 1049.630 4.000 ;
    END
  END io_m3_data_i[30]
  PIN io_m3_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1094.160 1100.000 1094.760 ;
    END
  END io_m3_data_i[31]
  PIN io_m3_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 1096.000 798.470 1100.000 ;
    END
  END io_m3_data_i[3]
  PIN io_m3_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END io_m3_data_i[4]
  PIN io_m3_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 1096.000 815.950 1100.000 ;
    END
  END io_m3_data_i[5]
  PIN io_m3_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END io_m3_data_i[6]
  PIN io_m3_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END io_m3_data_i[7]
  PIN io_m3_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END io_m3_data_i[8]
  PIN io_m3_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 1096.000 859.650 1100.000 ;
    END
  END io_m3_data_i[9]
  PIN io_spi_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 559.680 1100.000 560.280 ;
    END
  END io_spi_clk
  PIN io_spi_clk_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 1096.000 694.050 1100.000 ;
    END
  END io_spi_clk_en
  PIN io_spi_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 569.880 1100.000 570.480 ;
    END
  END io_spi_cs
  PIN io_spi_cs_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 912.600 4.000 913.200 ;
    END
  END io_spi_cs_en
  PIN io_spi_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 891.520 4.000 892.120 ;
    END
  END io_spi_irq
  PIN io_spi_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END io_spi_miso
  PIN io_spi_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 580.080 1100.000 580.680 ;
    END
  END io_spi_mosi
  PIN io_spi_mosi_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 631.760 1100.000 632.360 ;
    END
  END io_spi_mosi_en
  PIN io_uart_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.960 4.000 897.560 ;
    END
  END io_uart_irq
  PIN io_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END io_uart_rx
  PIN io_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 590.280 1100.000 590.880 ;
    END
  END io_uart_tx
  PIN io_uart_tx_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END io_uart_tx_en
  PIN io_wbm_m2s_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 25.200 1100.000 25.800 ;
    END
  END io_wbm_m2s_addr[0]
  PIN io_wbm_m2s_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 272.040 1100.000 272.640 ;
    END
  END io_wbm_m2s_addr[10]
  PIN io_wbm_m2s_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 292.440 1100.000 293.040 ;
    END
  END io_wbm_m2s_addr[11]
  PIN io_wbm_m2s_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 312.840 1100.000 313.440 ;
    END
  END io_wbm_m2s_addr[12]
  PIN io_wbm_m2s_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 333.240 1100.000 333.840 ;
    END
  END io_wbm_m2s_addr[13]
  PIN io_wbm_m2s_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 354.320 1100.000 354.920 ;
    END
  END io_wbm_m2s_addr[14]
  PIN io_wbm_m2s_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 374.720 1100.000 375.320 ;
    END
  END io_wbm_m2s_addr[15]
  PIN io_wbm_m2s_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 55.800 1100.000 56.400 ;
    END
  END io_wbm_m2s_addr[1]
  PIN io_wbm_m2s_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 86.400 1100.000 87.000 ;
    END
  END io_wbm_m2s_addr[2]
  PIN io_wbm_m2s_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 117.680 1100.000 118.280 ;
    END
  END io_wbm_m2s_addr[3]
  PIN io_wbm_m2s_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 148.280 1100.000 148.880 ;
    END
  END io_wbm_m2s_addr[4]
  PIN io_wbm_m2s_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 168.680 1100.000 169.280 ;
    END
  END io_wbm_m2s_addr[5]
  PIN io_wbm_m2s_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 189.760 1100.000 190.360 ;
    END
  END io_wbm_m2s_addr[6]
  PIN io_wbm_m2s_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 210.160 1100.000 210.760 ;
    END
  END io_wbm_m2s_addr[7]
  PIN io_wbm_m2s_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 230.560 1100.000 231.160 ;
    END
  END io_wbm_m2s_addr[8]
  PIN io_wbm_m2s_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 250.960 1100.000 251.560 ;
    END
  END io_wbm_m2s_addr[9]
  PIN io_wbm_m2s_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 35.400 1100.000 36.000 ;
    END
  END io_wbm_m2s_data[0]
  PIN io_wbm_m2s_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 282.240 1100.000 282.840 ;
    END
  END io_wbm_m2s_data[10]
  PIN io_wbm_m2s_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 302.640 1100.000 303.240 ;
    END
  END io_wbm_m2s_data[11]
  PIN io_wbm_m2s_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 323.040 1100.000 323.640 ;
    END
  END io_wbm_m2s_data[12]
  PIN io_wbm_m2s_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 344.120 1100.000 344.720 ;
    END
  END io_wbm_m2s_data[13]
  PIN io_wbm_m2s_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 364.520 1100.000 365.120 ;
    END
  END io_wbm_m2s_data[14]
  PIN io_wbm_m2s_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 384.920 1100.000 385.520 ;
    END
  END io_wbm_m2s_data[15]
  PIN io_wbm_m2s_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 395.120 1100.000 395.720 ;
    END
  END io_wbm_m2s_data[16]
  PIN io_wbm_m2s_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 405.320 1100.000 405.920 ;
    END
  END io_wbm_m2s_data[17]
  PIN io_wbm_m2s_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 415.520 1100.000 416.120 ;
    END
  END io_wbm_m2s_data[18]
  PIN io_wbm_m2s_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 425.720 1100.000 426.320 ;
    END
  END io_wbm_m2s_data[19]
  PIN io_wbm_m2s_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 66.000 1100.000 66.600 ;
    END
  END io_wbm_m2s_data[1]
  PIN io_wbm_m2s_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 436.600 1100.000 437.200 ;
    END
  END io_wbm_m2s_data[20]
  PIN io_wbm_m2s_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 446.800 1100.000 447.400 ;
    END
  END io_wbm_m2s_data[21]
  PIN io_wbm_m2s_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 457.000 1100.000 457.600 ;
    END
  END io_wbm_m2s_data[22]
  PIN io_wbm_m2s_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 467.200 1100.000 467.800 ;
    END
  END io_wbm_m2s_data[23]
  PIN io_wbm_m2s_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 477.400 1100.000 478.000 ;
    END
  END io_wbm_m2s_data[24]
  PIN io_wbm_m2s_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 487.600 1100.000 488.200 ;
    END
  END io_wbm_m2s_data[25]
  PIN io_wbm_m2s_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 497.800 1100.000 498.400 ;
    END
  END io_wbm_m2s_data[26]
  PIN io_wbm_m2s_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 508.000 1100.000 508.600 ;
    END
  END io_wbm_m2s_data[27]
  PIN io_wbm_m2s_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 518.880 1100.000 519.480 ;
    END
  END io_wbm_m2s_data[28]
  PIN io_wbm_m2s_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 529.080 1100.000 529.680 ;
    END
  END io_wbm_m2s_data[29]
  PIN io_wbm_m2s_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 97.280 1100.000 97.880 ;
    END
  END io_wbm_m2s_data[2]
  PIN io_wbm_m2s_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 539.280 1100.000 539.880 ;
    END
  END io_wbm_m2s_data[30]
  PIN io_wbm_m2s_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 549.480 1100.000 550.080 ;
    END
  END io_wbm_m2s_data[31]
  PIN io_wbm_m2s_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 127.880 1100.000 128.480 ;
    END
  END io_wbm_m2s_data[3]
  PIN io_wbm_m2s_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 158.480 1100.000 159.080 ;
    END
  END io_wbm_m2s_data[4]
  PIN io_wbm_m2s_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 179.560 1100.000 180.160 ;
    END
  END io_wbm_m2s_data[5]
  PIN io_wbm_m2s_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 199.960 1100.000 200.560 ;
    END
  END io_wbm_m2s_data[6]
  PIN io_wbm_m2s_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 220.360 1100.000 220.960 ;
    END
  END io_wbm_m2s_data[7]
  PIN io_wbm_m2s_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 240.760 1100.000 241.360 ;
    END
  END io_wbm_m2s_data[8]
  PIN io_wbm_m2s_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 261.840 1100.000 262.440 ;
    END
  END io_wbm_m2s_data[9]
  PIN io_wbm_m2s_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 45.600 1100.000 46.200 ;
    END
  END io_wbm_m2s_sel[0]
  PIN io_wbm_m2s_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 76.200 1100.000 76.800 ;
    END
  END io_wbm_m2s_sel[1]
  PIN io_wbm_m2s_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 107.480 1100.000 108.080 ;
    END
  END io_wbm_m2s_sel[2]
  PIN io_wbm_m2s_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 138.080 1100.000 138.680 ;
    END
  END io_wbm_m2s_sel[3]
  PIN io_wbm_m2s_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 4.800 1100.000 5.400 ;
    END
  END io_wbm_m2s_stb
  PIN io_wbm_m2s_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1096.000 15.000 1100.000 15.600 ;
    END
  END io_wbm_m2s_we
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1088.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1088.240 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1094.340 1088.085 ;
      LAYER met1 ;
        RECT 5.520 9.900 1095.650 1088.240 ;
      LAYER met2 ;
        RECT 4.790 1095.720 12.230 1097.365 ;
        RECT 13.070 1095.720 20.970 1097.365 ;
        RECT 21.810 1095.720 29.710 1097.365 ;
        RECT 30.550 1095.720 38.450 1097.365 ;
        RECT 39.290 1095.720 47.190 1097.365 ;
        RECT 48.030 1095.720 55.930 1097.365 ;
        RECT 56.770 1095.720 64.670 1097.365 ;
        RECT 65.510 1095.720 73.410 1097.365 ;
        RECT 74.250 1095.720 82.150 1097.365 ;
        RECT 82.990 1095.720 90.890 1097.365 ;
        RECT 91.730 1095.720 99.630 1097.365 ;
        RECT 100.470 1095.720 108.370 1097.365 ;
        RECT 109.210 1095.720 117.110 1097.365 ;
        RECT 117.950 1095.720 125.850 1097.365 ;
        RECT 126.690 1095.720 134.590 1097.365 ;
        RECT 135.430 1095.720 143.330 1097.365 ;
        RECT 144.170 1095.720 152.070 1097.365 ;
        RECT 152.910 1095.720 160.810 1097.365 ;
        RECT 161.650 1095.720 169.550 1097.365 ;
        RECT 170.390 1095.720 178.290 1097.365 ;
        RECT 179.130 1095.720 187.030 1097.365 ;
        RECT 187.870 1095.720 195.770 1097.365 ;
        RECT 196.610 1095.720 204.510 1097.365 ;
        RECT 205.350 1095.720 213.250 1097.365 ;
        RECT 214.090 1095.720 221.990 1097.365 ;
        RECT 222.830 1095.720 230.730 1097.365 ;
        RECT 231.570 1095.720 239.470 1097.365 ;
        RECT 240.310 1095.720 248.210 1097.365 ;
        RECT 249.050 1095.720 256.950 1097.365 ;
        RECT 257.790 1095.720 265.690 1097.365 ;
        RECT 266.530 1095.720 274.430 1097.365 ;
        RECT 275.270 1095.720 283.170 1097.365 ;
        RECT 284.010 1095.720 291.910 1097.365 ;
        RECT 292.750 1095.720 300.650 1097.365 ;
        RECT 301.490 1095.720 309.390 1097.365 ;
        RECT 310.230 1095.720 318.130 1097.365 ;
        RECT 318.970 1095.720 326.870 1097.365 ;
        RECT 327.710 1095.720 335.610 1097.365 ;
        RECT 336.450 1095.720 344.350 1097.365 ;
        RECT 345.190 1095.720 353.090 1097.365 ;
        RECT 353.930 1095.720 361.830 1097.365 ;
        RECT 362.670 1095.720 370.570 1097.365 ;
        RECT 371.410 1095.720 378.850 1097.365 ;
        RECT 379.690 1095.720 387.590 1097.365 ;
        RECT 388.430 1095.720 396.330 1097.365 ;
        RECT 397.170 1095.720 405.070 1097.365 ;
        RECT 405.910 1095.720 413.810 1097.365 ;
        RECT 414.650 1095.720 422.550 1097.365 ;
        RECT 423.390 1095.720 431.290 1097.365 ;
        RECT 432.130 1095.720 440.030 1097.365 ;
        RECT 440.870 1095.720 448.770 1097.365 ;
        RECT 449.610 1095.720 457.510 1097.365 ;
        RECT 458.350 1095.720 466.250 1097.365 ;
        RECT 467.090 1095.720 474.990 1097.365 ;
        RECT 475.830 1095.720 483.730 1097.365 ;
        RECT 484.570 1095.720 492.470 1097.365 ;
        RECT 493.310 1095.720 501.210 1097.365 ;
        RECT 502.050 1095.720 509.950 1097.365 ;
        RECT 510.790 1095.720 518.690 1097.365 ;
        RECT 519.530 1095.720 527.430 1097.365 ;
        RECT 528.270 1095.720 536.170 1097.365 ;
        RECT 537.010 1095.720 544.910 1097.365 ;
        RECT 545.750 1095.720 553.650 1097.365 ;
        RECT 554.490 1095.720 562.390 1097.365 ;
        RECT 563.230 1095.720 571.130 1097.365 ;
        RECT 571.970 1095.720 579.870 1097.365 ;
        RECT 580.710 1095.720 588.610 1097.365 ;
        RECT 589.450 1095.720 597.350 1097.365 ;
        RECT 598.190 1095.720 606.090 1097.365 ;
        RECT 606.930 1095.720 614.830 1097.365 ;
        RECT 615.670 1095.720 623.570 1097.365 ;
        RECT 624.410 1095.720 632.310 1097.365 ;
        RECT 633.150 1095.720 641.050 1097.365 ;
        RECT 641.890 1095.720 649.790 1097.365 ;
        RECT 650.630 1095.720 658.530 1097.365 ;
        RECT 659.370 1095.720 667.270 1097.365 ;
        RECT 668.110 1095.720 676.010 1097.365 ;
        RECT 676.850 1095.720 684.750 1097.365 ;
        RECT 685.590 1095.720 693.490 1097.365 ;
        RECT 694.330 1095.720 702.230 1097.365 ;
        RECT 703.070 1095.720 710.970 1097.365 ;
        RECT 711.810 1095.720 719.710 1097.365 ;
        RECT 720.550 1095.720 728.450 1097.365 ;
        RECT 729.290 1095.720 737.190 1097.365 ;
        RECT 738.030 1095.720 745.470 1097.365 ;
        RECT 746.310 1095.720 754.210 1097.365 ;
        RECT 755.050 1095.720 762.950 1097.365 ;
        RECT 763.790 1095.720 771.690 1097.365 ;
        RECT 772.530 1095.720 780.430 1097.365 ;
        RECT 781.270 1095.720 789.170 1097.365 ;
        RECT 790.010 1095.720 797.910 1097.365 ;
        RECT 798.750 1095.720 806.650 1097.365 ;
        RECT 807.490 1095.720 815.390 1097.365 ;
        RECT 816.230 1095.720 824.130 1097.365 ;
        RECT 824.970 1095.720 832.870 1097.365 ;
        RECT 833.710 1095.720 841.610 1097.365 ;
        RECT 842.450 1095.720 850.350 1097.365 ;
        RECT 851.190 1095.720 859.090 1097.365 ;
        RECT 859.930 1095.720 867.830 1097.365 ;
        RECT 868.670 1095.720 876.570 1097.365 ;
        RECT 877.410 1095.720 885.310 1097.365 ;
        RECT 886.150 1095.720 894.050 1097.365 ;
        RECT 894.890 1095.720 902.790 1097.365 ;
        RECT 903.630 1095.720 911.530 1097.365 ;
        RECT 912.370 1095.720 920.270 1097.365 ;
        RECT 921.110 1095.720 929.010 1097.365 ;
        RECT 929.850 1095.720 937.750 1097.365 ;
        RECT 938.590 1095.720 946.490 1097.365 ;
        RECT 947.330 1095.720 955.230 1097.365 ;
        RECT 956.070 1095.720 963.970 1097.365 ;
        RECT 964.810 1095.720 972.710 1097.365 ;
        RECT 973.550 1095.720 981.450 1097.365 ;
        RECT 982.290 1095.720 990.190 1097.365 ;
        RECT 991.030 1095.720 998.930 1097.365 ;
        RECT 999.770 1095.720 1007.670 1097.365 ;
        RECT 1008.510 1095.720 1016.410 1097.365 ;
        RECT 1017.250 1095.720 1025.150 1097.365 ;
        RECT 1025.990 1095.720 1033.890 1097.365 ;
        RECT 1034.730 1095.720 1042.630 1097.365 ;
        RECT 1043.470 1095.720 1051.370 1097.365 ;
        RECT 1052.210 1095.720 1060.110 1097.365 ;
        RECT 1060.950 1095.720 1068.850 1097.365 ;
        RECT 1069.690 1095.720 1077.590 1097.365 ;
        RECT 1078.430 1095.720 1086.330 1097.365 ;
        RECT 1087.170 1095.720 1095.070 1097.365 ;
        RECT 4.510 4.280 1095.620 1095.720 ;
        RECT 4.510 2.195 9.470 4.280 ;
        RECT 10.310 2.195 29.250 4.280 ;
        RECT 30.090 2.195 49.030 4.280 ;
        RECT 49.870 2.195 69.270 4.280 ;
        RECT 70.110 2.195 89.050 4.280 ;
        RECT 89.890 2.195 109.290 4.280 ;
        RECT 110.130 2.195 129.070 4.280 ;
        RECT 129.910 2.195 149.310 4.280 ;
        RECT 150.150 2.195 169.090 4.280 ;
        RECT 169.930 2.195 189.330 4.280 ;
        RECT 190.170 2.195 209.110 4.280 ;
        RECT 209.950 2.195 229.350 4.280 ;
        RECT 230.190 2.195 249.130 4.280 ;
        RECT 249.970 2.195 269.370 4.280 ;
        RECT 270.210 2.195 289.150 4.280 ;
        RECT 289.990 2.195 309.390 4.280 ;
        RECT 310.230 2.195 329.170 4.280 ;
        RECT 330.010 2.195 349.410 4.280 ;
        RECT 350.250 2.195 369.190 4.280 ;
        RECT 370.030 2.195 388.970 4.280 ;
        RECT 389.810 2.195 409.210 4.280 ;
        RECT 410.050 2.195 428.990 4.280 ;
        RECT 429.830 2.195 449.230 4.280 ;
        RECT 450.070 2.195 469.010 4.280 ;
        RECT 469.850 2.195 489.250 4.280 ;
        RECT 490.090 2.195 509.030 4.280 ;
        RECT 509.870 2.195 529.270 4.280 ;
        RECT 530.110 2.195 549.050 4.280 ;
        RECT 549.890 2.195 569.290 4.280 ;
        RECT 570.130 2.195 589.070 4.280 ;
        RECT 589.910 2.195 609.310 4.280 ;
        RECT 610.150 2.195 629.090 4.280 ;
        RECT 629.930 2.195 649.330 4.280 ;
        RECT 650.170 2.195 669.110 4.280 ;
        RECT 669.950 2.195 689.350 4.280 ;
        RECT 690.190 2.195 709.130 4.280 ;
        RECT 709.970 2.195 729.370 4.280 ;
        RECT 730.210 2.195 749.150 4.280 ;
        RECT 749.990 2.195 768.930 4.280 ;
        RECT 769.770 2.195 789.170 4.280 ;
        RECT 790.010 2.195 808.950 4.280 ;
        RECT 809.790 2.195 829.190 4.280 ;
        RECT 830.030 2.195 848.970 4.280 ;
        RECT 849.810 2.195 869.210 4.280 ;
        RECT 870.050 2.195 888.990 4.280 ;
        RECT 889.830 2.195 909.230 4.280 ;
        RECT 910.070 2.195 929.010 4.280 ;
        RECT 929.850 2.195 949.250 4.280 ;
        RECT 950.090 2.195 969.030 4.280 ;
        RECT 969.870 2.195 989.270 4.280 ;
        RECT 990.110 2.195 1009.050 4.280 ;
        RECT 1009.890 2.195 1029.290 4.280 ;
        RECT 1030.130 2.195 1049.070 4.280 ;
        RECT 1049.910 2.195 1069.310 4.280 ;
        RECT 1070.150 2.195 1089.090 4.280 ;
        RECT 1089.930 2.195 1095.620 4.280 ;
      LAYER met3 ;
        RECT 4.400 1096.480 1096.000 1097.345 ;
        RECT 4.000 1095.160 1096.000 1096.480 ;
        RECT 4.000 1093.760 1095.600 1095.160 ;
        RECT 4.000 1092.440 1096.000 1093.760 ;
        RECT 4.400 1091.040 1096.000 1092.440 ;
        RECT 4.000 1087.000 1096.000 1091.040 ;
        RECT 4.400 1085.600 1096.000 1087.000 ;
        RECT 4.000 1084.960 1096.000 1085.600 ;
        RECT 4.000 1083.560 1095.600 1084.960 ;
        RECT 4.000 1082.240 1096.000 1083.560 ;
        RECT 4.400 1080.840 1096.000 1082.240 ;
        RECT 4.000 1076.800 1096.000 1080.840 ;
        RECT 4.400 1075.400 1096.000 1076.800 ;
        RECT 4.000 1074.760 1096.000 1075.400 ;
        RECT 4.000 1073.360 1095.600 1074.760 ;
        RECT 4.000 1071.360 1096.000 1073.360 ;
        RECT 4.400 1069.960 1096.000 1071.360 ;
        RECT 4.000 1065.920 1096.000 1069.960 ;
        RECT 4.400 1064.560 1096.000 1065.920 ;
        RECT 4.400 1064.520 1095.600 1064.560 ;
        RECT 4.000 1063.160 1095.600 1064.520 ;
        RECT 4.000 1061.160 1096.000 1063.160 ;
        RECT 4.400 1059.760 1096.000 1061.160 ;
        RECT 4.000 1055.720 1096.000 1059.760 ;
        RECT 4.400 1054.360 1096.000 1055.720 ;
        RECT 4.400 1054.320 1095.600 1054.360 ;
        RECT 4.000 1052.960 1095.600 1054.320 ;
        RECT 4.000 1050.280 1096.000 1052.960 ;
        RECT 4.400 1048.880 1096.000 1050.280 ;
        RECT 4.000 1044.840 1096.000 1048.880 ;
        RECT 4.400 1044.160 1096.000 1044.840 ;
        RECT 4.400 1043.440 1095.600 1044.160 ;
        RECT 4.000 1042.760 1095.600 1043.440 ;
        RECT 4.000 1040.080 1096.000 1042.760 ;
        RECT 4.400 1038.680 1096.000 1040.080 ;
        RECT 4.000 1034.640 1096.000 1038.680 ;
        RECT 4.400 1033.960 1096.000 1034.640 ;
        RECT 4.400 1033.240 1095.600 1033.960 ;
        RECT 4.000 1032.560 1095.600 1033.240 ;
        RECT 4.000 1029.200 1096.000 1032.560 ;
        RECT 4.400 1027.800 1096.000 1029.200 ;
        RECT 4.000 1023.760 1096.000 1027.800 ;
        RECT 4.400 1022.360 1095.600 1023.760 ;
        RECT 4.000 1019.000 1096.000 1022.360 ;
        RECT 4.400 1017.600 1096.000 1019.000 ;
        RECT 4.000 1013.560 1096.000 1017.600 ;
        RECT 4.400 1012.880 1096.000 1013.560 ;
        RECT 4.400 1012.160 1095.600 1012.880 ;
        RECT 4.000 1011.480 1095.600 1012.160 ;
        RECT 4.000 1008.120 1096.000 1011.480 ;
        RECT 4.400 1006.720 1096.000 1008.120 ;
        RECT 4.000 1002.680 1096.000 1006.720 ;
        RECT 4.400 1001.280 1095.600 1002.680 ;
        RECT 4.000 997.920 1096.000 1001.280 ;
        RECT 4.400 996.520 1096.000 997.920 ;
        RECT 4.000 992.480 1096.000 996.520 ;
        RECT 4.400 991.080 1095.600 992.480 ;
        RECT 4.000 987.040 1096.000 991.080 ;
        RECT 4.400 985.640 1096.000 987.040 ;
        RECT 4.000 982.280 1096.000 985.640 ;
        RECT 4.000 981.600 1095.600 982.280 ;
        RECT 4.400 980.880 1095.600 981.600 ;
        RECT 4.400 980.200 1096.000 980.880 ;
        RECT 4.000 976.840 1096.000 980.200 ;
        RECT 4.400 975.440 1096.000 976.840 ;
        RECT 4.000 972.080 1096.000 975.440 ;
        RECT 4.000 971.400 1095.600 972.080 ;
        RECT 4.400 970.680 1095.600 971.400 ;
        RECT 4.400 970.000 1096.000 970.680 ;
        RECT 4.000 965.960 1096.000 970.000 ;
        RECT 4.400 964.560 1096.000 965.960 ;
        RECT 4.000 961.880 1096.000 964.560 ;
        RECT 4.000 960.520 1095.600 961.880 ;
        RECT 4.400 960.480 1095.600 960.520 ;
        RECT 4.400 959.120 1096.000 960.480 ;
        RECT 4.000 955.760 1096.000 959.120 ;
        RECT 4.400 954.360 1096.000 955.760 ;
        RECT 4.000 951.680 1096.000 954.360 ;
        RECT 4.000 950.320 1095.600 951.680 ;
        RECT 4.400 950.280 1095.600 950.320 ;
        RECT 4.400 948.920 1096.000 950.280 ;
        RECT 4.000 944.880 1096.000 948.920 ;
        RECT 4.400 943.480 1096.000 944.880 ;
        RECT 4.000 941.480 1096.000 943.480 ;
        RECT 4.000 940.120 1095.600 941.480 ;
        RECT 4.400 940.080 1095.600 940.120 ;
        RECT 4.400 938.720 1096.000 940.080 ;
        RECT 4.000 934.680 1096.000 938.720 ;
        RECT 4.400 933.280 1096.000 934.680 ;
        RECT 4.000 930.600 1096.000 933.280 ;
        RECT 4.000 929.240 1095.600 930.600 ;
        RECT 4.400 929.200 1095.600 929.240 ;
        RECT 4.400 927.840 1096.000 929.200 ;
        RECT 4.000 923.800 1096.000 927.840 ;
        RECT 4.400 922.400 1096.000 923.800 ;
        RECT 4.000 920.400 1096.000 922.400 ;
        RECT 4.000 919.040 1095.600 920.400 ;
        RECT 4.400 919.000 1095.600 919.040 ;
        RECT 4.400 917.640 1096.000 919.000 ;
        RECT 4.000 913.600 1096.000 917.640 ;
        RECT 4.400 912.200 1096.000 913.600 ;
        RECT 4.000 910.200 1096.000 912.200 ;
        RECT 4.000 908.800 1095.600 910.200 ;
        RECT 4.000 908.160 1096.000 908.800 ;
        RECT 4.400 906.760 1096.000 908.160 ;
        RECT 4.000 902.720 1096.000 906.760 ;
        RECT 4.400 901.320 1096.000 902.720 ;
        RECT 4.000 900.000 1096.000 901.320 ;
        RECT 4.000 898.600 1095.600 900.000 ;
        RECT 4.000 897.960 1096.000 898.600 ;
        RECT 4.400 896.560 1096.000 897.960 ;
        RECT 4.000 892.520 1096.000 896.560 ;
        RECT 4.400 891.120 1096.000 892.520 ;
        RECT 4.000 889.800 1096.000 891.120 ;
        RECT 4.000 888.400 1095.600 889.800 ;
        RECT 4.000 887.080 1096.000 888.400 ;
        RECT 4.400 885.680 1096.000 887.080 ;
        RECT 4.000 881.640 1096.000 885.680 ;
        RECT 4.400 880.240 1096.000 881.640 ;
        RECT 4.000 879.600 1096.000 880.240 ;
        RECT 4.000 878.200 1095.600 879.600 ;
        RECT 4.000 876.880 1096.000 878.200 ;
        RECT 4.400 875.480 1096.000 876.880 ;
        RECT 4.000 871.440 1096.000 875.480 ;
        RECT 4.400 870.040 1096.000 871.440 ;
        RECT 4.000 869.400 1096.000 870.040 ;
        RECT 4.000 868.000 1095.600 869.400 ;
        RECT 4.000 866.000 1096.000 868.000 ;
        RECT 4.400 864.600 1096.000 866.000 ;
        RECT 4.000 860.560 1096.000 864.600 ;
        RECT 4.400 859.200 1096.000 860.560 ;
        RECT 4.400 859.160 1095.600 859.200 ;
        RECT 4.000 857.800 1095.600 859.160 ;
        RECT 4.000 855.800 1096.000 857.800 ;
        RECT 4.400 854.400 1096.000 855.800 ;
        RECT 4.000 850.360 1096.000 854.400 ;
        RECT 4.400 848.960 1096.000 850.360 ;
        RECT 4.000 848.320 1096.000 848.960 ;
        RECT 4.000 846.920 1095.600 848.320 ;
        RECT 4.000 844.920 1096.000 846.920 ;
        RECT 4.400 843.520 1096.000 844.920 ;
        RECT 4.000 839.480 1096.000 843.520 ;
        RECT 4.400 838.120 1096.000 839.480 ;
        RECT 4.400 838.080 1095.600 838.120 ;
        RECT 4.000 836.720 1095.600 838.080 ;
        RECT 4.000 834.720 1096.000 836.720 ;
        RECT 4.400 833.320 1096.000 834.720 ;
        RECT 4.000 829.280 1096.000 833.320 ;
        RECT 4.400 827.920 1096.000 829.280 ;
        RECT 4.400 827.880 1095.600 827.920 ;
        RECT 4.000 826.520 1095.600 827.880 ;
        RECT 4.000 823.840 1096.000 826.520 ;
        RECT 4.400 822.440 1096.000 823.840 ;
        RECT 4.000 818.400 1096.000 822.440 ;
        RECT 4.400 817.720 1096.000 818.400 ;
        RECT 4.400 817.000 1095.600 817.720 ;
        RECT 4.000 816.320 1095.600 817.000 ;
        RECT 4.000 813.640 1096.000 816.320 ;
        RECT 4.400 812.240 1096.000 813.640 ;
        RECT 4.000 808.200 1096.000 812.240 ;
        RECT 4.400 807.520 1096.000 808.200 ;
        RECT 4.400 806.800 1095.600 807.520 ;
        RECT 4.000 806.120 1095.600 806.800 ;
        RECT 4.000 802.760 1096.000 806.120 ;
        RECT 4.400 801.360 1096.000 802.760 ;
        RECT 4.000 797.320 1096.000 801.360 ;
        RECT 4.400 795.920 1095.600 797.320 ;
        RECT 4.000 792.560 1096.000 795.920 ;
        RECT 4.400 791.160 1096.000 792.560 ;
        RECT 4.000 787.120 1096.000 791.160 ;
        RECT 4.400 785.720 1095.600 787.120 ;
        RECT 4.000 781.680 1096.000 785.720 ;
        RECT 4.400 780.280 1096.000 781.680 ;
        RECT 4.000 776.920 1096.000 780.280 ;
        RECT 4.400 775.520 1095.600 776.920 ;
        RECT 4.000 771.480 1096.000 775.520 ;
        RECT 4.400 770.080 1096.000 771.480 ;
        RECT 4.000 766.040 1096.000 770.080 ;
        RECT 4.400 764.640 1095.600 766.040 ;
        RECT 4.000 760.600 1096.000 764.640 ;
        RECT 4.400 759.200 1096.000 760.600 ;
        RECT 4.000 755.840 1096.000 759.200 ;
        RECT 4.400 754.440 1095.600 755.840 ;
        RECT 4.000 750.400 1096.000 754.440 ;
        RECT 4.400 749.000 1096.000 750.400 ;
        RECT 4.000 745.640 1096.000 749.000 ;
        RECT 4.000 744.960 1095.600 745.640 ;
        RECT 4.400 744.240 1095.600 744.960 ;
        RECT 4.400 743.560 1096.000 744.240 ;
        RECT 4.000 739.520 1096.000 743.560 ;
        RECT 4.400 738.120 1096.000 739.520 ;
        RECT 4.000 735.440 1096.000 738.120 ;
        RECT 4.000 734.760 1095.600 735.440 ;
        RECT 4.400 734.040 1095.600 734.760 ;
        RECT 4.400 733.360 1096.000 734.040 ;
        RECT 4.000 729.320 1096.000 733.360 ;
        RECT 4.400 727.920 1096.000 729.320 ;
        RECT 4.000 725.240 1096.000 727.920 ;
        RECT 4.000 723.880 1095.600 725.240 ;
        RECT 4.400 723.840 1095.600 723.880 ;
        RECT 4.400 722.480 1096.000 723.840 ;
        RECT 4.000 718.440 1096.000 722.480 ;
        RECT 4.400 717.040 1096.000 718.440 ;
        RECT 4.000 715.040 1096.000 717.040 ;
        RECT 4.000 713.680 1095.600 715.040 ;
        RECT 4.400 713.640 1095.600 713.680 ;
        RECT 4.400 712.280 1096.000 713.640 ;
        RECT 4.000 708.240 1096.000 712.280 ;
        RECT 4.400 706.840 1096.000 708.240 ;
        RECT 4.000 704.840 1096.000 706.840 ;
        RECT 4.000 703.440 1095.600 704.840 ;
        RECT 4.000 702.800 1096.000 703.440 ;
        RECT 4.400 701.400 1096.000 702.800 ;
        RECT 4.000 697.360 1096.000 701.400 ;
        RECT 4.400 695.960 1096.000 697.360 ;
        RECT 4.000 694.640 1096.000 695.960 ;
        RECT 4.000 693.240 1095.600 694.640 ;
        RECT 4.000 692.600 1096.000 693.240 ;
        RECT 4.400 691.200 1096.000 692.600 ;
        RECT 4.000 687.160 1096.000 691.200 ;
        RECT 4.400 685.760 1096.000 687.160 ;
        RECT 4.000 684.440 1096.000 685.760 ;
        RECT 4.000 683.040 1095.600 684.440 ;
        RECT 4.000 681.720 1096.000 683.040 ;
        RECT 4.400 680.320 1096.000 681.720 ;
        RECT 4.000 676.280 1096.000 680.320 ;
        RECT 4.400 674.880 1096.000 676.280 ;
        RECT 4.000 673.560 1096.000 674.880 ;
        RECT 4.000 672.160 1095.600 673.560 ;
        RECT 4.000 671.520 1096.000 672.160 ;
        RECT 4.400 670.120 1096.000 671.520 ;
        RECT 4.000 666.080 1096.000 670.120 ;
        RECT 4.400 664.680 1096.000 666.080 ;
        RECT 4.000 663.360 1096.000 664.680 ;
        RECT 4.000 661.960 1095.600 663.360 ;
        RECT 4.000 660.640 1096.000 661.960 ;
        RECT 4.400 659.240 1096.000 660.640 ;
        RECT 4.000 655.200 1096.000 659.240 ;
        RECT 4.400 653.800 1096.000 655.200 ;
        RECT 4.000 653.160 1096.000 653.800 ;
        RECT 4.000 651.760 1095.600 653.160 ;
        RECT 4.000 650.440 1096.000 651.760 ;
        RECT 4.400 649.040 1096.000 650.440 ;
        RECT 4.000 645.000 1096.000 649.040 ;
        RECT 4.400 643.600 1096.000 645.000 ;
        RECT 4.000 642.960 1096.000 643.600 ;
        RECT 4.000 641.560 1095.600 642.960 ;
        RECT 4.000 639.560 1096.000 641.560 ;
        RECT 4.400 638.160 1096.000 639.560 ;
        RECT 4.000 634.120 1096.000 638.160 ;
        RECT 4.400 632.760 1096.000 634.120 ;
        RECT 4.400 632.720 1095.600 632.760 ;
        RECT 4.000 631.360 1095.600 632.720 ;
        RECT 4.000 629.360 1096.000 631.360 ;
        RECT 4.400 627.960 1096.000 629.360 ;
        RECT 4.000 623.920 1096.000 627.960 ;
        RECT 4.400 622.560 1096.000 623.920 ;
        RECT 4.400 622.520 1095.600 622.560 ;
        RECT 4.000 621.160 1095.600 622.520 ;
        RECT 4.000 618.480 1096.000 621.160 ;
        RECT 4.400 617.080 1096.000 618.480 ;
        RECT 4.000 613.720 1096.000 617.080 ;
        RECT 4.400 612.360 1096.000 613.720 ;
        RECT 4.400 612.320 1095.600 612.360 ;
        RECT 4.000 610.960 1095.600 612.320 ;
        RECT 4.000 608.280 1096.000 610.960 ;
        RECT 4.400 606.880 1096.000 608.280 ;
        RECT 4.000 602.840 1096.000 606.880 ;
        RECT 4.400 602.160 1096.000 602.840 ;
        RECT 4.400 601.440 1095.600 602.160 ;
        RECT 4.000 600.760 1095.600 601.440 ;
        RECT 4.000 597.400 1096.000 600.760 ;
        RECT 4.400 596.000 1096.000 597.400 ;
        RECT 4.000 592.640 1096.000 596.000 ;
        RECT 4.400 591.280 1096.000 592.640 ;
        RECT 4.400 591.240 1095.600 591.280 ;
        RECT 4.000 589.880 1095.600 591.240 ;
        RECT 4.000 587.200 1096.000 589.880 ;
        RECT 4.400 585.800 1096.000 587.200 ;
        RECT 4.000 581.760 1096.000 585.800 ;
        RECT 4.400 581.080 1096.000 581.760 ;
        RECT 4.400 580.360 1095.600 581.080 ;
        RECT 4.000 579.680 1095.600 580.360 ;
        RECT 4.000 576.320 1096.000 579.680 ;
        RECT 4.400 574.920 1096.000 576.320 ;
        RECT 4.000 571.560 1096.000 574.920 ;
        RECT 4.400 570.880 1096.000 571.560 ;
        RECT 4.400 570.160 1095.600 570.880 ;
        RECT 4.000 569.480 1095.600 570.160 ;
        RECT 4.000 566.120 1096.000 569.480 ;
        RECT 4.400 564.720 1096.000 566.120 ;
        RECT 4.000 560.680 1096.000 564.720 ;
        RECT 4.400 559.280 1095.600 560.680 ;
        RECT 4.000 555.240 1096.000 559.280 ;
        RECT 4.400 553.840 1096.000 555.240 ;
        RECT 4.000 550.480 1096.000 553.840 ;
        RECT 4.400 549.080 1095.600 550.480 ;
        RECT 4.000 545.040 1096.000 549.080 ;
        RECT 4.400 543.640 1096.000 545.040 ;
        RECT 4.000 540.280 1096.000 543.640 ;
        RECT 4.000 539.600 1095.600 540.280 ;
        RECT 4.400 538.880 1095.600 539.600 ;
        RECT 4.400 538.200 1096.000 538.880 ;
        RECT 4.000 534.160 1096.000 538.200 ;
        RECT 4.400 532.760 1096.000 534.160 ;
        RECT 4.000 530.080 1096.000 532.760 ;
        RECT 4.000 529.400 1095.600 530.080 ;
        RECT 4.400 528.680 1095.600 529.400 ;
        RECT 4.400 528.000 1096.000 528.680 ;
        RECT 4.000 523.960 1096.000 528.000 ;
        RECT 4.400 522.560 1096.000 523.960 ;
        RECT 4.000 519.880 1096.000 522.560 ;
        RECT 4.000 518.520 1095.600 519.880 ;
        RECT 4.400 518.480 1095.600 518.520 ;
        RECT 4.400 517.120 1096.000 518.480 ;
        RECT 4.000 513.080 1096.000 517.120 ;
        RECT 4.400 511.680 1096.000 513.080 ;
        RECT 4.000 509.000 1096.000 511.680 ;
        RECT 4.000 508.320 1095.600 509.000 ;
        RECT 4.400 507.600 1095.600 508.320 ;
        RECT 4.400 506.920 1096.000 507.600 ;
        RECT 4.000 502.880 1096.000 506.920 ;
        RECT 4.400 501.480 1096.000 502.880 ;
        RECT 4.000 498.800 1096.000 501.480 ;
        RECT 4.000 497.440 1095.600 498.800 ;
        RECT 4.400 497.400 1095.600 497.440 ;
        RECT 4.400 496.040 1096.000 497.400 ;
        RECT 4.000 492.000 1096.000 496.040 ;
        RECT 4.400 490.600 1096.000 492.000 ;
        RECT 4.000 488.600 1096.000 490.600 ;
        RECT 4.000 487.240 1095.600 488.600 ;
        RECT 4.400 487.200 1095.600 487.240 ;
        RECT 4.400 485.840 1096.000 487.200 ;
        RECT 4.000 481.800 1096.000 485.840 ;
        RECT 4.400 480.400 1096.000 481.800 ;
        RECT 4.000 478.400 1096.000 480.400 ;
        RECT 4.000 477.000 1095.600 478.400 ;
        RECT 4.000 476.360 1096.000 477.000 ;
        RECT 4.400 474.960 1096.000 476.360 ;
        RECT 4.000 471.600 1096.000 474.960 ;
        RECT 4.400 470.200 1096.000 471.600 ;
        RECT 4.000 468.200 1096.000 470.200 ;
        RECT 4.000 466.800 1095.600 468.200 ;
        RECT 4.000 466.160 1096.000 466.800 ;
        RECT 4.400 464.760 1096.000 466.160 ;
        RECT 4.000 460.720 1096.000 464.760 ;
        RECT 4.400 459.320 1096.000 460.720 ;
        RECT 4.000 458.000 1096.000 459.320 ;
        RECT 4.000 456.600 1095.600 458.000 ;
        RECT 4.000 455.280 1096.000 456.600 ;
        RECT 4.400 453.880 1096.000 455.280 ;
        RECT 4.000 450.520 1096.000 453.880 ;
        RECT 4.400 449.120 1096.000 450.520 ;
        RECT 4.000 447.800 1096.000 449.120 ;
        RECT 4.000 446.400 1095.600 447.800 ;
        RECT 4.000 445.080 1096.000 446.400 ;
        RECT 4.400 443.680 1096.000 445.080 ;
        RECT 4.000 439.640 1096.000 443.680 ;
        RECT 4.400 438.240 1096.000 439.640 ;
        RECT 4.000 437.600 1096.000 438.240 ;
        RECT 4.000 436.200 1095.600 437.600 ;
        RECT 4.000 434.200 1096.000 436.200 ;
        RECT 4.400 432.800 1096.000 434.200 ;
        RECT 4.000 429.440 1096.000 432.800 ;
        RECT 4.400 428.040 1096.000 429.440 ;
        RECT 4.000 426.720 1096.000 428.040 ;
        RECT 4.000 425.320 1095.600 426.720 ;
        RECT 4.000 424.000 1096.000 425.320 ;
        RECT 4.400 422.600 1096.000 424.000 ;
        RECT 4.000 418.560 1096.000 422.600 ;
        RECT 4.400 417.160 1096.000 418.560 ;
        RECT 4.000 416.520 1096.000 417.160 ;
        RECT 4.000 415.120 1095.600 416.520 ;
        RECT 4.000 413.120 1096.000 415.120 ;
        RECT 4.400 411.720 1096.000 413.120 ;
        RECT 4.000 408.360 1096.000 411.720 ;
        RECT 4.400 406.960 1096.000 408.360 ;
        RECT 4.000 406.320 1096.000 406.960 ;
        RECT 4.000 404.920 1095.600 406.320 ;
        RECT 4.000 402.920 1096.000 404.920 ;
        RECT 4.400 401.520 1096.000 402.920 ;
        RECT 4.000 397.480 1096.000 401.520 ;
        RECT 4.400 396.120 1096.000 397.480 ;
        RECT 4.400 396.080 1095.600 396.120 ;
        RECT 4.000 394.720 1095.600 396.080 ;
        RECT 4.000 392.040 1096.000 394.720 ;
        RECT 4.400 390.640 1096.000 392.040 ;
        RECT 4.000 387.280 1096.000 390.640 ;
        RECT 4.400 385.920 1096.000 387.280 ;
        RECT 4.400 385.880 1095.600 385.920 ;
        RECT 4.000 384.520 1095.600 385.880 ;
        RECT 4.000 381.840 1096.000 384.520 ;
        RECT 4.400 380.440 1096.000 381.840 ;
        RECT 4.000 376.400 1096.000 380.440 ;
        RECT 4.400 375.720 1096.000 376.400 ;
        RECT 4.400 375.000 1095.600 375.720 ;
        RECT 4.000 374.320 1095.600 375.000 ;
        RECT 4.000 370.960 1096.000 374.320 ;
        RECT 4.400 369.560 1096.000 370.960 ;
        RECT 4.000 366.200 1096.000 369.560 ;
        RECT 4.400 365.520 1096.000 366.200 ;
        RECT 4.400 364.800 1095.600 365.520 ;
        RECT 4.000 364.120 1095.600 364.800 ;
        RECT 4.000 360.760 1096.000 364.120 ;
        RECT 4.400 359.360 1096.000 360.760 ;
        RECT 4.000 355.320 1096.000 359.360 ;
        RECT 4.400 353.920 1095.600 355.320 ;
        RECT 4.000 349.880 1096.000 353.920 ;
        RECT 4.400 348.480 1096.000 349.880 ;
        RECT 4.000 345.120 1096.000 348.480 ;
        RECT 4.400 343.720 1095.600 345.120 ;
        RECT 4.000 339.680 1096.000 343.720 ;
        RECT 4.400 338.280 1096.000 339.680 ;
        RECT 4.000 334.240 1096.000 338.280 ;
        RECT 4.400 332.840 1095.600 334.240 ;
        RECT 4.000 328.800 1096.000 332.840 ;
        RECT 4.400 327.400 1096.000 328.800 ;
        RECT 4.000 324.040 1096.000 327.400 ;
        RECT 4.400 322.640 1095.600 324.040 ;
        RECT 4.000 318.600 1096.000 322.640 ;
        RECT 4.400 317.200 1096.000 318.600 ;
        RECT 4.000 313.840 1096.000 317.200 ;
        RECT 4.000 313.160 1095.600 313.840 ;
        RECT 4.400 312.440 1095.600 313.160 ;
        RECT 4.400 311.760 1096.000 312.440 ;
        RECT 4.000 308.400 1096.000 311.760 ;
        RECT 4.400 307.000 1096.000 308.400 ;
        RECT 4.000 303.640 1096.000 307.000 ;
        RECT 4.000 302.960 1095.600 303.640 ;
        RECT 4.400 302.240 1095.600 302.960 ;
        RECT 4.400 301.560 1096.000 302.240 ;
        RECT 4.000 297.520 1096.000 301.560 ;
        RECT 4.400 296.120 1096.000 297.520 ;
        RECT 4.000 293.440 1096.000 296.120 ;
        RECT 4.000 292.080 1095.600 293.440 ;
        RECT 4.400 292.040 1095.600 292.080 ;
        RECT 4.400 290.680 1096.000 292.040 ;
        RECT 4.000 287.320 1096.000 290.680 ;
        RECT 4.400 285.920 1096.000 287.320 ;
        RECT 4.000 283.240 1096.000 285.920 ;
        RECT 4.000 281.880 1095.600 283.240 ;
        RECT 4.400 281.840 1095.600 281.880 ;
        RECT 4.400 280.480 1096.000 281.840 ;
        RECT 4.000 276.440 1096.000 280.480 ;
        RECT 4.400 275.040 1096.000 276.440 ;
        RECT 4.000 273.040 1096.000 275.040 ;
        RECT 4.000 271.640 1095.600 273.040 ;
        RECT 4.000 271.000 1096.000 271.640 ;
        RECT 4.400 269.600 1096.000 271.000 ;
        RECT 4.000 266.240 1096.000 269.600 ;
        RECT 4.400 264.840 1096.000 266.240 ;
        RECT 4.000 262.840 1096.000 264.840 ;
        RECT 4.000 261.440 1095.600 262.840 ;
        RECT 4.000 260.800 1096.000 261.440 ;
        RECT 4.400 259.400 1096.000 260.800 ;
        RECT 4.000 255.360 1096.000 259.400 ;
        RECT 4.400 253.960 1096.000 255.360 ;
        RECT 4.000 251.960 1096.000 253.960 ;
        RECT 4.000 250.560 1095.600 251.960 ;
        RECT 4.000 249.920 1096.000 250.560 ;
        RECT 4.400 248.520 1096.000 249.920 ;
        RECT 4.000 245.160 1096.000 248.520 ;
        RECT 4.400 243.760 1096.000 245.160 ;
        RECT 4.000 241.760 1096.000 243.760 ;
        RECT 4.000 240.360 1095.600 241.760 ;
        RECT 4.000 239.720 1096.000 240.360 ;
        RECT 4.400 238.320 1096.000 239.720 ;
        RECT 4.000 234.280 1096.000 238.320 ;
        RECT 4.400 232.880 1096.000 234.280 ;
        RECT 4.000 231.560 1096.000 232.880 ;
        RECT 4.000 230.160 1095.600 231.560 ;
        RECT 4.000 228.840 1096.000 230.160 ;
        RECT 4.400 227.440 1096.000 228.840 ;
        RECT 4.000 224.080 1096.000 227.440 ;
        RECT 4.400 222.680 1096.000 224.080 ;
        RECT 4.000 221.360 1096.000 222.680 ;
        RECT 4.000 219.960 1095.600 221.360 ;
        RECT 4.000 218.640 1096.000 219.960 ;
        RECT 4.400 217.240 1096.000 218.640 ;
        RECT 4.000 213.200 1096.000 217.240 ;
        RECT 4.400 211.800 1096.000 213.200 ;
        RECT 4.000 211.160 1096.000 211.800 ;
        RECT 4.000 209.760 1095.600 211.160 ;
        RECT 4.000 207.760 1096.000 209.760 ;
        RECT 4.400 206.360 1096.000 207.760 ;
        RECT 4.000 203.000 1096.000 206.360 ;
        RECT 4.400 201.600 1096.000 203.000 ;
        RECT 4.000 200.960 1096.000 201.600 ;
        RECT 4.000 199.560 1095.600 200.960 ;
        RECT 4.000 197.560 1096.000 199.560 ;
        RECT 4.400 196.160 1096.000 197.560 ;
        RECT 4.000 192.120 1096.000 196.160 ;
        RECT 4.400 190.760 1096.000 192.120 ;
        RECT 4.400 190.720 1095.600 190.760 ;
        RECT 4.000 189.360 1095.600 190.720 ;
        RECT 4.000 186.680 1096.000 189.360 ;
        RECT 4.400 185.280 1096.000 186.680 ;
        RECT 4.000 181.920 1096.000 185.280 ;
        RECT 4.400 180.560 1096.000 181.920 ;
        RECT 4.400 180.520 1095.600 180.560 ;
        RECT 4.000 179.160 1095.600 180.520 ;
        RECT 4.000 176.480 1096.000 179.160 ;
        RECT 4.400 175.080 1096.000 176.480 ;
        RECT 4.000 171.040 1096.000 175.080 ;
        RECT 4.400 169.680 1096.000 171.040 ;
        RECT 4.400 169.640 1095.600 169.680 ;
        RECT 4.000 168.280 1095.600 169.640 ;
        RECT 4.000 165.600 1096.000 168.280 ;
        RECT 4.400 164.200 1096.000 165.600 ;
        RECT 4.000 160.840 1096.000 164.200 ;
        RECT 4.400 159.480 1096.000 160.840 ;
        RECT 4.400 159.440 1095.600 159.480 ;
        RECT 4.000 158.080 1095.600 159.440 ;
        RECT 4.000 155.400 1096.000 158.080 ;
        RECT 4.400 154.000 1096.000 155.400 ;
        RECT 4.000 149.960 1096.000 154.000 ;
        RECT 4.400 149.280 1096.000 149.960 ;
        RECT 4.400 148.560 1095.600 149.280 ;
        RECT 4.000 147.880 1095.600 148.560 ;
        RECT 4.000 145.200 1096.000 147.880 ;
        RECT 4.400 143.800 1096.000 145.200 ;
        RECT 4.000 139.760 1096.000 143.800 ;
        RECT 4.400 139.080 1096.000 139.760 ;
        RECT 4.400 138.360 1095.600 139.080 ;
        RECT 4.000 137.680 1095.600 138.360 ;
        RECT 4.000 134.320 1096.000 137.680 ;
        RECT 4.400 132.920 1096.000 134.320 ;
        RECT 4.000 128.880 1096.000 132.920 ;
        RECT 4.400 127.480 1095.600 128.880 ;
        RECT 4.000 124.120 1096.000 127.480 ;
        RECT 4.400 122.720 1096.000 124.120 ;
        RECT 4.000 118.680 1096.000 122.720 ;
        RECT 4.400 117.280 1095.600 118.680 ;
        RECT 4.000 113.240 1096.000 117.280 ;
        RECT 4.400 111.840 1096.000 113.240 ;
        RECT 4.000 108.480 1096.000 111.840 ;
        RECT 4.000 107.800 1095.600 108.480 ;
        RECT 4.400 107.080 1095.600 107.800 ;
        RECT 4.400 106.400 1096.000 107.080 ;
        RECT 4.000 103.040 1096.000 106.400 ;
        RECT 4.400 101.640 1096.000 103.040 ;
        RECT 4.000 98.280 1096.000 101.640 ;
        RECT 4.000 97.600 1095.600 98.280 ;
        RECT 4.400 96.880 1095.600 97.600 ;
        RECT 4.400 96.200 1096.000 96.880 ;
        RECT 4.000 92.160 1096.000 96.200 ;
        RECT 4.400 90.760 1096.000 92.160 ;
        RECT 4.000 87.400 1096.000 90.760 ;
        RECT 4.000 86.720 1095.600 87.400 ;
        RECT 4.400 86.000 1095.600 86.720 ;
        RECT 4.400 85.320 1096.000 86.000 ;
        RECT 4.000 81.960 1096.000 85.320 ;
        RECT 4.400 80.560 1096.000 81.960 ;
        RECT 4.000 77.200 1096.000 80.560 ;
        RECT 4.000 76.520 1095.600 77.200 ;
        RECT 4.400 75.800 1095.600 76.520 ;
        RECT 4.400 75.120 1096.000 75.800 ;
        RECT 4.000 71.080 1096.000 75.120 ;
        RECT 4.400 69.680 1096.000 71.080 ;
        RECT 4.000 67.000 1096.000 69.680 ;
        RECT 4.000 65.640 1095.600 67.000 ;
        RECT 4.400 65.600 1095.600 65.640 ;
        RECT 4.400 64.240 1096.000 65.600 ;
        RECT 4.000 60.880 1096.000 64.240 ;
        RECT 4.400 59.480 1096.000 60.880 ;
        RECT 4.000 56.800 1096.000 59.480 ;
        RECT 4.000 55.440 1095.600 56.800 ;
        RECT 4.400 55.400 1095.600 55.440 ;
        RECT 4.400 54.040 1096.000 55.400 ;
        RECT 4.000 50.000 1096.000 54.040 ;
        RECT 4.400 48.600 1096.000 50.000 ;
        RECT 4.000 46.600 1096.000 48.600 ;
        RECT 4.000 45.200 1095.600 46.600 ;
        RECT 4.000 44.560 1096.000 45.200 ;
        RECT 4.400 43.160 1096.000 44.560 ;
        RECT 4.000 39.800 1096.000 43.160 ;
        RECT 4.400 38.400 1096.000 39.800 ;
        RECT 4.000 36.400 1096.000 38.400 ;
        RECT 4.000 35.000 1095.600 36.400 ;
        RECT 4.000 34.360 1096.000 35.000 ;
        RECT 4.400 32.960 1096.000 34.360 ;
        RECT 4.000 28.920 1096.000 32.960 ;
        RECT 4.400 27.520 1096.000 28.920 ;
        RECT 4.000 26.200 1096.000 27.520 ;
        RECT 4.000 24.800 1095.600 26.200 ;
        RECT 4.000 23.480 1096.000 24.800 ;
        RECT 4.400 22.080 1096.000 23.480 ;
        RECT 4.000 18.720 1096.000 22.080 ;
        RECT 4.400 17.320 1096.000 18.720 ;
        RECT 4.000 16.000 1096.000 17.320 ;
        RECT 4.000 14.600 1095.600 16.000 ;
        RECT 4.000 13.280 1096.000 14.600 ;
        RECT 4.400 11.880 1096.000 13.280 ;
        RECT 4.000 7.840 1096.000 11.880 ;
        RECT 4.400 6.440 1096.000 7.840 ;
        RECT 4.000 5.800 1096.000 6.440 ;
        RECT 4.000 4.400 1095.600 5.800 ;
        RECT 4.000 3.080 1096.000 4.400 ;
        RECT 4.400 2.215 1096.000 3.080 ;
      LAYER met4 ;
        RECT 59.175 134.135 97.440 1085.785 ;
        RECT 99.840 134.135 174.240 1085.785 ;
        RECT 176.640 134.135 251.040 1085.785 ;
        RECT 253.440 134.135 327.840 1085.785 ;
        RECT 330.240 134.135 404.640 1085.785 ;
        RECT 407.040 134.135 481.440 1085.785 ;
        RECT 483.840 134.135 558.240 1085.785 ;
        RECT 560.640 134.135 635.040 1085.785 ;
        RECT 637.440 134.135 711.840 1085.785 ;
        RECT 714.240 134.135 788.640 1085.785 ;
        RECT 791.040 134.135 865.440 1085.785 ;
        RECT 867.840 134.135 942.240 1085.785 ;
        RECT 944.640 134.135 1019.040 1085.785 ;
        RECT 1021.440 134.135 1088.985 1085.785 ;
  END
END WB_InterConnect
END LIBRARY

