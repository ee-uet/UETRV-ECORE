magic
tech sky130A
magscale 1 2
timestamp 1647680207
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2048 98808 97424
<< metal2 >>
rect 1674 99200 1730 100000
rect 4986 99200 5042 100000
rect 8298 99200 8354 100000
rect 11610 99200 11666 100000
rect 14922 99200 14978 100000
rect 18326 99200 18382 100000
rect 21638 99200 21694 100000
rect 24950 99200 25006 100000
rect 28262 99200 28318 100000
rect 31666 99200 31722 100000
rect 34978 99200 35034 100000
rect 38290 99200 38346 100000
rect 41602 99200 41658 100000
rect 45006 99200 45062 100000
rect 48318 99200 48374 100000
rect 51630 99200 51686 100000
rect 54942 99200 54998 100000
rect 58254 99200 58310 100000
rect 61658 99200 61714 100000
rect 64970 99200 65026 100000
rect 68282 99200 68338 100000
rect 71594 99200 71650 100000
rect 74998 99200 75054 100000
rect 78310 99200 78366 100000
rect 81622 99200 81678 100000
rect 84934 99200 84990 100000
rect 88338 99200 88394 100000
rect 91650 99200 91706 100000
rect 94962 99200 95018 100000
rect 98274 99200 98330 100000
rect 2318 0 2374 800
rect 7010 0 7066 800
rect 11794 0 11850 800
rect 16578 0 16634 800
rect 21362 0 21418 800
rect 26054 0 26110 800
rect 30838 0 30894 800
rect 35622 0 35678 800
rect 40406 0 40462 800
rect 45098 0 45154 800
rect 49882 0 49938 800
rect 54666 0 54722 800
rect 59450 0 59506 800
rect 64142 0 64198 800
rect 68926 0 68982 800
rect 73710 0 73766 800
rect 78494 0 78550 800
rect 83186 0 83242 800
rect 87970 0 88026 800
rect 92754 0 92810 800
rect 97538 0 97594 800
<< obsm2 >>
rect 1398 99144 1618 99362
rect 1786 99144 4930 99362
rect 5098 99144 8242 99362
rect 8410 99144 11554 99362
rect 11722 99144 14866 99362
rect 15034 99144 18270 99362
rect 18438 99144 21582 99362
rect 21750 99144 24894 99362
rect 25062 99144 28206 99362
rect 28374 99144 31610 99362
rect 31778 99144 34922 99362
rect 35090 99144 38234 99362
rect 38402 99144 41546 99362
rect 41714 99144 44950 99362
rect 45118 99144 48262 99362
rect 48430 99144 51574 99362
rect 51742 99144 54886 99362
rect 55054 99144 58198 99362
rect 58366 99144 61602 99362
rect 61770 99144 64914 99362
rect 65082 99144 68226 99362
rect 68394 99144 71538 99362
rect 71706 99144 74942 99362
rect 75110 99144 78254 99362
rect 78422 99144 81566 99362
rect 81734 99144 84878 99362
rect 85046 99144 88282 99362
rect 88450 99144 91594 99362
rect 91762 99144 94906 99362
rect 95074 99144 98218 99362
rect 1398 856 98330 99144
rect 1398 734 2262 856
rect 2430 734 6954 856
rect 7122 734 11738 856
rect 11906 734 16522 856
rect 16690 734 21306 856
rect 21474 734 25998 856
rect 26166 734 30782 856
rect 30950 734 35566 856
rect 35734 734 40350 856
rect 40518 734 45042 856
rect 45210 734 49826 856
rect 49994 734 54610 856
rect 54778 734 59394 856
rect 59562 734 64086 856
rect 64254 734 68870 856
rect 69038 734 73654 856
rect 73822 734 78438 856
rect 78606 734 83130 856
rect 83298 734 87914 856
rect 88082 734 92698 856
rect 92866 734 97482 856
rect 97650 734 98330 856
<< metal3 >>
rect 99200 98064 100000 98184
rect 0 96568 800 96688
rect 99200 94664 100000 94784
rect 99200 91128 100000 91248
rect 0 89904 800 90024
rect 99200 87728 100000 87848
rect 99200 84328 100000 84448
rect 0 83240 800 83360
rect 99200 80792 100000 80912
rect 99200 77392 100000 77512
rect 0 76576 800 76696
rect 99200 73992 100000 74112
rect 99200 70456 100000 70576
rect 0 69912 800 70032
rect 99200 67056 100000 67176
rect 99200 63656 100000 63776
rect 0 63248 800 63368
rect 99200 60120 100000 60240
rect 0 56584 800 56704
rect 99200 56720 100000 56840
rect 99200 53320 100000 53440
rect 0 49920 800 50040
rect 99200 49784 100000 49904
rect 99200 46384 100000 46504
rect 0 43256 800 43376
rect 99200 42984 100000 43104
rect 99200 39448 100000 39568
rect 0 36592 800 36712
rect 99200 36048 100000 36168
rect 99200 32648 100000 32768
rect 0 29928 800 30048
rect 99200 29112 100000 29232
rect 99200 25712 100000 25832
rect 0 23264 800 23384
rect 99200 22312 100000 22432
rect 99200 18776 100000 18896
rect 0 16600 800 16720
rect 99200 15376 100000 15496
rect 99200 11976 100000 12096
rect 0 9936 800 10056
rect 99200 8440 100000 8560
rect 99200 5040 100000 5160
rect 0 3272 800 3392
rect 99200 1640 100000 1760
<< obsm3 >>
rect 800 97984 99120 98157
rect 800 96768 99200 97984
rect 880 96488 99200 96768
rect 800 94864 99200 96488
rect 800 94584 99120 94864
rect 800 91328 99200 94584
rect 800 91048 99120 91328
rect 800 90104 99200 91048
rect 880 89824 99200 90104
rect 800 87928 99200 89824
rect 800 87648 99120 87928
rect 800 84528 99200 87648
rect 800 84248 99120 84528
rect 800 83440 99200 84248
rect 880 83160 99200 83440
rect 800 80992 99200 83160
rect 800 80712 99120 80992
rect 800 77592 99200 80712
rect 800 77312 99120 77592
rect 800 76776 99200 77312
rect 880 76496 99200 76776
rect 800 74192 99200 76496
rect 800 73912 99120 74192
rect 800 70656 99200 73912
rect 800 70376 99120 70656
rect 800 70112 99200 70376
rect 880 69832 99200 70112
rect 800 67256 99200 69832
rect 800 66976 99120 67256
rect 800 63856 99200 66976
rect 800 63576 99120 63856
rect 800 63448 99200 63576
rect 880 63168 99200 63448
rect 800 60320 99200 63168
rect 800 60040 99120 60320
rect 800 56920 99200 60040
rect 800 56784 99120 56920
rect 880 56640 99120 56784
rect 880 56504 99200 56640
rect 800 53520 99200 56504
rect 800 53240 99120 53520
rect 800 50120 99200 53240
rect 880 49984 99200 50120
rect 880 49840 99120 49984
rect 800 49704 99120 49840
rect 800 46584 99200 49704
rect 800 46304 99120 46584
rect 800 43456 99200 46304
rect 880 43184 99200 43456
rect 880 43176 99120 43184
rect 800 42904 99120 43176
rect 800 39648 99200 42904
rect 800 39368 99120 39648
rect 800 36792 99200 39368
rect 880 36512 99200 36792
rect 800 36248 99200 36512
rect 800 35968 99120 36248
rect 800 32848 99200 35968
rect 800 32568 99120 32848
rect 800 30128 99200 32568
rect 880 29848 99200 30128
rect 800 29312 99200 29848
rect 800 29032 99120 29312
rect 800 25912 99200 29032
rect 800 25632 99120 25912
rect 800 23464 99200 25632
rect 880 23184 99200 23464
rect 800 22512 99200 23184
rect 800 22232 99120 22512
rect 800 18976 99200 22232
rect 800 18696 99120 18976
rect 800 16800 99200 18696
rect 880 16520 99200 16800
rect 800 15576 99200 16520
rect 800 15296 99120 15576
rect 800 12176 99200 15296
rect 800 11896 99120 12176
rect 800 10136 99200 11896
rect 880 9856 99200 10136
rect 800 8640 99200 9856
rect 800 8360 99120 8640
rect 800 5240 99200 8360
rect 800 4960 99120 5240
rect 800 3472 99200 4960
rect 880 3192 99200 3472
rect 800 1840 99200 3192
rect 800 1667 99120 1840
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 46059 2619 50208 97069
rect 50688 2619 65568 97069
rect 66048 2619 80928 97069
rect 81408 2619 90837 97069
<< labels >>
rlabel metal2 s 2318 0 2374 800 6 clock
port 1 nsew signal input
rlabel metal2 s 8298 99200 8354 100000 6 io_ba_match
port 2 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 io_motor_irq
port 3 nsew signal output
rlabel metal2 s 1674 99200 1730 100000 6 io_pwm_high
port 4 nsew signal output
rlabel metal2 s 4986 99200 5042 100000 6 io_pwm_low
port 5 nsew signal output
rlabel metal3 s 99200 1640 100000 1760 6 io_qei_ch_a
port 6 nsew signal input
rlabel metal2 s 11610 99200 11666 100000 6 io_qei_ch_b
port 7 nsew signal input
rlabel metal3 s 99200 5040 100000 5160 6 io_wbs_ack_o
port 8 nsew signal output
rlabel metal3 s 99200 15376 100000 15496 6 io_wbs_data_o[0]
port 9 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 io_wbs_data_o[10]
port 10 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 io_wbs_data_o[11]
port 11 nsew signal output
rlabel metal2 s 54942 99200 54998 100000 6 io_wbs_data_o[12]
port 12 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 io_wbs_data_o[13]
port 13 nsew signal output
rlabel metal2 s 58254 99200 58310 100000 6 io_wbs_data_o[14]
port 14 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 io_wbs_data_o[15]
port 15 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 io_wbs_data_o[16]
port 16 nsew signal output
rlabel metal3 s 99200 67056 100000 67176 6 io_wbs_data_o[17]
port 17 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 io_wbs_data_o[18]
port 18 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 io_wbs_data_o[19]
port 19 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 io_wbs_data_o[1]
port 20 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 io_wbs_data_o[20]
port 21 nsew signal output
rlabel metal2 s 78310 99200 78366 100000 6 io_wbs_data_o[21]
port 22 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 io_wbs_data_o[22]
port 23 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 io_wbs_data_o[23]
port 24 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 io_wbs_data_o[24]
port 25 nsew signal output
rlabel metal2 s 88338 99200 88394 100000 6 io_wbs_data_o[25]
port 26 nsew signal output
rlabel metal3 s 99200 84328 100000 84448 6 io_wbs_data_o[26]
port 27 nsew signal output
rlabel metal2 s 91650 99200 91706 100000 6 io_wbs_data_o[27]
port 28 nsew signal output
rlabel metal2 s 94962 99200 95018 100000 6 io_wbs_data_o[28]
port 29 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 io_wbs_data_o[29]
port 30 nsew signal output
rlabel metal2 s 18326 99200 18382 100000 6 io_wbs_data_o[2]
port 31 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 io_wbs_data_o[30]
port 32 nsew signal output
rlabel metal3 s 99200 94664 100000 94784 6 io_wbs_data_o[31]
port 33 nsew signal output
rlabel metal2 s 21638 99200 21694 100000 6 io_wbs_data_o[3]
port 34 nsew signal output
rlabel metal2 s 28262 99200 28318 100000 6 io_wbs_data_o[4]
port 35 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 io_wbs_data_o[5]
port 36 nsew signal output
rlabel metal3 s 99200 32648 100000 32768 6 io_wbs_data_o[6]
port 37 nsew signal output
rlabel metal2 s 38290 99200 38346 100000 6 io_wbs_data_o[7]
port 38 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 io_wbs_data_o[8]
port 39 nsew signal output
rlabel metal3 s 99200 46384 100000 46504 6 io_wbs_data_o[9]
port 40 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 io_wbs_m2s_addr[0]
port 41 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 io_wbs_m2s_addr[10]
port 42 nsew signal input
rlabel metal3 s 99200 53320 100000 53440 6 io_wbs_m2s_addr[11]
port 43 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 io_wbs_m2s_addr[12]
port 44 nsew signal input
rlabel metal3 s 99200 56720 100000 56840 6 io_wbs_m2s_addr[13]
port 45 nsew signal input
rlabel metal2 s 61658 99200 61714 100000 6 io_wbs_m2s_addr[14]
port 46 nsew signal input
rlabel metal2 s 68282 99200 68338 100000 6 io_wbs_m2s_addr[15]
port 47 nsew signal input
rlabel metal3 s 99200 18776 100000 18896 6 io_wbs_m2s_addr[1]
port 48 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 io_wbs_m2s_addr[2]
port 49 nsew signal input
rlabel metal2 s 24950 99200 25006 100000 6 io_wbs_m2s_addr[3]
port 50 nsew signal input
rlabel metal2 s 31666 99200 31722 100000 6 io_wbs_m2s_addr[4]
port 51 nsew signal input
rlabel metal3 s 99200 29112 100000 29232 6 io_wbs_m2s_addr[5]
port 52 nsew signal input
rlabel metal3 s 99200 36048 100000 36168 6 io_wbs_m2s_addr[6]
port 53 nsew signal input
rlabel metal2 s 41602 99200 41658 100000 6 io_wbs_m2s_addr[7]
port 54 nsew signal input
rlabel metal2 s 45006 99200 45062 100000 6 io_wbs_m2s_addr[8]
port 55 nsew signal input
rlabel metal3 s 99200 49784 100000 49904 6 io_wbs_m2s_addr[9]
port 56 nsew signal input
rlabel metal2 s 14922 99200 14978 100000 6 io_wbs_m2s_data[0]
port 57 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 io_wbs_m2s_data[10]
port 58 nsew signal input
rlabel metal2 s 51630 99200 51686 100000 6 io_wbs_m2s_data[11]
port 59 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 io_wbs_m2s_data[12]
port 60 nsew signal input
rlabel metal3 s 99200 60120 100000 60240 6 io_wbs_m2s_data[13]
port 61 nsew signal input
rlabel metal2 s 64970 99200 65026 100000 6 io_wbs_m2s_data[14]
port 62 nsew signal input
rlabel metal3 s 99200 63656 100000 63776 6 io_wbs_m2s_data[15]
port 63 nsew signal input
rlabel metal2 s 71594 99200 71650 100000 6 io_wbs_m2s_data[16]
port 64 nsew signal input
rlabel metal2 s 74998 99200 75054 100000 6 io_wbs_m2s_data[17]
port 65 nsew signal input
rlabel metal3 s 99200 70456 100000 70576 6 io_wbs_m2s_data[18]
port 66 nsew signal input
rlabel metal3 s 99200 73992 100000 74112 6 io_wbs_m2s_data[19]
port 67 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 io_wbs_m2s_data[1]
port 68 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 io_wbs_m2s_data[20]
port 69 nsew signal input
rlabel metal3 s 99200 77392 100000 77512 6 io_wbs_m2s_data[21]
port 70 nsew signal input
rlabel metal2 s 81622 99200 81678 100000 6 io_wbs_m2s_data[22]
port 71 nsew signal input
rlabel metal2 s 84934 99200 84990 100000 6 io_wbs_m2s_data[23]
port 72 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 io_wbs_m2s_data[24]
port 73 nsew signal input
rlabel metal3 s 99200 80792 100000 80912 6 io_wbs_m2s_data[25]
port 74 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 io_wbs_m2s_data[26]
port 75 nsew signal input
rlabel metal3 s 99200 87728 100000 87848 6 io_wbs_m2s_data[27]
port 76 nsew signal input
rlabel metal3 s 99200 91128 100000 91248 6 io_wbs_m2s_data[28]
port 77 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 io_wbs_m2s_data[29]
port 78 nsew signal input
rlabel metal3 s 99200 25712 100000 25832 6 io_wbs_m2s_data[2]
port 79 nsew signal input
rlabel metal2 s 98274 99200 98330 100000 6 io_wbs_m2s_data[30]
port 80 nsew signal input
rlabel metal3 s 99200 98064 100000 98184 6 io_wbs_m2s_data[31]
port 81 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 io_wbs_m2s_data[3]
port 82 nsew signal input
rlabel metal2 s 34978 99200 35034 100000 6 io_wbs_m2s_data[4]
port 83 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 io_wbs_m2s_data[5]
port 84 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 io_wbs_m2s_data[6]
port 85 nsew signal input
rlabel metal3 s 99200 39448 100000 39568 6 io_wbs_m2s_data[7]
port 86 nsew signal input
rlabel metal3 s 99200 42984 100000 43104 6 io_wbs_m2s_data[8]
port 87 nsew signal input
rlabel metal2 s 48318 99200 48374 100000 6 io_wbs_m2s_data[9]
port 88 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 io_wbs_m2s_sel[0]
port 89 nsew signal input
rlabel metal3 s 99200 22312 100000 22432 6 io_wbs_m2s_sel[1]
port 90 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 io_wbs_m2s_sel[2]
port 91 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 io_wbs_m2s_sel[3]
port 92 nsew signal input
rlabel metal3 s 99200 8440 100000 8560 6 io_wbs_m2s_stb
port 93 nsew signal input
rlabel metal3 s 99200 11976 100000 12096 6 io_wbs_m2s_we
port 94 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 reset
port 95 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 97 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 97 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 97 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17432058
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/Motor_Top/runs/Motor_Top/results/finishing/Motor_Top.magic.gds
string GDS_START 1020774
<< end >>

