magic
tech sky130A
magscale 1 2
timestamp 1647505418
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 1104 2128 28888 27792
<< metal2 >>
rect 662 29200 718 30000
rect 1306 29200 1362 30000
rect 2594 29200 2650 30000
rect 3882 29200 3938 30000
rect 4526 29200 4582 30000
rect 5814 29200 5870 30000
rect 7102 29200 7158 30000
rect 8390 29200 8446 30000
rect 9034 29200 9090 30000
rect 10322 29200 10378 30000
rect 11610 29200 11666 30000
rect 12898 29200 12954 30000
rect 13542 29200 13598 30000
rect 14830 29200 14886 30000
rect 16118 29200 16174 30000
rect 17406 29200 17462 30000
rect 18050 29200 18106 30000
rect 19338 29200 19394 30000
rect 20626 29200 20682 30000
rect 21270 29200 21326 30000
rect 22558 29200 22614 30000
rect 23846 29200 23902 30000
rect 25134 29200 25190 30000
rect 25778 29200 25834 30000
rect 27066 29200 27122 30000
rect 28354 29200 28410 30000
rect 29642 29200 29698 30000
rect 18 0 74 800
rect 662 0 718 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 28998 0 29054 800
rect 29642 0 29698 800
<< obsm2 >>
rect 1418 29144 2538 29345
rect 2706 29144 3826 29345
rect 3994 29144 4470 29345
rect 4638 29144 5758 29345
rect 5926 29144 7046 29345
rect 7214 29144 8334 29345
rect 8502 29144 8978 29345
rect 9146 29144 10266 29345
rect 10434 29144 11554 29345
rect 11722 29144 12842 29345
rect 13010 29144 13486 29345
rect 13654 29144 14774 29345
rect 14942 29144 16062 29345
rect 16230 29144 17350 29345
rect 17518 29144 17994 29345
rect 18162 29144 19282 29345
rect 19450 29144 20570 29345
rect 20738 29144 21214 29345
rect 21382 29144 22502 29345
rect 22670 29144 23790 29345
rect 23958 29144 25078 29345
rect 25246 29144 25722 29345
rect 25890 29144 27010 29345
rect 27178 29144 28298 29345
rect 1398 856 28410 29144
rect 1398 711 1894 856
rect 2062 711 3182 856
rect 3350 711 3826 856
rect 3994 711 5114 856
rect 5282 711 6402 856
rect 6570 711 7690 856
rect 7858 711 8334 856
rect 8502 711 9622 856
rect 9790 711 10910 856
rect 11078 711 12198 856
rect 12366 711 12842 856
rect 13010 711 14130 856
rect 14298 711 15418 856
rect 15586 711 16706 856
rect 16874 711 17350 856
rect 17518 711 18638 856
rect 18806 711 19926 856
rect 20094 711 20570 856
rect 20738 711 21858 856
rect 22026 711 23146 856
rect 23314 711 24434 856
rect 24602 711 25078 856
rect 25246 711 26366 856
rect 26534 711 27654 856
rect 27822 711 28410 856
<< metal3 >>
rect 0 29248 800 29368
rect 29200 29248 30000 29368
rect 0 27888 800 28008
rect 29200 27888 30000 28008
rect 0 26528 800 26648
rect 29200 26528 30000 26648
rect 0 25848 800 25968
rect 29200 25168 30000 25288
rect 0 24488 800 24608
rect 29200 24488 30000 24608
rect 0 23128 800 23248
rect 29200 23128 30000 23248
rect 0 21768 800 21888
rect 29200 21768 30000 21888
rect 0 21088 800 21208
rect 29200 21088 30000 21208
rect 0 19728 800 19848
rect 29200 19728 30000 19848
rect 0 18368 800 18488
rect 29200 18368 30000 18488
rect 0 17008 800 17128
rect 29200 17008 30000 17128
rect 0 16328 800 16448
rect 29200 16328 30000 16448
rect 0 14968 800 15088
rect 29200 14968 30000 15088
rect 0 13608 800 13728
rect 29200 13608 30000 13728
rect 0 12928 800 13048
rect 29200 12248 30000 12368
rect 0 11568 800 11688
rect 29200 11568 30000 11688
rect 0 10208 800 10328
rect 29200 10208 30000 10328
rect 0 8848 800 8968
rect 29200 8848 30000 8968
rect 0 8168 800 8288
rect 29200 7488 30000 7608
rect 0 6808 800 6928
rect 29200 6808 30000 6928
rect 0 5448 800 5568
rect 29200 5448 30000 5568
rect 0 4088 800 4208
rect 29200 4088 30000 4208
rect 0 3408 800 3528
rect 29200 3408 30000 3528
rect 0 2048 800 2168
rect 29200 2048 30000 2168
rect 0 688 800 808
rect 29200 688 30000 808
<< obsm3 >>
rect 880 29168 29120 29341
rect 800 28088 29200 29168
rect 880 27808 29120 28088
rect 800 26728 29200 27808
rect 880 26448 29120 26728
rect 800 26048 29200 26448
rect 880 25768 29200 26048
rect 800 25368 29200 25768
rect 800 25088 29120 25368
rect 800 24688 29200 25088
rect 880 24408 29120 24688
rect 800 23328 29200 24408
rect 880 23048 29120 23328
rect 800 21968 29200 23048
rect 880 21688 29120 21968
rect 800 21288 29200 21688
rect 880 21008 29120 21288
rect 800 19928 29200 21008
rect 880 19648 29120 19928
rect 800 18568 29200 19648
rect 880 18288 29120 18568
rect 800 17208 29200 18288
rect 880 16928 29120 17208
rect 800 16528 29200 16928
rect 880 16248 29120 16528
rect 800 15168 29200 16248
rect 880 14888 29120 15168
rect 800 13808 29200 14888
rect 880 13528 29120 13808
rect 800 13128 29200 13528
rect 880 12848 29200 13128
rect 800 12448 29200 12848
rect 800 12168 29120 12448
rect 800 11768 29200 12168
rect 880 11488 29120 11768
rect 800 10408 29200 11488
rect 880 10128 29120 10408
rect 800 9048 29200 10128
rect 880 8768 29120 9048
rect 800 8368 29200 8768
rect 880 8088 29200 8368
rect 800 7688 29200 8088
rect 800 7408 29120 7688
rect 800 7008 29200 7408
rect 880 6728 29120 7008
rect 800 5648 29200 6728
rect 880 5368 29120 5648
rect 800 4288 29200 5368
rect 880 4008 29120 4288
rect 800 3608 29200 4008
rect 880 3328 29120 3608
rect 800 2248 29200 3328
rect 880 1968 29120 2248
rect 800 888 29200 1968
rect 880 715 29120 888
<< metal4 >>
rect 5576 2128 5896 27792
rect 10208 2128 10528 27792
rect 14840 2128 15160 27792
rect 19472 2128 19792 27792
rect 24104 2128 24424 27792
<< obsm4 >>
rect 11099 3435 14760 21317
rect 15240 3435 19392 21317
rect 19872 3435 21101 21317
<< labels >>
rlabel metal2 s 9034 29200 9090 30000 6 clock
port 1 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 io_rxd
port 2 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 io_txd
port 3 nsew signal output
rlabel metal2 s 16118 29200 16174 30000 6 io_uartInt
port 4 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 io_uart_select
port 5 nsew signal input
rlabel metal3 s 29200 10208 30000 10328 6 io_wbs_ack_o
port 6 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 io_wbs_data_o[0]
port 7 nsew signal output
rlabel metal2 s 19338 29200 19394 30000 6 io_wbs_data_o[10]
port 8 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 io_wbs_data_o[11]
port 9 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 io_wbs_data_o[12]
port 10 nsew signal output
rlabel metal3 s 29200 23128 30000 23248 6 io_wbs_data_o[13]
port 11 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 io_wbs_data_o[14]
port 12 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 io_wbs_data_o[15]
port 13 nsew signal output
rlabel metal3 s 29200 5448 30000 5568 6 io_wbs_data_o[16]
port 14 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 io_wbs_data_o[17]
port 15 nsew signal output
rlabel metal3 s 29200 14968 30000 15088 6 io_wbs_data_o[18]
port 16 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 io_wbs_data_o[19]
port 17 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 io_wbs_data_o[1]
port 18 nsew signal output
rlabel metal2 s 25778 29200 25834 30000 6 io_wbs_data_o[20]
port 19 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 io_wbs_data_o[21]
port 20 nsew signal output
rlabel metal3 s 29200 4088 30000 4208 6 io_wbs_data_o[22]
port 21 nsew signal output
rlabel metal3 s 29200 16328 30000 16448 6 io_wbs_data_o[23]
port 22 nsew signal output
rlabel metal3 s 29200 26528 30000 26648 6 io_wbs_data_o[24]
port 23 nsew signal output
rlabel metal2 s 3882 29200 3938 30000 6 io_wbs_data_o[25]
port 24 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 io_wbs_data_o[26]
port 25 nsew signal output
rlabel metal2 s 21270 29200 21326 30000 6 io_wbs_data_o[27]
port 26 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 io_wbs_data_o[28]
port 27 nsew signal output
rlabel metal2 s 28354 29200 28410 30000 6 io_wbs_data_o[29]
port 28 nsew signal output
rlabel metal3 s 29200 27888 30000 28008 6 io_wbs_data_o[2]
port 29 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 io_wbs_data_o[30]
port 30 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 io_wbs_data_o[31]
port 31 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 io_wbs_data_o[3]
port 32 nsew signal output
rlabel metal3 s 29200 29248 30000 29368 6 io_wbs_data_o[4]
port 33 nsew signal output
rlabel metal2 s 25134 29200 25190 30000 6 io_wbs_data_o[5]
port 34 nsew signal output
rlabel metal3 s 29200 688 30000 808 6 io_wbs_data_o[6]
port 35 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_wbs_data_o[7]
port 36 nsew signal output
rlabel metal3 s 29200 12248 30000 12368 6 io_wbs_data_o[8]
port 37 nsew signal output
rlabel metal3 s 29200 8848 30000 8968 6 io_wbs_data_o[9]
port 38 nsew signal output
rlabel metal2 s 10322 29200 10378 30000 6 io_wbs_m2s_addr[0]
port 39 nsew signal input
rlabel metal2 s 11610 29200 11666 30000 6 io_wbs_m2s_addr[10]
port 40 nsew signal input
rlabel metal3 s 29200 21768 30000 21888 6 io_wbs_m2s_addr[11]
port 41 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 io_wbs_m2s_addr[12]
port 42 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 io_wbs_m2s_addr[13]
port 43 nsew signal input
rlabel metal3 s 29200 24488 30000 24608 6 io_wbs_m2s_addr[14]
port 44 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 io_wbs_m2s_addr[15]
port 45 nsew signal input
rlabel metal2 s 17406 29200 17462 30000 6 io_wbs_m2s_addr[16]
port 46 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 io_wbs_m2s_addr[17]
port 47 nsew signal input
rlabel metal2 s 8390 29200 8446 30000 6 io_wbs_m2s_addr[18]
port 48 nsew signal input
rlabel metal2 s 12898 29200 12954 30000 6 io_wbs_m2s_addr[19]
port 49 nsew signal input
rlabel metal3 s 29200 25168 30000 25288 6 io_wbs_m2s_addr[1]
port 50 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 io_wbs_m2s_addr[20]
port 51 nsew signal input
rlabel metal2 s 14830 29200 14886 30000 6 io_wbs_m2s_addr[21]
port 52 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 io_wbs_m2s_addr[22]
port 53 nsew signal input
rlabel metal3 s 29200 6808 30000 6928 6 io_wbs_m2s_addr[23]
port 54 nsew signal input
rlabel metal3 s 29200 18368 30000 18488 6 io_wbs_m2s_addr[24]
port 55 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 io_wbs_m2s_addr[25]
port 56 nsew signal input
rlabel metal2 s 18050 29200 18106 30000 6 io_wbs_m2s_addr[26]
port 57 nsew signal input
rlabel metal2 s 5814 29200 5870 30000 6 io_wbs_m2s_addr[27]
port 58 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 io_wbs_m2s_addr[28]
port 59 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 io_wbs_m2s_addr[29]
port 60 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 io_wbs_m2s_addr[2]
port 61 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 io_wbs_m2s_addr[30]
port 62 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_wbs_m2s_addr[31]
port 63 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 io_wbs_m2s_addr[3]
port 64 nsew signal input
rlabel metal3 s 0 688 800 808 6 io_wbs_m2s_addr[4]
port 65 nsew signal input
rlabel metal3 s 29200 7488 30000 7608 6 io_wbs_m2s_addr[5]
port 66 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 io_wbs_m2s_addr[6]
port 67 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_wbs_m2s_addr[7]
port 68 nsew signal input
rlabel metal3 s 29200 2048 30000 2168 6 io_wbs_m2s_addr[8]
port 69 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 io_wbs_m2s_addr[9]
port 70 nsew signal input
rlabel metal3 s 29200 11568 30000 11688 6 io_wbs_m2s_data[0]
port 71 nsew signal input
rlabel metal3 s 29200 19728 30000 19848 6 io_wbs_m2s_data[10]
port 72 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 io_wbs_m2s_data[11]
port 73 nsew signal input
rlabel metal3 s 29200 21088 30000 21208 6 io_wbs_m2s_data[12]
port 74 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_wbs_m2s_data[13]
port 75 nsew signal input
rlabel metal2 s 662 29200 718 30000 6 io_wbs_m2s_data[14]
port 76 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 io_wbs_m2s_data[15]
port 77 nsew signal input
rlabel metal2 s 18 0 74 800 6 io_wbs_m2s_data[16]
port 78 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 io_wbs_m2s_data[17]
port 79 nsew signal input
rlabel metal2 s 4526 29200 4582 30000 6 io_wbs_m2s_data[18]
port 80 nsew signal input
rlabel metal2 s 13542 29200 13598 30000 6 io_wbs_m2s_data[19]
port 81 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 io_wbs_m2s_data[1]
port 82 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 io_wbs_m2s_data[20]
port 83 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 io_wbs_m2s_data[21]
port 84 nsew signal input
rlabel metal2 s 662 0 718 800 6 io_wbs_m2s_data[22]
port 85 nsew signal input
rlabel metal2 s 27066 29200 27122 30000 6 io_wbs_m2s_data[23]
port 86 nsew signal input
rlabel metal2 s 20626 29200 20682 30000 6 io_wbs_m2s_data[24]
port 87 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 io_wbs_m2s_data[25]
port 88 nsew signal input
rlabel metal2 s 29642 29200 29698 30000 6 io_wbs_m2s_data[26]
port 89 nsew signal input
rlabel metal3 s 29200 3408 30000 3528 6 io_wbs_m2s_data[27]
port 90 nsew signal input
rlabel metal2 s 1306 29200 1362 30000 6 io_wbs_m2s_data[28]
port 91 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 io_wbs_m2s_data[29]
port 92 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 io_wbs_m2s_data[2]
port 93 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 io_wbs_m2s_data[30]
port 94 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 io_wbs_m2s_data[31]
port 95 nsew signal input
rlabel metal3 s 29200 17008 30000 17128 6 io_wbs_m2s_data[3]
port 96 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_wbs_m2s_data[4]
port 97 nsew signal input
rlabel metal2 s 23846 29200 23902 30000 6 io_wbs_m2s_data[5]
port 98 nsew signal input
rlabel metal2 s 22558 29200 22614 30000 6 io_wbs_m2s_data[6]
port 99 nsew signal input
rlabel metal2 s 2594 29200 2650 30000 6 io_wbs_m2s_data[7]
port 100 nsew signal input
rlabel metal2 s 7102 29200 7158 30000 6 io_wbs_m2s_data[8]
port 101 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 io_wbs_m2s_data[9]
port 102 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 io_wbs_m2s_stb
port 103 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 io_wbs_m2s_we
port 104 nsew signal input
rlabel metal3 s 29200 13608 30000 13728 6 reset
port 105 nsew signal input
rlabel metal4 s 5576 2128 5896 27792 6 vccd1
port 106 nsew power input
rlabel metal4 s 14840 2128 15160 27792 6 vccd1
port 106 nsew power input
rlabel metal4 s 24104 2128 24424 27792 6 vccd1
port 106 nsew power input
rlabel metal4 s 10208 2128 10528 27792 6 vssd1
port 107 nsew ground input
rlabel metal4 s 19472 2128 19792 27792 6 vssd1
port 107 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2221828
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/UART/runs/UART/results/finishing/UART.magic.gds
string GDS_START 408722
<< end >>

