IntxLNK/ h o m e / a l i 1 1 2 0 0 0 / D e s k t o p / m p w / p d k / o p e n _ p d k s / s o u r c e s / s k y 1 3 0 _ s r a m _ m a c r o s / s k y 1 3 0 _ s r a m _ 2 k b y t e _ 1 r w 1 r _ 3 2 x 5 1 2 _ 8 / s k y 1 3 0 _ s r a m _ 2 k b y t e _ 1 r w 1 r _ 3 2 x 5 1 2 _ 8 . l e f 