VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO UART
  CLASS BLOCK ;
  FOREIGN UART ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 146.000 45.450 150.000 ;
    END
  END clock
  PIN io_rxd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END io_rxd
  PIN io_txd
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END io_txd
  PIN io_uartInt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 146.000 80.870 150.000 ;
    END
  END io_uartInt
  PIN io_uart_select
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_uart_select
  PIN io_wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 51.040 150.000 51.640 ;
    END
  END io_wbs_ack_o
  PIN io_wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END io_wbs_data_o[0]
  PIN io_wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 146.000 96.970 150.000 ;
    END
  END io_wbs_data_o[10]
  PIN io_wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END io_wbs_data_o[11]
  PIN io_wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END io_wbs_data_o[12]
  PIN io_wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 115.640 150.000 116.240 ;
    END
  END io_wbs_data_o[13]
  PIN io_wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END io_wbs_data_o[14]
  PIN io_wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END io_wbs_data_o[15]
  PIN io_wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 27.240 150.000 27.840 ;
    END
  END io_wbs_data_o[16]
  PIN io_wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_wbs_data_o[17]
  PIN io_wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.840 150.000 75.440 ;
    END
  END io_wbs_data_o[18]
  PIN io_wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_wbs_data_o[19]
  PIN io_wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END io_wbs_data_o[1]
  PIN io_wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 146.000 129.170 150.000 ;
    END
  END io_wbs_data_o[20]
  PIN io_wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END io_wbs_data_o[21]
  PIN io_wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 20.440 150.000 21.040 ;
    END
  END io_wbs_data_o[22]
  PIN io_wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 81.640 150.000 82.240 ;
    END
  END io_wbs_data_o[23]
  PIN io_wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 132.640 150.000 133.240 ;
    END
  END io_wbs_data_o[24]
  PIN io_wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 146.000 19.690 150.000 ;
    END
  END io_wbs_data_o[25]
  PIN io_wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END io_wbs_data_o[26]
  PIN io_wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 146.000 106.630 150.000 ;
    END
  END io_wbs_data_o[27]
  PIN io_wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END io_wbs_data_o[28]
  PIN io_wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 146.000 142.050 150.000 ;
    END
  END io_wbs_data_o[29]
  PIN io_wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 139.440 150.000 140.040 ;
    END
  END io_wbs_data_o[2]
  PIN io_wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_wbs_data_o[30]
  PIN io_wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END io_wbs_data_o[31]
  PIN io_wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_wbs_data_o[3]
  PIN io_wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 146.240 150.000 146.840 ;
    END
  END io_wbs_data_o[4]
  PIN io_wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 146.000 125.950 150.000 ;
    END
  END io_wbs_data_o[5]
  PIN io_wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 3.440 150.000 4.040 ;
    END
  END io_wbs_data_o[6]
  PIN io_wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_wbs_data_o[7]
  PIN io_wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 61.240 150.000 61.840 ;
    END
  END io_wbs_data_o[8]
  PIN io_wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 44.240 150.000 44.840 ;
    END
  END io_wbs_data_o[9]
  PIN io_wbs_m2s_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 146.000 51.890 150.000 ;
    END
  END io_wbs_m2s_addr[0]
  PIN io_wbs_m2s_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 146.000 58.330 150.000 ;
    END
  END io_wbs_m2s_addr[10]
  PIN io_wbs_m2s_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 108.840 150.000 109.440 ;
    END
  END io_wbs_m2s_addr[11]
  PIN io_wbs_m2s_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END io_wbs_m2s_addr[12]
  PIN io_wbs_m2s_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END io_wbs_m2s_addr[13]
  PIN io_wbs_m2s_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 122.440 150.000 123.040 ;
    END
  END io_wbs_m2s_addr[14]
  PIN io_wbs_m2s_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END io_wbs_m2s_addr[15]
  PIN io_wbs_m2s_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 146.000 87.310 150.000 ;
    END
  END io_wbs_m2s_addr[16]
  PIN io_wbs_m2s_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END io_wbs_m2s_addr[17]
  PIN io_wbs_m2s_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 146.000 42.230 150.000 ;
    END
  END io_wbs_m2s_addr[18]
  PIN io_wbs_m2s_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 146.000 64.770 150.000 ;
    END
  END io_wbs_m2s_addr[19]
  PIN io_wbs_m2s_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 125.840 150.000 126.440 ;
    END
  END io_wbs_m2s_addr[1]
  PIN io_wbs_m2s_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END io_wbs_m2s_addr[20]
  PIN io_wbs_m2s_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 146.000 74.430 150.000 ;
    END
  END io_wbs_m2s_addr[21]
  PIN io_wbs_m2s_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END io_wbs_m2s_addr[22]
  PIN io_wbs_m2s_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 34.040 150.000 34.640 ;
    END
  END io_wbs_m2s_addr[23]
  PIN io_wbs_m2s_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 91.840 150.000 92.440 ;
    END
  END io_wbs_m2s_addr[24]
  PIN io_wbs_m2s_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END io_wbs_m2s_addr[25]
  PIN io_wbs_m2s_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 146.000 90.530 150.000 ;
    END
  END io_wbs_m2s_addr[26]
  PIN io_wbs_m2s_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 146.000 29.350 150.000 ;
    END
  END io_wbs_m2s_addr[27]
  PIN io_wbs_m2s_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END io_wbs_m2s_addr[28]
  PIN io_wbs_m2s_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END io_wbs_m2s_addr[29]
  PIN io_wbs_m2s_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END io_wbs_m2s_addr[2]
  PIN io_wbs_m2s_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END io_wbs_m2s_addr[30]
  PIN io_wbs_m2s_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_wbs_m2s_addr[31]
  PIN io_wbs_m2s_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END io_wbs_m2s_addr[3]
  PIN io_wbs_m2s_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END io_wbs_m2s_addr[4]
  PIN io_wbs_m2s_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 37.440 150.000 38.040 ;
    END
  END io_wbs_m2s_addr[5]
  PIN io_wbs_m2s_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END io_wbs_m2s_addr[6]
  PIN io_wbs_m2s_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_wbs_m2s_addr[7]
  PIN io_wbs_m2s_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 10.240 150.000 10.840 ;
    END
  END io_wbs_m2s_addr[8]
  PIN io_wbs_m2s_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_wbs_m2s_addr[9]
  PIN io_wbs_m2s_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 57.840 150.000 58.440 ;
    END
  END io_wbs_m2s_data[0]
  PIN io_wbs_m2s_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 98.640 150.000 99.240 ;
    END
  END io_wbs_m2s_data[10]
  PIN io_wbs_m2s_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END io_wbs_m2s_data[11]
  PIN io_wbs_m2s_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 105.440 150.000 106.040 ;
    END
  END io_wbs_m2s_data[12]
  PIN io_wbs_m2s_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END io_wbs_m2s_data[13]
  PIN io_wbs_m2s_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 146.000 3.590 150.000 ;
    END
  END io_wbs_m2s_data[14]
  PIN io_wbs_m2s_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_wbs_m2s_data[15]
  PIN io_wbs_m2s_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_wbs_m2s_data[16]
  PIN io_wbs_m2s_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END io_wbs_m2s_data[17]
  PIN io_wbs_m2s_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 146.000 22.910 150.000 ;
    END
  END io_wbs_m2s_data[18]
  PIN io_wbs_m2s_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 146.000 67.990 150.000 ;
    END
  END io_wbs_m2s_data[19]
  PIN io_wbs_m2s_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END io_wbs_m2s_data[1]
  PIN io_wbs_m2s_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_wbs_m2s_data[20]
  PIN io_wbs_m2s_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END io_wbs_m2s_data[21]
  PIN io_wbs_m2s_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END io_wbs_m2s_data[22]
  PIN io_wbs_m2s_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 146.000 135.610 150.000 ;
    END
  END io_wbs_m2s_data[23]
  PIN io_wbs_m2s_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 146.000 103.410 150.000 ;
    END
  END io_wbs_m2s_data[24]
  PIN io_wbs_m2s_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END io_wbs_m2s_data[25]
  PIN io_wbs_m2s_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 146.000 148.490 150.000 ;
    END
  END io_wbs_m2s_data[26]
  PIN io_wbs_m2s_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 17.040 150.000 17.640 ;
    END
  END io_wbs_m2s_data[27]
  PIN io_wbs_m2s_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 146.000 6.810 150.000 ;
    END
  END io_wbs_m2s_data[28]
  PIN io_wbs_m2s_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_wbs_m2s_data[29]
  PIN io_wbs_m2s_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END io_wbs_m2s_data[2]
  PIN io_wbs_m2s_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END io_wbs_m2s_data[30]
  PIN io_wbs_m2s_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END io_wbs_m2s_data[31]
  PIN io_wbs_m2s_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 85.040 150.000 85.640 ;
    END
  END io_wbs_m2s_data[3]
  PIN io_wbs_m2s_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END io_wbs_m2s_data[4]
  PIN io_wbs_m2s_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 146.000 119.510 150.000 ;
    END
  END io_wbs_m2s_data[5]
  PIN io_wbs_m2s_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 146.000 113.070 150.000 ;
    END
  END io_wbs_m2s_data[6]
  PIN io_wbs_m2s_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 146.000 13.250 150.000 ;
    END
  END io_wbs_m2s_data[7]
  PIN io_wbs_m2s_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 146.000 35.790 150.000 ;
    END
  END io_wbs_m2s_data[8]
  PIN io_wbs_m2s_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END io_wbs_m2s_data[9]
  PIN io_wbs_m2s_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END io_wbs_m2s_stb
  PIN io_wbs_m2s_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END io_wbs_m2s_we
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 68.040 150.000 68.640 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.880 10.640 29.480 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.200 10.640 75.800 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.520 10.640 122.120 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.360 10.640 98.960 138.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 144.440 138.960 ;
      LAYER met2 ;
        RECT 7.090 145.720 12.690 146.725 ;
        RECT 13.530 145.720 19.130 146.725 ;
        RECT 19.970 145.720 22.350 146.725 ;
        RECT 23.190 145.720 28.790 146.725 ;
        RECT 29.630 145.720 35.230 146.725 ;
        RECT 36.070 145.720 41.670 146.725 ;
        RECT 42.510 145.720 44.890 146.725 ;
        RECT 45.730 145.720 51.330 146.725 ;
        RECT 52.170 145.720 57.770 146.725 ;
        RECT 58.610 145.720 64.210 146.725 ;
        RECT 65.050 145.720 67.430 146.725 ;
        RECT 68.270 145.720 73.870 146.725 ;
        RECT 74.710 145.720 80.310 146.725 ;
        RECT 81.150 145.720 86.750 146.725 ;
        RECT 87.590 145.720 89.970 146.725 ;
        RECT 90.810 145.720 96.410 146.725 ;
        RECT 97.250 145.720 102.850 146.725 ;
        RECT 103.690 145.720 106.070 146.725 ;
        RECT 106.910 145.720 112.510 146.725 ;
        RECT 113.350 145.720 118.950 146.725 ;
        RECT 119.790 145.720 125.390 146.725 ;
        RECT 126.230 145.720 128.610 146.725 ;
        RECT 129.450 145.720 135.050 146.725 ;
        RECT 135.890 145.720 141.490 146.725 ;
        RECT 6.990 4.280 142.050 145.720 ;
        RECT 6.990 3.555 9.470 4.280 ;
        RECT 10.310 3.555 15.910 4.280 ;
        RECT 16.750 3.555 19.130 4.280 ;
        RECT 19.970 3.555 25.570 4.280 ;
        RECT 26.410 3.555 32.010 4.280 ;
        RECT 32.850 3.555 38.450 4.280 ;
        RECT 39.290 3.555 41.670 4.280 ;
        RECT 42.510 3.555 48.110 4.280 ;
        RECT 48.950 3.555 54.550 4.280 ;
        RECT 55.390 3.555 60.990 4.280 ;
        RECT 61.830 3.555 64.210 4.280 ;
        RECT 65.050 3.555 70.650 4.280 ;
        RECT 71.490 3.555 77.090 4.280 ;
        RECT 77.930 3.555 83.530 4.280 ;
        RECT 84.370 3.555 86.750 4.280 ;
        RECT 87.590 3.555 93.190 4.280 ;
        RECT 94.030 3.555 99.630 4.280 ;
        RECT 100.470 3.555 102.850 4.280 ;
        RECT 103.690 3.555 109.290 4.280 ;
        RECT 110.130 3.555 115.730 4.280 ;
        RECT 116.570 3.555 122.170 4.280 ;
        RECT 123.010 3.555 125.390 4.280 ;
        RECT 126.230 3.555 131.830 4.280 ;
        RECT 132.670 3.555 138.270 4.280 ;
        RECT 139.110 3.555 142.050 4.280 ;
      LAYER met3 ;
        RECT 4.400 145.840 145.600 146.705 ;
        RECT 4.000 140.440 146.000 145.840 ;
        RECT 4.400 139.040 145.600 140.440 ;
        RECT 4.000 133.640 146.000 139.040 ;
        RECT 4.400 132.240 145.600 133.640 ;
        RECT 4.000 130.240 146.000 132.240 ;
        RECT 4.400 128.840 146.000 130.240 ;
        RECT 4.000 126.840 146.000 128.840 ;
        RECT 4.000 125.440 145.600 126.840 ;
        RECT 4.000 123.440 146.000 125.440 ;
        RECT 4.400 122.040 145.600 123.440 ;
        RECT 4.000 116.640 146.000 122.040 ;
        RECT 4.400 115.240 145.600 116.640 ;
        RECT 4.000 109.840 146.000 115.240 ;
        RECT 4.400 108.440 145.600 109.840 ;
        RECT 4.000 106.440 146.000 108.440 ;
        RECT 4.400 105.040 145.600 106.440 ;
        RECT 4.000 99.640 146.000 105.040 ;
        RECT 4.400 98.240 145.600 99.640 ;
        RECT 4.000 92.840 146.000 98.240 ;
        RECT 4.400 91.440 145.600 92.840 ;
        RECT 4.000 86.040 146.000 91.440 ;
        RECT 4.400 84.640 145.600 86.040 ;
        RECT 4.000 82.640 146.000 84.640 ;
        RECT 4.400 81.240 145.600 82.640 ;
        RECT 4.000 75.840 146.000 81.240 ;
        RECT 4.400 74.440 145.600 75.840 ;
        RECT 4.000 69.040 146.000 74.440 ;
        RECT 4.400 67.640 145.600 69.040 ;
        RECT 4.000 65.640 146.000 67.640 ;
        RECT 4.400 64.240 146.000 65.640 ;
        RECT 4.000 62.240 146.000 64.240 ;
        RECT 4.000 60.840 145.600 62.240 ;
        RECT 4.000 58.840 146.000 60.840 ;
        RECT 4.400 57.440 145.600 58.840 ;
        RECT 4.000 52.040 146.000 57.440 ;
        RECT 4.400 50.640 145.600 52.040 ;
        RECT 4.000 45.240 146.000 50.640 ;
        RECT 4.400 43.840 145.600 45.240 ;
        RECT 4.000 41.840 146.000 43.840 ;
        RECT 4.400 40.440 146.000 41.840 ;
        RECT 4.000 38.440 146.000 40.440 ;
        RECT 4.000 37.040 145.600 38.440 ;
        RECT 4.000 35.040 146.000 37.040 ;
        RECT 4.400 33.640 145.600 35.040 ;
        RECT 4.000 28.240 146.000 33.640 ;
        RECT 4.400 26.840 145.600 28.240 ;
        RECT 4.000 21.440 146.000 26.840 ;
        RECT 4.400 20.040 145.600 21.440 ;
        RECT 4.000 18.040 146.000 20.040 ;
        RECT 4.400 16.640 145.600 18.040 ;
        RECT 4.000 11.240 146.000 16.640 ;
        RECT 4.400 9.840 145.600 11.240 ;
        RECT 4.000 4.440 146.000 9.840 ;
        RECT 4.400 3.575 145.600 4.440 ;
      LAYER met4 ;
        RECT 55.495 17.175 73.800 106.585 ;
        RECT 76.200 17.175 96.960 106.585 ;
        RECT 99.360 17.175 105.505 106.585 ;
  END
END UART
END LIBRARY

