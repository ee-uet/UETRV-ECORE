magic
tech sky130A
magscale 1 2
timestamp 1647678698
<< obsli1 >>
rect 1104 2159 78844 77809
<< obsm1 >>
rect 1104 1980 78844 77840
<< metal2 >>
rect 1766 79200 1822 80000
rect 5354 79200 5410 80000
rect 9034 79200 9090 80000
rect 12622 79200 12678 80000
rect 16302 79200 16358 80000
rect 19890 79200 19946 80000
rect 23570 79200 23626 80000
rect 27158 79200 27214 80000
rect 30838 79200 30894 80000
rect 34426 79200 34482 80000
rect 38106 79200 38162 80000
rect 41786 79200 41842 80000
rect 45374 79200 45430 80000
rect 49054 79200 49110 80000
rect 52642 79200 52698 80000
rect 56322 79200 56378 80000
rect 59910 79200 59966 80000
rect 63590 79200 63646 80000
rect 67178 79200 67234 80000
rect 70858 79200 70914 80000
rect 74446 79200 74502 80000
rect 78126 79200 78182 80000
rect 1674 0 1730 800
rect 4986 0 5042 800
rect 8298 0 8354 800
rect 11610 0 11666 800
rect 15014 0 15070 800
rect 18326 0 18382 800
rect 21638 0 21694 800
rect 24950 0 25006 800
rect 28354 0 28410 800
rect 31666 0 31722 800
rect 34978 0 35034 800
rect 38290 0 38346 800
rect 41694 0 41750 800
rect 45006 0 45062 800
rect 48318 0 48374 800
rect 51630 0 51686 800
rect 55034 0 55090 800
rect 58346 0 58402 800
rect 61658 0 61714 800
rect 64970 0 65026 800
rect 68374 0 68430 800
rect 71686 0 71742 800
rect 74998 0 75054 800
rect 78310 0 78366 800
<< obsm2 >>
rect 1398 79144 1710 79200
rect 1878 79144 5298 79200
rect 5466 79144 8978 79200
rect 9146 79144 12566 79200
rect 12734 79144 16246 79200
rect 16414 79144 19834 79200
rect 20002 79144 23514 79200
rect 23682 79144 27102 79200
rect 27270 79144 30782 79200
rect 30950 79144 34370 79200
rect 34538 79144 38050 79200
rect 38218 79144 41730 79200
rect 41898 79144 45318 79200
rect 45486 79144 48998 79200
rect 49166 79144 52586 79200
rect 52754 79144 56266 79200
rect 56434 79144 59854 79200
rect 60022 79144 63534 79200
rect 63702 79144 67122 79200
rect 67290 79144 70802 79200
rect 70970 79144 74390 79200
rect 74558 79144 78070 79200
rect 78238 79144 78366 79200
rect 1398 856 78366 79144
rect 1398 734 1618 856
rect 1786 734 4930 856
rect 5098 734 8242 856
rect 8410 734 11554 856
rect 11722 734 14958 856
rect 15126 734 18270 856
rect 18438 734 21582 856
rect 21750 734 24894 856
rect 25062 734 28298 856
rect 28466 734 31610 856
rect 31778 734 34922 856
rect 35090 734 38234 856
rect 38402 734 41638 856
rect 41806 734 44950 856
rect 45118 734 48262 856
rect 48430 734 51574 856
rect 51742 734 54978 856
rect 55146 734 58290 856
rect 58458 734 61602 856
rect 61770 734 64914 856
rect 65082 734 68318 856
rect 68486 734 71630 856
rect 71798 734 74942 856
rect 75110 734 78254 856
<< metal3 >>
rect 0 78344 800 78464
rect 79200 78072 80000 78192
rect 0 75216 800 75336
rect 79200 74536 80000 74656
rect 0 72224 800 72344
rect 79200 71136 80000 71256
rect 0 69096 800 69216
rect 79200 67600 80000 67720
rect 0 65968 800 66088
rect 79200 64200 80000 64320
rect 0 62976 800 63096
rect 79200 60664 80000 60784
rect 0 59848 800 59968
rect 79200 57264 80000 57384
rect 0 56856 800 56976
rect 0 53728 800 53848
rect 79200 53728 80000 53848
rect 0 50600 800 50720
rect 79200 50192 80000 50312
rect 0 47608 800 47728
rect 79200 46792 80000 46912
rect 0 44480 800 44600
rect 79200 43256 80000 43376
rect 0 41488 800 41608
rect 79200 39856 80000 39976
rect 0 38360 800 38480
rect 79200 36320 80000 36440
rect 0 35232 800 35352
rect 79200 32920 80000 33040
rect 0 32240 800 32360
rect 79200 29384 80000 29504
rect 0 29112 800 29232
rect 0 25984 800 26104
rect 79200 25848 80000 25968
rect 0 22992 800 23112
rect 79200 22448 80000 22568
rect 0 19864 800 19984
rect 79200 18912 80000 19032
rect 0 16872 800 16992
rect 79200 15512 80000 15632
rect 0 13744 800 13864
rect 79200 11976 80000 12096
rect 0 10616 800 10736
rect 79200 8576 80000 8696
rect 0 7624 800 7744
rect 79200 5040 80000 5160
rect 0 4496 800 4616
rect 0 1504 800 1624
rect 79200 1640 80000 1760
<< obsm3 >>
rect 880 78272 79200 78437
rect 880 78264 79120 78272
rect 800 77992 79120 78264
rect 800 75416 79200 77992
rect 880 75136 79200 75416
rect 800 74736 79200 75136
rect 800 74456 79120 74736
rect 800 72424 79200 74456
rect 880 72144 79200 72424
rect 800 71336 79200 72144
rect 800 71056 79120 71336
rect 800 69296 79200 71056
rect 880 69016 79200 69296
rect 800 67800 79200 69016
rect 800 67520 79120 67800
rect 800 66168 79200 67520
rect 880 65888 79200 66168
rect 800 64400 79200 65888
rect 800 64120 79120 64400
rect 800 63176 79200 64120
rect 880 62896 79200 63176
rect 800 60864 79200 62896
rect 800 60584 79120 60864
rect 800 60048 79200 60584
rect 880 59768 79200 60048
rect 800 57464 79200 59768
rect 800 57184 79120 57464
rect 800 57056 79200 57184
rect 880 56776 79200 57056
rect 800 53928 79200 56776
rect 880 53648 79120 53928
rect 800 50800 79200 53648
rect 880 50520 79200 50800
rect 800 50392 79200 50520
rect 800 50112 79120 50392
rect 800 47808 79200 50112
rect 880 47528 79200 47808
rect 800 46992 79200 47528
rect 800 46712 79120 46992
rect 800 44680 79200 46712
rect 880 44400 79200 44680
rect 800 43456 79200 44400
rect 800 43176 79120 43456
rect 800 41688 79200 43176
rect 880 41408 79200 41688
rect 800 40056 79200 41408
rect 800 39776 79120 40056
rect 800 38560 79200 39776
rect 880 38280 79200 38560
rect 800 36520 79200 38280
rect 800 36240 79120 36520
rect 800 35432 79200 36240
rect 880 35152 79200 35432
rect 800 33120 79200 35152
rect 800 32840 79120 33120
rect 800 32440 79200 32840
rect 880 32160 79200 32440
rect 800 29584 79200 32160
rect 800 29312 79120 29584
rect 880 29304 79120 29312
rect 880 29032 79200 29304
rect 800 26184 79200 29032
rect 880 26048 79200 26184
rect 880 25904 79120 26048
rect 800 25768 79120 25904
rect 800 23192 79200 25768
rect 880 22912 79200 23192
rect 800 22648 79200 22912
rect 800 22368 79120 22648
rect 800 20064 79200 22368
rect 880 19784 79200 20064
rect 800 19112 79200 19784
rect 800 18832 79120 19112
rect 800 17072 79200 18832
rect 880 16792 79200 17072
rect 800 15712 79200 16792
rect 800 15432 79120 15712
rect 800 13944 79200 15432
rect 880 13664 79200 13944
rect 800 12176 79200 13664
rect 800 11896 79120 12176
rect 800 10816 79200 11896
rect 880 10536 79200 10816
rect 800 8776 79200 10536
rect 800 8496 79120 8776
rect 800 7824 79200 8496
rect 880 7544 79200 7824
rect 800 5240 79200 7544
rect 800 4960 79120 5240
rect 800 4696 79200 4960
rect 880 4416 79200 4696
rect 800 1840 79200 4416
rect 800 1704 79120 1840
rect 880 1560 79120 1704
rect 880 1531 79200 1560
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
<< obsm4 >>
rect 20299 2211 34848 77621
rect 35328 2211 50208 77621
rect 50688 2211 65568 77621
rect 66048 2211 72989 77621
<< labels >>
rlabel metal2 s 1674 0 1730 800 6 clock
port 1 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 io_ba_match
port 2 nsew signal input
rlabel metal3 s 79200 1640 80000 1760 6 io_motor_irq
port 3 nsew signal output
rlabel metal2 s 1766 79200 1822 80000 6 io_pwm_high
port 4 nsew signal output
rlabel metal2 s 5354 79200 5410 80000 6 io_pwm_low
port 5 nsew signal output
rlabel metal3 s 79200 5040 80000 5160 6 io_qei_ch_a
port 6 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 io_qei_ch_b
port 7 nsew signal input
rlabel metal3 s 79200 8576 80000 8696 6 io_wbs_ack_o
port 8 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 io_wbs_data_o[0]
port 9 nsew signal output
rlabel metal2 s 38106 79200 38162 80000 6 io_wbs_data_o[10]
port 10 nsew signal output
rlabel metal3 s 79200 39856 80000 39976 6 io_wbs_data_o[11]
port 11 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 io_wbs_data_o[12]
port 12 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 io_wbs_data_o[13]
port 13 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 io_wbs_data_o[14]
port 14 nsew signal output
rlabel metal3 s 79200 46792 80000 46912 6 io_wbs_data_o[15]
port 15 nsew signal output
rlabel metal2 s 45374 79200 45430 80000 6 io_wbs_data_o[16]
port 16 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 io_wbs_data_o[17]
port 17 nsew signal output
rlabel metal3 s 0 69096 800 69216 6 io_wbs_data_o[18]
port 18 nsew signal output
rlabel metal2 s 52642 79200 52698 80000 6 io_wbs_data_o[19]
port 19 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 io_wbs_data_o[1]
port 20 nsew signal output
rlabel metal3 s 79200 53728 80000 53848 6 io_wbs_data_o[20]
port 21 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 io_wbs_data_o[21]
port 22 nsew signal output
rlabel metal2 s 59910 79200 59966 80000 6 io_wbs_data_o[22]
port 23 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 io_wbs_data_o[23]
port 24 nsew signal output
rlabel metal3 s 79200 64200 80000 64320 6 io_wbs_data_o[24]
port 25 nsew signal output
rlabel metal2 s 67178 79200 67234 80000 6 io_wbs_data_o[25]
port 26 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 io_wbs_data_o[26]
port 27 nsew signal output
rlabel metal3 s 79200 67600 80000 67720 6 io_wbs_data_o[27]
port 28 nsew signal output
rlabel metal3 s 79200 71136 80000 71256 6 io_wbs_data_o[28]
port 29 nsew signal output
rlabel metal3 s 0 75216 800 75336 6 io_wbs_data_o[29]
port 30 nsew signal output
rlabel metal3 s 79200 11976 80000 12096 6 io_wbs_data_o[2]
port 31 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 io_wbs_data_o[30]
port 32 nsew signal output
rlabel metal2 s 78126 79200 78182 80000 6 io_wbs_data_o[31]
port 33 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 io_wbs_data_o[3]
port 34 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 io_wbs_data_o[4]
port 35 nsew signal output
rlabel metal2 s 12622 79200 12678 80000 6 io_wbs_data_o[5]
port 36 nsew signal output
rlabel metal3 s 79200 22448 80000 22568 6 io_wbs_data_o[6]
port 37 nsew signal output
rlabel metal3 s 0 35232 800 35352 6 io_wbs_data_o[7]
port 38 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 io_wbs_data_o[8]
port 39 nsew signal output
rlabel metal3 s 79200 25848 80000 25968 6 io_wbs_data_o[9]
port 40 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 io_wbs_m2s_addr[0]
port 41 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 io_wbs_m2s_addr[10]
port 42 nsew signal input
rlabel metal3 s 79200 43256 80000 43376 6 io_wbs_m2s_addr[11]
port 43 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 io_wbs_m2s_addr[12]
port 44 nsew signal input
rlabel metal2 s 41786 79200 41842 80000 6 io_wbs_m2s_addr[13]
port 45 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 io_wbs_m2s_addr[14]
port 46 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 io_wbs_m2s_addr[15]
port 47 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 io_wbs_m2s_addr[1]
port 48 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 io_wbs_m2s_addr[2]
port 49 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 io_wbs_m2s_addr[3]
port 50 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 io_wbs_m2s_addr[4]
port 51 nsew signal input
rlabel metal2 s 16302 79200 16358 80000 6 io_wbs_m2s_addr[5]
port 52 nsew signal input
rlabel metal2 s 23570 79200 23626 80000 6 io_wbs_m2s_addr[6]
port 53 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 io_wbs_m2s_addr[7]
port 54 nsew signal input
rlabel metal2 s 30838 79200 30894 80000 6 io_wbs_m2s_addr[8]
port 55 nsew signal input
rlabel metal3 s 79200 29384 80000 29504 6 io_wbs_m2s_addr[9]
port 56 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 io_wbs_m2s_data[0]
port 57 nsew signal input
rlabel metal3 s 79200 36320 80000 36440 6 io_wbs_m2s_data[10]
port 58 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 io_wbs_m2s_data[11]
port 59 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 io_wbs_m2s_data[12]
port 60 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 io_wbs_m2s_data[13]
port 61 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 io_wbs_m2s_data[14]
port 62 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 io_wbs_m2s_data[15]
port 63 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 io_wbs_m2s_data[16]
port 64 nsew signal input
rlabel metal2 s 49054 79200 49110 80000 6 io_wbs_m2s_data[17]
port 65 nsew signal input
rlabel metal3 s 79200 50192 80000 50312 6 io_wbs_m2s_data[18]
port 66 nsew signal input
rlabel metal2 s 56322 79200 56378 80000 6 io_wbs_m2s_data[19]
port 67 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 io_wbs_m2s_data[1]
port 68 nsew signal input
rlabel metal3 s 79200 57264 80000 57384 6 io_wbs_m2s_data[20]
port 69 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 io_wbs_m2s_data[21]
port 70 nsew signal input
rlabel metal2 s 63590 79200 63646 80000 6 io_wbs_m2s_data[22]
port 71 nsew signal input
rlabel metal3 s 79200 60664 80000 60784 6 io_wbs_m2s_data[23]
port 72 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 io_wbs_m2s_data[24]
port 73 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 io_wbs_m2s_data[25]
port 74 nsew signal input
rlabel metal2 s 70858 79200 70914 80000 6 io_wbs_m2s_data[26]
port 75 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 io_wbs_m2s_data[27]
port 76 nsew signal input
rlabel metal3 s 79200 74536 80000 74656 6 io_wbs_m2s_data[28]
port 77 nsew signal input
rlabel metal2 s 74446 79200 74502 80000 6 io_wbs_m2s_data[29]
port 78 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 io_wbs_m2s_data[2]
port 79 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 io_wbs_m2s_data[30]
port 80 nsew signal input
rlabel metal3 s 79200 78072 80000 78192 6 io_wbs_m2s_data[31]
port 81 nsew signal input
rlabel metal3 s 0 32240 800 32360 6 io_wbs_m2s_data[3]
port 82 nsew signal input
rlabel metal3 s 79200 18912 80000 19032 6 io_wbs_m2s_data[4]
port 83 nsew signal input
rlabel metal2 s 19890 79200 19946 80000 6 io_wbs_m2s_data[5]
port 84 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 io_wbs_m2s_data[6]
port 85 nsew signal input
rlabel metal2 s 27158 79200 27214 80000 6 io_wbs_m2s_data[7]
port 86 nsew signal input
rlabel metal2 s 34426 79200 34482 80000 6 io_wbs_m2s_data[8]
port 87 nsew signal input
rlabel metal3 s 79200 32920 80000 33040 6 io_wbs_m2s_data[9]
port 88 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 io_wbs_m2s_sel[0]
port 89 nsew signal input
rlabel metal2 s 9034 79200 9090 80000 6 io_wbs_m2s_sel[1]
port 90 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 io_wbs_m2s_sel[2]
port 91 nsew signal input
rlabel metal3 s 79200 15512 80000 15632 6 io_wbs_m2s_sel[3]
port 92 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 io_wbs_m2s_stb
port 93 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 io_wbs_m2s_we
port 94 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 reset
port 95 nsew signal input
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 96 nsew power input
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 96 nsew power input
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 96 nsew power input
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 97 nsew ground input
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 97 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16498720
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/Motor_Top/runs/Motor_Top/results/finishing/Motor_Top.magic.gds
string GDS_START 1023248
<< end >>

