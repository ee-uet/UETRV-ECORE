VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Motor_Top
  CLASS BLOCK ;
  FOREIGN Motor_Top ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 550.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 546.000 30.730 550.000 ;
    END
  END clock
  PIN io_ba_match
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END io_ba_match
  PIN io_motor_gpio_pwm_high
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END io_motor_gpio_pwm_high
  PIN io_motor_gpio_pwm_high_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END io_motor_gpio_pwm_high_en
  PIN io_motor_gpio_pwm_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END io_motor_gpio_pwm_low
  PIN io_motor_gpio_pwm_low_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END io_motor_gpio_pwm_low_en
  PIN io_motor_gpio_qei_ch_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END io_motor_gpio_qei_ch_a
  PIN io_motor_gpio_qei_ch_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END io_motor_gpio_qei_ch_b
  PIN io_motor_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END io_motor_irq
  PIN io_wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 34.040 550.000 34.640 ;
    END
  END io_wbs_ack_o
  PIN io_wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 102.720 550.000 103.320 ;
    END
  END io_wbs_data_o[0]
  PIN io_wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END io_wbs_data_o[10]
  PIN io_wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END io_wbs_data_o[11]
  PIN io_wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 546.000 213.810 550.000 ;
    END
  END io_wbs_data_o[12]
  PIN io_wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END io_wbs_data_o[13]
  PIN io_wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 514.800 550.000 515.400 ;
    END
  END io_wbs_data_o[14]
  PIN io_wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 546.000 274.990 550.000 ;
    END
  END io_wbs_data_o[15]
  PIN io_wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END io_wbs_data_o[16]
  PIN io_wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END io_wbs_data_o[17]
  PIN io_wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END io_wbs_data_o[18]
  PIN io_wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 546.000 336.170 550.000 ;
    END
  END io_wbs_data_o[19]
  PIN io_wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 171.400 550.000 172.000 ;
    END
  END io_wbs_data_o[1]
  PIN io_wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END io_wbs_data_o[20]
  PIN io_wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 546.000 397.350 550.000 ;
    END
  END io_wbs_data_o[21]
  PIN io_wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END io_wbs_data_o[22]
  PIN io_wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END io_wbs_data_o[23]
  PIN io_wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END io_wbs_data_o[24]
  PIN io_wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END io_wbs_data_o[25]
  PIN io_wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END io_wbs_data_o[26]
  PIN io_wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 546.000 458.530 550.000 ;
    END
  END io_wbs_data_o[27]
  PIN io_wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END io_wbs_data_o[28]
  PIN io_wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END io_wbs_data_o[29]
  PIN io_wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END io_wbs_data_o[2]
  PIN io_wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 546.000 519.710 550.000 ;
    END
  END io_wbs_data_o[30]
  PIN io_wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END io_wbs_data_o[31]
  PIN io_wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 546.000 152.630 550.000 ;
    END
  END io_wbs_data_o[3]
  PIN io_wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 240.080 550.000 240.680 ;
    END
  END io_wbs_data_o[4]
  PIN io_wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 308.760 550.000 309.360 ;
    END
  END io_wbs_data_o[5]
  PIN io_wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END io_wbs_data_o[6]
  PIN io_wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END io_wbs_data_o[7]
  PIN io_wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 377.440 550.000 378.040 ;
    END
  END io_wbs_data_o[8]
  PIN io_wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 446.120 550.000 446.720 ;
    END
  END io_wbs_data_o[9]
  PIN io_wbs_m2s_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END io_wbs_m2s_addr[0]
  PIN io_wbs_m2s_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END io_wbs_m2s_addr[10]
  PIN io_wbs_m2s_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END io_wbs_m2s_addr[11]
  PIN io_wbs_m2s_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END io_wbs_m2s_addr[12]
  PIN io_wbs_m2s_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END io_wbs_m2s_addr[13]
  PIN io_wbs_m2s_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END io_wbs_m2s_addr[14]
  PIN io_wbs_m2s_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_wbs_m2s_addr[15]
  PIN io_wbs_m2s_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END io_wbs_m2s_addr[1]
  PIN io_wbs_m2s_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END io_wbs_m2s_addr[2]
  PIN io_wbs_m2s_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END io_wbs_m2s_addr[3]
  PIN io_wbs_m2s_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_wbs_m2s_addr[4]
  PIN io_wbs_m2s_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END io_wbs_m2s_addr[5]
  PIN io_wbs_m2s_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END io_wbs_m2s_addr[6]
  PIN io_wbs_m2s_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END io_wbs_m2s_addr[7]
  PIN io_wbs_m2s_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END io_wbs_m2s_addr[8]
  PIN io_wbs_m2s_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END io_wbs_m2s_addr[9]
  PIN io_wbs_m2s_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END io_wbs_m2s_data[0]
  PIN io_wbs_m2s_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END io_wbs_m2s_data[10]
  PIN io_wbs_m2s_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END io_wbs_m2s_data[11]
  PIN io_wbs_m2s_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END io_wbs_m2s_data[12]
  PIN io_wbs_m2s_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END io_wbs_m2s_data[13]
  PIN io_wbs_m2s_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END io_wbs_m2s_data[14]
  PIN io_wbs_m2s_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END io_wbs_m2s_data[15]
  PIN io_wbs_m2s_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END io_wbs_m2s_data[16]
  PIN io_wbs_m2s_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END io_wbs_m2s_data[17]
  PIN io_wbs_m2s_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END io_wbs_m2s_data[18]
  PIN io_wbs_m2s_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END io_wbs_m2s_data[19]
  PIN io_wbs_m2s_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END io_wbs_m2s_data[1]
  PIN io_wbs_m2s_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END io_wbs_m2s_data[20]
  PIN io_wbs_m2s_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END io_wbs_m2s_data[21]
  PIN io_wbs_m2s_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END io_wbs_m2s_data[22]
  PIN io_wbs_m2s_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END io_wbs_m2s_data[23]
  PIN io_wbs_m2s_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END io_wbs_m2s_data[24]
  PIN io_wbs_m2s_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END io_wbs_m2s_data[25]
  PIN io_wbs_m2s_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END io_wbs_m2s_data[26]
  PIN io_wbs_m2s_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END io_wbs_m2s_data[27]
  PIN io_wbs_m2s_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.160 4.000 414.760 ;
    END
  END io_wbs_m2s_data[28]
  PIN io_wbs_m2s_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 422.320 4.000 422.920 ;
    END
  END io_wbs_m2s_data[29]
  PIN io_wbs_m2s_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END io_wbs_m2s_data[2]
  PIN io_wbs_m2s_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END io_wbs_m2s_data[30]
  PIN io_wbs_m2s_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END io_wbs_m2s_data[31]
  PIN io_wbs_m2s_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_wbs_m2s_data[3]
  PIN io_wbs_m2s_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END io_wbs_m2s_data[4]
  PIN io_wbs_m2s_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END io_wbs_m2s_data[5]
  PIN io_wbs_m2s_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_wbs_m2s_data[6]
  PIN io_wbs_m2s_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END io_wbs_m2s_data[7]
  PIN io_wbs_m2s_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END io_wbs_m2s_data[8]
  PIN io_wbs_m2s_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END io_wbs_m2s_data[9]
  PIN io_wbs_m2s_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END io_wbs_m2s_sel[0]
  PIN io_wbs_m2s_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END io_wbs_m2s_sel[1]
  PIN io_wbs_m2s_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END io_wbs_m2s_sel[2]
  PIN io_wbs_m2s_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END io_wbs_m2s_sel[3]
  PIN io_wbs_m2s_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END io_wbs_m2s_stb
  PIN io_wbs_m2s_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END io_wbs_m2s_we
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 546.000 91.450 550.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 538.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 538.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 544.180 538.645 ;
      LAYER met1 ;
        RECT 5.520 9.900 544.180 538.800 ;
      LAYER met2 ;
        RECT 6.990 545.720 30.170 546.450 ;
        RECT 31.010 545.720 90.890 546.450 ;
        RECT 91.730 545.720 152.070 546.450 ;
        RECT 152.910 545.720 213.250 546.450 ;
        RECT 214.090 545.720 274.430 546.450 ;
        RECT 275.270 545.720 335.610 546.450 ;
        RECT 336.450 545.720 396.790 546.450 ;
        RECT 397.630 545.720 457.970 546.450 ;
        RECT 458.810 545.720 519.150 546.450 ;
        RECT 519.990 545.720 541.330 546.450 ;
        RECT 6.990 4.280 541.330 545.720 ;
        RECT 6.990 4.000 20.970 4.280 ;
        RECT 21.810 4.000 63.290 4.280 ;
        RECT 64.130 4.000 105.610 4.280 ;
        RECT 106.450 4.000 147.930 4.280 ;
        RECT 148.770 4.000 190.250 4.280 ;
        RECT 191.090 4.000 232.570 4.280 ;
        RECT 233.410 4.000 274.890 4.280 ;
        RECT 275.730 4.000 317.210 4.280 ;
        RECT 318.050 4.000 359.530 4.280 ;
        RECT 360.370 4.000 401.850 4.280 ;
        RECT 402.690 4.000 444.170 4.280 ;
        RECT 445.010 4.000 486.490 4.280 ;
        RECT 487.330 4.000 528.810 4.280 ;
        RECT 529.650 4.000 541.330 4.280 ;
      LAYER met3 ;
        RECT 4.400 545.000 546.000 545.865 ;
        RECT 4.000 538.240 546.000 545.000 ;
        RECT 4.400 536.840 546.000 538.240 ;
        RECT 4.000 530.080 546.000 536.840 ;
        RECT 4.400 528.680 546.000 530.080 ;
        RECT 4.000 521.920 546.000 528.680 ;
        RECT 4.400 520.520 546.000 521.920 ;
        RECT 4.000 515.800 546.000 520.520 ;
        RECT 4.000 514.400 545.600 515.800 ;
        RECT 4.000 513.760 546.000 514.400 ;
        RECT 4.400 512.360 546.000 513.760 ;
        RECT 4.000 505.600 546.000 512.360 ;
        RECT 4.400 504.200 546.000 505.600 ;
        RECT 4.000 497.440 546.000 504.200 ;
        RECT 4.400 496.040 546.000 497.440 ;
        RECT 4.000 489.280 546.000 496.040 ;
        RECT 4.400 487.880 546.000 489.280 ;
        RECT 4.000 481.120 546.000 487.880 ;
        RECT 4.400 479.720 546.000 481.120 ;
        RECT 4.000 472.960 546.000 479.720 ;
        RECT 4.400 471.560 546.000 472.960 ;
        RECT 4.000 464.800 546.000 471.560 ;
        RECT 4.400 463.400 546.000 464.800 ;
        RECT 4.000 456.640 546.000 463.400 ;
        RECT 4.400 455.240 546.000 456.640 ;
        RECT 4.000 448.480 546.000 455.240 ;
        RECT 4.400 447.120 546.000 448.480 ;
        RECT 4.400 447.080 545.600 447.120 ;
        RECT 4.000 445.720 545.600 447.080 ;
        RECT 4.000 439.640 546.000 445.720 ;
        RECT 4.400 438.240 546.000 439.640 ;
        RECT 4.000 431.480 546.000 438.240 ;
        RECT 4.400 430.080 546.000 431.480 ;
        RECT 4.000 423.320 546.000 430.080 ;
        RECT 4.400 421.920 546.000 423.320 ;
        RECT 4.000 415.160 546.000 421.920 ;
        RECT 4.400 413.760 546.000 415.160 ;
        RECT 4.000 407.000 546.000 413.760 ;
        RECT 4.400 405.600 546.000 407.000 ;
        RECT 4.000 398.840 546.000 405.600 ;
        RECT 4.400 397.440 546.000 398.840 ;
        RECT 4.000 390.680 546.000 397.440 ;
        RECT 4.400 389.280 546.000 390.680 ;
        RECT 4.000 382.520 546.000 389.280 ;
        RECT 4.400 381.120 546.000 382.520 ;
        RECT 4.000 378.440 546.000 381.120 ;
        RECT 4.000 377.040 545.600 378.440 ;
        RECT 4.000 374.360 546.000 377.040 ;
        RECT 4.400 372.960 546.000 374.360 ;
        RECT 4.000 366.200 546.000 372.960 ;
        RECT 4.400 364.800 546.000 366.200 ;
        RECT 4.000 358.040 546.000 364.800 ;
        RECT 4.400 356.640 546.000 358.040 ;
        RECT 4.000 349.880 546.000 356.640 ;
        RECT 4.400 348.480 546.000 349.880 ;
        RECT 4.000 341.720 546.000 348.480 ;
        RECT 4.400 340.320 546.000 341.720 ;
        RECT 4.000 332.880 546.000 340.320 ;
        RECT 4.400 331.480 546.000 332.880 ;
        RECT 4.000 324.720 546.000 331.480 ;
        RECT 4.400 323.320 546.000 324.720 ;
        RECT 4.000 316.560 546.000 323.320 ;
        RECT 4.400 315.160 546.000 316.560 ;
        RECT 4.000 309.760 546.000 315.160 ;
        RECT 4.000 308.400 545.600 309.760 ;
        RECT 4.400 308.360 545.600 308.400 ;
        RECT 4.400 307.000 546.000 308.360 ;
        RECT 4.000 300.240 546.000 307.000 ;
        RECT 4.400 298.840 546.000 300.240 ;
        RECT 4.000 292.080 546.000 298.840 ;
        RECT 4.400 290.680 546.000 292.080 ;
        RECT 4.000 283.920 546.000 290.680 ;
        RECT 4.400 282.520 546.000 283.920 ;
        RECT 4.000 275.760 546.000 282.520 ;
        RECT 4.400 274.360 546.000 275.760 ;
        RECT 4.000 267.600 546.000 274.360 ;
        RECT 4.400 266.200 546.000 267.600 ;
        RECT 4.000 259.440 546.000 266.200 ;
        RECT 4.400 258.040 546.000 259.440 ;
        RECT 4.000 251.280 546.000 258.040 ;
        RECT 4.400 249.880 546.000 251.280 ;
        RECT 4.000 243.120 546.000 249.880 ;
        RECT 4.400 241.720 546.000 243.120 ;
        RECT 4.000 241.080 546.000 241.720 ;
        RECT 4.000 239.680 545.600 241.080 ;
        RECT 4.000 234.960 546.000 239.680 ;
        RECT 4.400 233.560 546.000 234.960 ;
        RECT 4.000 226.800 546.000 233.560 ;
        RECT 4.400 225.400 546.000 226.800 ;
        RECT 4.000 217.960 546.000 225.400 ;
        RECT 4.400 216.560 546.000 217.960 ;
        RECT 4.000 209.800 546.000 216.560 ;
        RECT 4.400 208.400 546.000 209.800 ;
        RECT 4.000 201.640 546.000 208.400 ;
        RECT 4.400 200.240 546.000 201.640 ;
        RECT 4.000 193.480 546.000 200.240 ;
        RECT 4.400 192.080 546.000 193.480 ;
        RECT 4.000 185.320 546.000 192.080 ;
        RECT 4.400 183.920 546.000 185.320 ;
        RECT 4.000 177.160 546.000 183.920 ;
        RECT 4.400 175.760 546.000 177.160 ;
        RECT 4.000 172.400 546.000 175.760 ;
        RECT 4.000 171.000 545.600 172.400 ;
        RECT 4.000 169.000 546.000 171.000 ;
        RECT 4.400 167.600 546.000 169.000 ;
        RECT 4.000 160.840 546.000 167.600 ;
        RECT 4.400 159.440 546.000 160.840 ;
        RECT 4.000 152.680 546.000 159.440 ;
        RECT 4.400 151.280 546.000 152.680 ;
        RECT 4.000 144.520 546.000 151.280 ;
        RECT 4.400 143.120 546.000 144.520 ;
        RECT 4.000 136.360 546.000 143.120 ;
        RECT 4.400 134.960 546.000 136.360 ;
        RECT 4.000 128.200 546.000 134.960 ;
        RECT 4.400 126.800 546.000 128.200 ;
        RECT 4.000 120.040 546.000 126.800 ;
        RECT 4.400 118.640 546.000 120.040 ;
        RECT 4.000 111.200 546.000 118.640 ;
        RECT 4.400 109.800 546.000 111.200 ;
        RECT 4.000 103.720 546.000 109.800 ;
        RECT 4.000 103.040 545.600 103.720 ;
        RECT 4.400 102.320 545.600 103.040 ;
        RECT 4.400 101.640 546.000 102.320 ;
        RECT 4.000 94.880 546.000 101.640 ;
        RECT 4.400 93.480 546.000 94.880 ;
        RECT 4.000 86.720 546.000 93.480 ;
        RECT 4.400 85.320 546.000 86.720 ;
        RECT 4.000 78.560 546.000 85.320 ;
        RECT 4.400 77.160 546.000 78.560 ;
        RECT 4.000 70.400 546.000 77.160 ;
        RECT 4.400 69.000 546.000 70.400 ;
        RECT 4.000 62.240 546.000 69.000 ;
        RECT 4.400 60.840 546.000 62.240 ;
        RECT 4.000 54.080 546.000 60.840 ;
        RECT 4.400 52.680 546.000 54.080 ;
        RECT 4.000 45.920 546.000 52.680 ;
        RECT 4.400 44.520 546.000 45.920 ;
        RECT 4.000 37.760 546.000 44.520 ;
        RECT 4.400 36.360 546.000 37.760 ;
        RECT 4.000 35.040 546.000 36.360 ;
        RECT 4.000 33.640 545.600 35.040 ;
        RECT 4.000 29.600 546.000 33.640 ;
        RECT 4.400 28.200 546.000 29.600 ;
        RECT 4.000 21.440 546.000 28.200 ;
        RECT 4.400 20.040 546.000 21.440 ;
        RECT 4.000 13.280 546.000 20.040 ;
        RECT 4.400 11.880 546.000 13.280 ;
        RECT 4.000 5.120 546.000 11.880 ;
        RECT 4.400 4.255 546.000 5.120 ;
      LAYER met4 ;
        RECT 50.895 11.735 97.440 458.825 ;
        RECT 99.840 11.735 174.240 458.825 ;
        RECT 176.640 11.735 251.040 458.825 ;
        RECT 253.440 11.735 303.305 458.825 ;
  END
END Motor_Top
END LIBRARY

