* NGSPICE file created from UART.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

.subckt UART clock io_rxd io_txd io_uartInt io_uart_select io_wbs_ack_o io_wbs_data_o[0]
+ io_wbs_data_o[10] io_wbs_data_o[11] io_wbs_data_o[12] io_wbs_data_o[13] io_wbs_data_o[14]
+ io_wbs_data_o[15] io_wbs_data_o[16] io_wbs_data_o[17] io_wbs_data_o[18] io_wbs_data_o[19]
+ io_wbs_data_o[1] io_wbs_data_o[20] io_wbs_data_o[21] io_wbs_data_o[22] io_wbs_data_o[23]
+ io_wbs_data_o[24] io_wbs_data_o[25] io_wbs_data_o[26] io_wbs_data_o[27] io_wbs_data_o[28]
+ io_wbs_data_o[29] io_wbs_data_o[2] io_wbs_data_o[30] io_wbs_data_o[31] io_wbs_data_o[3]
+ io_wbs_data_o[4] io_wbs_data_o[5] io_wbs_data_o[6] io_wbs_data_o[7] io_wbs_data_o[8]
+ io_wbs_data_o[9] io_wbs_m2s_addr[0] io_wbs_m2s_addr[10] io_wbs_m2s_addr[11] io_wbs_m2s_addr[12]
+ io_wbs_m2s_addr[13] io_wbs_m2s_addr[14] io_wbs_m2s_addr[15] io_wbs_m2s_addr[1] io_wbs_m2s_addr[2]
+ io_wbs_m2s_addr[3] io_wbs_m2s_addr[4] io_wbs_m2s_addr[5] io_wbs_m2s_addr[6] io_wbs_m2s_addr[7]
+ io_wbs_m2s_addr[8] io_wbs_m2s_addr[9] io_wbs_m2s_data[0] io_wbs_m2s_data[10] io_wbs_m2s_data[11]
+ io_wbs_m2s_data[12] io_wbs_m2s_data[13] io_wbs_m2s_data[14] io_wbs_m2s_data[15]
+ io_wbs_m2s_data[16] io_wbs_m2s_data[17] io_wbs_m2s_data[18] io_wbs_m2s_data[19]
+ io_wbs_m2s_data[1] io_wbs_m2s_data[20] io_wbs_m2s_data[21] io_wbs_m2s_data[22] io_wbs_m2s_data[23]
+ io_wbs_m2s_data[24] io_wbs_m2s_data[25] io_wbs_m2s_data[26] io_wbs_m2s_data[27]
+ io_wbs_m2s_data[28] io_wbs_m2s_data[29] io_wbs_m2s_data[2] io_wbs_m2s_data[30] io_wbs_m2s_data[31]
+ io_wbs_m2s_data[3] io_wbs_m2s_data[4] io_wbs_m2s_data[5] io_wbs_m2s_data[6] io_wbs_m2s_data[7]
+ io_wbs_m2s_data[8] io_wbs_m2s_data[9] io_wbs_m2s_stb io_wbs_m2s_we reset vccd1 vssd1
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0985_ _1145_/Q vssd1 vssd1 vccd1 vccd1 _0999_/B sky130_fd_sc_hd__inv_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0770_ _1097_/Q _1098_/Q _0770_/S vssd1 vssd1 vccd1 vccd1 _0771_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0968_ _1142_/Q _1141_/Q _0971_/S vssd1 vssd1 vccd1 vccd1 _0969_/B sky130_fd_sc_hd__mux2_1
X_0899_ _1037_/C _1044_/B _0898_/Y vssd1 vssd1 vccd1 vccd1 _0914_/A sky130_fd_sc_hd__o21bai_2
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0822_ _0822_/A vssd1 vssd1 vccd1 vccd1 _0822_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0684_ input6/X input5/X vssd1 vssd1 vccd1 vccd1 _0708_/B sky130_fd_sc_hd__or2b_1
X_0753_ _0753_/A vssd1 vssd1 vccd1 vccd1 _1091_/D sky130_fd_sc_hd__clkbuf_1
X_1098_ _1106_/CLK _1098_/D vssd1 vssd1 vccd1 vccd1 _1098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0829__C1 _0584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1021_ _1152_/Q vssd1 vssd1 vccd1 vccd1 _1021_/Y sky130_fd_sc_hd__inv_2
X_0805_ _0798_/X _0803_/X _0804_/X vssd1 vssd1 vccd1 vccd1 _1109_/D sky130_fd_sc_hd__o21a_1
X_0667_ input12/X _0657_/X _0666_/X _0664_/X vssd1 vssd1 vccd1 vccd1 _1066_/D sky130_fd_sc_hd__o211a_1
X_0598_ input11/X _1049_/Q _0622_/S vssd1 vssd1 vccd1 vccd1 _0599_/B sky130_fd_sc_hd__mux2_1
X_0736_ input3/X input4/X input2/X vssd1 vssd1 vccd1 vccd1 _0856_/C sky130_fd_sc_hd__and3b_1
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input18_A io_wbs_m2s_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1004_ _1023_/A _0988_/X _0825_/Y _0822_/A vssd1 vssd1 vccd1 vccd1 _1004_/X sky130_fd_sc_hd__a31o_1
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0719_ input14/X _1083_/Q _0726_/S vssd1 vssd1 vccd1 vccd1 _0720_/B sky130_fd_sc_hd__mux2_1
X_1163__36 vssd1 vssd1 vccd1 vccd1 _1163__36/HI io_wbs_data_o[11] sky130_fd_sc_hd__conb_1
Xoutput31 _1124_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_clock clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _1156_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0984_ _0980_/X _0983_/Y _0887_/X vssd1 vssd1 vccd1 vccd1 _1144_/D sky130_fd_sc_hd__o21a_1
XFILLER_42_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0967_ _0967_/A vssd1 vssd1 vccd1 vccd1 _1140_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1042__A0 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0898_ _1107_/Q input1/X vssd1 vssd1 vccd1 vccd1 _0898_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__0608__A0 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0821_ _0821_/A _0821_/B _0821_/C vssd1 vssd1 vccd1 vccd1 _0821_/X sky130_fd_sc_hd__or3_1
X_0752_ _0752_/A _0752_/B vssd1 vssd1 vccd1 vccd1 _0753_/A sky130_fd_sc_hd__or2_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0683_ _0683_/A _0683_/B vssd1 vssd1 vccd1 vccd1 _1073_/D sky130_fd_sc_hd__nor2_1
X_1097_ _1106_/CLK _1097_/D vssd1 vssd1 vccd1 vccd1 _1097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1169__42 vssd1 vssd1 vccd1 vccd1 _1169__42/HI io_wbs_data_o[17] sky130_fd_sc_hd__conb_1
X_1020_ _1018_/Y _1019_/X _0887_/X vssd1 vssd1 vccd1 vccd1 _1151_/D sky130_fd_sc_hd__o21a_1
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0735_ _1088_/Q vssd1 vssd1 vccd1 vccd1 _0799_/B sky130_fd_sc_hd__clkbuf_2
X_0804_ _0887_/A vssd1 vssd1 vccd1 vccd1 _0804_/X sky130_fd_sc_hd__clkbuf_2
X_0666_ _1066_/Q _0672_/B vssd1 vssd1 vccd1 vccd1 _0666_/X sky130_fd_sc_hd__or2_1
X_0597_ _0619_/S vssd1 vssd1 vccd1 vccd1 _0622_/S sky130_fd_sc_hd__buf_2
X_1149_ _1149_/CLK _1149_/D vssd1 vssd1 vccd1 vccd1 _1149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1003_ _0997_/Y _0988_/X _1148_/Q vssd1 vssd1 vccd1 vccd1 _1003_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__0977__C1 _0922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0718_ _0718_/A vssd1 vssd1 vccd1 vccd1 _1082_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_11_0_clock clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _1117_/CLK sky130_fd_sc_hd__clkbuf_2
X_0649_ _0722_/A vssd1 vssd1 vccd1 vccd1 _0699_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput32 _1125_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0671__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0983_ _0981_/Y _1023_/B _1144_/Q vssd1 vssd1 vccd1 vccd1 _0983_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0897_ _1126_/Q vssd1 vssd1 vccd1 vccd1 _0902_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0966_ _0972_/A _0966_/B vssd1 vssd1 vccd1 vccd1 _0967_/A sky130_fd_sc_hd__and2_1
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0820_ _0820_/A _0820_/B vssd1 vssd1 vccd1 vccd1 _0821_/C sky130_fd_sc_hd__nor2_1
X_0751_ input14/X _1091_/Q _0765_/S vssd1 vssd1 vccd1 vccd1 _0752_/B sky130_fd_sc_hd__mux2_1
X_0682_ _0682_/A _0682_/B _0682_/C _0737_/A vssd1 vssd1 vccd1 vccd1 _0683_/B sky130_fd_sc_hd__or4_1
X_1096_ _1117_/CLK _1096_/D vssd1 vssd1 vccd1 vccd1 _1096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0949_ _0971_/S vssd1 vssd1 vccd1 vccd1 _0962_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0765__A0 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0734_ _0734_/A vssd1 vssd1 vccd1 vccd1 _1087_/D sky130_fd_sc_hd__clkbuf_1
X_0803_ _0820_/A _0801_/X _0808_/B vssd1 vssd1 vccd1 vccd1 _0803_/X sky130_fd_sc_hd__o21ba_1
X_0665_ input11/X _0657_/X _0663_/X _0664_/X vssd1 vssd1 vccd1 vccd1 _1065_/D sky130_fd_sc_hd__o211a_1
X_0596_ _0682_/A _0708_/A vssd1 vssd1 vccd1 vccd1 _0619_/S sky130_fd_sc_hd__or2_1
X_1148_ _1156_/CLK _1148_/D vssd1 vssd1 vccd1 vccd1 _1148_/Q sky130_fd_sc_hd__dfxtp_1
X_1079_ _1158_/CLK _1079_/D vssd1 vssd1 vccd1 vccd1 _1079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1002_ _1148_/Q _1147_/Q _1007_/A _0988_/A vssd1 vssd1 vccd1 vccd1 _1002_/X sky130_fd_sc_hd__or4b_1
XFILLER_19_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0729__A0 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0717_ _0720_/A _0717_/B vssd1 vssd1 vccd1 vccd1 _0718_/A sky130_fd_sc_hd__and2_1
X_0648_ _0648_/A vssd1 vssd1 vccd1 vccd1 _1063_/D sky130_fd_sc_hd__clkbuf_1
X_0579_ _0922_/A _0579_/B _0579_/C vssd1 vssd1 vccd1 vccd1 _0580_/A sky130_fd_sc_hd__and3_1
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput22 _1097_/Q vssd1 vssd1 vccd1 vccd1 io_txd sky130_fd_sc_hd__buf_2
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_clock clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 _1110_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0982_ _0988_/A vssd1 vssd1 vccd1 vccd1 _1023_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0896_ _0878_/B _0894_/X _0895_/X _0843_/X vssd1 vssd1 vccd1 vccd1 _1125_/D sky130_fd_sc_hd__o211a_1
X_0965_ _1141_/Q _1140_/Q _0971_/S vssd1 vssd1 vccd1 vccd1 _0966_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0681_ input18/X _0657_/A _0680_/X _0674_/X vssd1 vssd1 vccd1 vccd1 _1072_/D sky130_fd_sc_hd__o211a_1
X_0750_ _0750_/A vssd1 vssd1 vccd1 vccd1 _1090_/D sky130_fd_sc_hd__clkbuf_1
X_1095_ _1095_/CLK _1095_/D vssd1 vssd1 vccd1 vccd1 _1095_/Q sky130_fd_sc_hd__dfxtp_2
X_0948_ _1006_/B _0948_/B vssd1 vssd1 vccd1 vccd1 _0971_/S sky130_fd_sc_hd__nand2_2
X_0879_ _0877_/X _0878_/X _0804_/X vssd1 vssd1 vccd1 vccd1 _1121_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0802_ _1109_/Q _1108_/Q _0802_/C vssd1 vssd1 vccd1 vccd1 _0808_/B sky130_fd_sc_hd__or3_1
X_0733_ _0740_/A _0733_/B vssd1 vssd1 vccd1 vccd1 _0734_/A sky130_fd_sc_hd__and2_1
X_0664_ _0922_/A vssd1 vssd1 vccd1 vccd1 _0664_/X sky130_fd_sc_hd__clkbuf_2
X_0595_ _0686_/A _0682_/C _0737_/A vssd1 vssd1 vccd1 vccd1 _0708_/A sky130_fd_sc_hd__or3_1
X_1147_ _1156_/CLK _1147_/D vssd1 vssd1 vccd1 vccd1 _1147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1078_ _1158_/CLK _1078_/D vssd1 vssd1 vccd1 vccd1 _1078_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0692__A0 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _0998_/X _1000_/Y _0887_/X vssd1 vssd1 vccd1 vccd1 _1147_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0716_ input13/X _1082_/Q _0726_/S vssd1 vssd1 vccd1 vccd1 _0717_/B sky130_fd_sc_hd__mux2_1
X_0578_ _1045_/Q _0802_/C _0820_/A _1046_/Q vssd1 vssd1 vccd1 vccd1 _0579_/C sky130_fd_sc_hd__or4b_1
X_0647_ _0647_/A _0647_/B vssd1 vssd1 vccd1 vccd1 _0648_/A sky130_fd_sc_hd__and2_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_clock clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 _1141_/CLK sky130_fd_sc_hd__clkbuf_2
Xoutput23 _0525_/X vssd1 vssd1 vccd1 vccd1 io_uartInt sky130_fd_sc_hd__buf_2
XANTENNA_input16_A io_wbs_m2s_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input8_A io_wbs_m2s_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0685__C_N input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0981_ _1143_/Q vssd1 vssd1 vccd1 vccd1 _0981_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_clock clock vssd1 vssd1 vccd1 vccd1 clkbuf_0_clock/X sky130_fd_sc_hd__clkbuf_16
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0964_ _0964_/A vssd1 vssd1 vccd1 vccd1 _1139_/D sky130_fd_sc_hd__clkbuf_1
X_0895_ _1072_/Q _0895_/B vssd1 vssd1 vccd1 vccd1 _0895_/X sky130_fd_sc_hd__or2_1
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0680_ _1072_/Q _0680_/B vssd1 vssd1 vccd1 vccd1 _0680_/X sky130_fd_sc_hd__or2_1
XFILLER_13_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1094_ _1143_/CLK _1094_/D vssd1 vssd1 vccd1 vccd1 _1094_/Q sky130_fd_sc_hd__dfxtp_1
X_0947_ _1037_/A _0947_/B vssd1 vssd1 vccd1 vccd1 _0948_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0878_ _1068_/Q _0878_/B vssd1 vssd1 vccd1 vccd1 _0878_/X sky130_fd_sc_hd__and2_1
XFILLER_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0736__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0801_ _0807_/B _0801_/B vssd1 vssd1 vccd1 vccd1 _0801_/X sky130_fd_sc_hd__or2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0663_ _1065_/Q _0672_/B vssd1 vssd1 vccd1 vccd1 _0663_/X sky130_fd_sc_hd__or2_1
X_1175__48 vssd1 vssd1 vccd1 vccd1 _1175__48/HI io_wbs_data_o[23] sky130_fd_sc_hd__conb_1
X_0732_ input18/X _1087_/Q _0732_/S vssd1 vssd1 vccd1 vccd1 _0733_/B sky130_fd_sc_hd__mux2_1
X_0594_ _0686_/B vssd1 vssd1 vccd1 vccd1 _0737_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1146_ _1152_/CLK _1146_/D vssd1 vssd1 vccd1 vccd1 _1146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1077_ _1121_/CLK _1077_/D vssd1 vssd1 vccd1 vccd1 _1077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_1_0_clock clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 _1137_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1000_ _0999_/X _1023_/B _1147_/Q vssd1 vssd1 vccd1 vccd1 _1000_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0715_ _0715_/A vssd1 vssd1 vccd1 vccd1 _1081_/D sky130_fd_sc_hd__clkbuf_1
X_0577_ _1073_/Q _0821_/A _0770_/S _0566_/Y _1046_/Q vssd1 vssd1 vccd1 vccd1 _0579_/B
+ sky130_fd_sc_hd__a221o_1
X_0646_ _1063_/Q _1141_/Q _0646_/S vssd1 vssd1 vccd1 vccd1 _0647_/B sky130_fd_sc_hd__mux2_1
X_1129_ _1149_/CLK _1129_/D vssd1 vssd1 vccd1 vccd1 _1129_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0665__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput24 _1096_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0629_ _1058_/Q _1136_/Q _0629_/S vssd1 vssd1 vccd1 vccd1 _0630_/B sky130_fd_sc_hd__mux2_1
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0980_ _1044_/A _0801_/X _0987_/C _0999_/C vssd1 vssd1 vccd1 vccd1 _0980_/X sky130_fd_sc_hd__o211a_1
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0894_ _1095_/Q _0853_/X _0893_/X vssd1 vssd1 vccd1 vccd1 _0894_/X sky130_fd_sc_hd__o21a_1
X_0963_ _0972_/A _0963_/B vssd1 vssd1 vccd1 vccd1 _0964_/A sky130_fd_sc_hd__and2_1
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1093_ _1143_/CLK _1093_/D vssd1 vssd1 vccd1 vccd1 _1093_/Q sky130_fd_sc_hd__dfxtp_2
X_0946_ _0992_/A _1007_/B _0946_/C vssd1 vssd1 vccd1 vccd1 _1006_/B sky130_fd_sc_hd__nor3_2
XANTENNA__0759__B1 _0584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0877_ _1091_/Q _0853_/X _0859_/X _0876_/X vssd1 vssd1 vccd1 vccd1 _0877_/X sky130_fd_sc_hd__o211a_1
XANTENNA__0736__C input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0731_ _0731_/A vssd1 vssd1 vccd1 vccd1 _1086_/D sky130_fd_sc_hd__clkbuf_1
X_0800_ _0800_/A _1088_/Q vssd1 vssd1 vccd1 vccd1 _0801_/B sky130_fd_sc_hd__and2_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0662_ _0680_/B vssd1 vssd1 vccd1 vccd1 _0672_/B sky130_fd_sc_hd__clkbuf_1
X_0593_ _0850_/B _0593_/B vssd1 vssd1 vccd1 vccd1 _0686_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1145_ _1152_/CLK _1145_/D vssd1 vssd1 vccd1 vccd1 _1145_/Q sky130_fd_sc_hd__dfxtp_1
X_1076_ _1135_/CLK _1076_/D vssd1 vssd1 vccd1 vccd1 _1076_/Q sky130_fd_sc_hd__dfxtp_1
X_0929_ _1131_/Q _0934_/C _0929_/C vssd1 vssd1 vccd1 vccd1 _0929_/X sky130_fd_sc_hd__and3_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0840__C1 _0584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0645_ _0645_/A vssd1 vssd1 vccd1 vccd1 _1062_/D sky130_fd_sc_hd__clkbuf_1
X_0714_ _0720_/A _0714_/B vssd1 vssd1 vccd1 vccd1 _0715_/A sky130_fd_sc_hd__and2_1
X_0576_ _0802_/C vssd1 vssd1 vccd1 vccd1 _0821_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__0848__A _0960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1128_ _1159_/CLK _1128_/D vssd1 vssd1 vccd1 vccd1 _1128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1059_ _1137_/CLK _1059_/D vssd1 vssd1 vccd1 vccd1 _1059_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput25 _1118_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[0] sky130_fd_sc_hd__buf_2
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0850__B _0850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0628_ _0628_/A vssd1 vssd1 vccd1 vccd1 _1057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0559_ _0559_/A vssd1 vssd1 vccd1 vccd1 _1104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input21_A reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0951__A _0960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0861__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0962_ _1140_/Q _1139_/Q _0962_/S vssd1 vssd1 vccd1 vccd1 _0963_/B sky130_fd_sc_hd__mux2_1
X_0893_ _1079_/Q _0865_/A _0866_/A _1064_/Q _0867_/A vssd1 vssd1 vccd1 vccd1 _0893_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1092_ _1143_/CLK _1092_/D vssd1 vssd1 vccd1 vccd1 _1092_/Q sky130_fd_sc_hd__dfxtp_1
X_0945_ _0941_/C _0943_/Y _0944_/X _0922_/X vssd1 vssd1 vccd1 vccd1 _1134_/D sky130_fd_sc_hd__o211a_1
X_0876_ _1075_/Q _0865_/X _0866_/X _1060_/Q _0867_/X vssd1 vssd1 vccd1 vccd1 _0876_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0695__A0 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0730_ _0740_/A _0730_/B vssd1 vssd1 vccd1 vccd1 _0731_/A sky130_fd_sc_hd__and2_1
X_0661_ _0858_/A _0737_/A _0861_/B _0861_/C vssd1 vssd1 vccd1 vccd1 _0680_/B sky130_fd_sc_hd__and4bb_1
X_0592_ input4/X input3/X input2/X vssd1 vssd1 vccd1 vccd1 _0682_/C sky130_fd_sc_hd__nand3b_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1144_ _1152_/CLK _1144_/D vssd1 vssd1 vccd1 vccd1 _1144_/Q sky130_fd_sc_hd__dfxtp_1
X_1075_ _1135_/CLK _1075_/D vssd1 vssd1 vccd1 vccd1 _1075_/Q sky130_fd_sc_hd__dfxtp_1
X_1166__39 vssd1 vssd1 vccd1 vccd1 _1166__39/HI io_wbs_data_o[14] sky130_fd_sc_hd__conb_1
X_0928_ _0934_/C _0914_/A _0929_/C _1131_/Q vssd1 vssd1 vccd1 vccd1 _0931_/B sky130_fd_sc_hd__a31o_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0859_ _0895_/B vssd1 vssd1 vccd1 vccd1 _0859_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1180__53 vssd1 vssd1 vccd1 vccd1 _1180__53/HI io_wbs_data_o[28] sky130_fd_sc_hd__conb_1
XANTENNA__0954__A _0960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0713_ input12/X _1081_/Q _0726_/S vssd1 vssd1 vccd1 vccd1 _0714_/B sky130_fd_sc_hd__mux2_1
X_0644_ _0647_/A _0644_/B vssd1 vssd1 vccd1 vccd1 _0645_/A sky130_fd_sc_hd__and2_1
X_0575_ _0845_/A vssd1 vssd1 vccd1 vccd1 _0922_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1127_ _1159_/CLK _1127_/D vssd1 vssd1 vccd1 vccd1 _1127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1058_ _1137_/CLK _1058_/D vssd1 vssd1 vccd1 vccd1 _1058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput26 _1119_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0558_ _0557_/X _1105_/Q _0558_/S vssd1 vssd1 vccd1 vccd1 _0559_/A sky130_fd_sc_hd__mux2_1
X_0627_ _0630_/A _0627_/B vssd1 vssd1 vccd1 vccd1 _0628_/A sky130_fd_sc_hd__and2_1
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input14_A io_wbs_m2s_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1039__A0 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input6_A io_wbs_m2s_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0961_ _0961_/A vssd1 vssd1 vccd1 vccd1 _1138_/D sky130_fd_sc_hd__clkbuf_1
X_0892_ _0890_/X _0891_/X _0887_/X vssd1 vssd1 vccd1 vccd1 _1124_/D sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_3_4_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0957__A _0960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1091_ _1110_/CLK _1091_/D vssd1 vssd1 vccd1 vccd1 _1091_/Q sky130_fd_sc_hd__dfxtp_2
X_0944_ _1133_/Q _0914_/X _0934_/X _1134_/Q vssd1 vssd1 vccd1 vccd1 _0944_/X sky130_fd_sc_hd__a31o_1
X_0875_ _0878_/B _0873_/X _0874_/X _0843_/X vssd1 vssd1 vccd1 vccd1 _1120_/D sky130_fd_sc_hd__o211a_1
XANTENNA__0850__A_N _0593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0591_ input8/X input7/X _0591_/C input9/X vssd1 vssd1 vccd1 vccd1 _0686_/A sky130_fd_sc_hd__or4_2
X_0660_ input2/X input4/X vssd1 vssd1 vccd1 vccd1 _0861_/C sky130_fd_sc_hd__and2_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1143_ _1143_/CLK _1143_/D vssd1 vssd1 vccd1 vccd1 _1143_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0677__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1074_ _1135_/CLK _1074_/D vssd1 vssd1 vccd1 vccd1 _1074_/Q sky130_fd_sc_hd__dfxtp_1
X_0927_ _0908_/A _0925_/X _0926_/Y _0584_/A vssd1 vssd1 vccd1 vccd1 _1130_/D sky130_fd_sc_hd__a211oi_1
X_0789_ _0785_/Y _0832_/A _0758_/Y _1130_/Q _0788_/X vssd1 vssd1 vccd1 vccd1 _0789_/Y
+ sky130_fd_sc_hd__a221oi_1
X_0858_ _0858_/A _0858_/B _0858_/C _0861_/D vssd1 vssd1 vccd1 vccd1 _0895_/B sky130_fd_sc_hd__or4b_2
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0643_ _1062_/Q _1140_/Q _0646_/S vssd1 vssd1 vccd1 vccd1 _0644_/B sky130_fd_sc_hd__mux2_1
X_0712_ _0732_/S vssd1 vssd1 vccd1 vccd1 _0726_/S sky130_fd_sc_hd__clkbuf_2
X_0574_ _0566_/Y _0794_/B _0820_/A _0569_/X _0887_/A vssd1 vssd1 vccd1 vccd1 _1045_/D
+ sky130_fd_sc_hd__o311a_1
X_1126_ _1149_/CLK _1126_/D vssd1 vssd1 vccd1 vccd1 _1126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1057_ _1135_/CLK _1057_/D vssd1 vssd1 vccd1 vccd1 _1057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput27 _1120_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0557_ _1054_/Q _1104_/Q _0557_/S vssd1 vssd1 vccd1 vccd1 _0557_/X sky130_fd_sc_hd__mux2_1
X_0626_ _1057_/Q _1135_/Q _0629_/S vssd1 vssd1 vccd1 vccd1 _0627_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1109_ _1110_/CLK _1109_/D vssd1 vssd1 vccd1 vccd1 _1109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0713__A0 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0609_ _0752_/A _0609_/B vssd1 vssd1 vccd1 vccd1 _0610_/A sky130_fd_sc_hd__or2_1
XFILLER_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0960_ _0960_/A _0960_/B vssd1 vssd1 vccd1 vccd1 _0961_/A sky130_fd_sc_hd__and2_1
X_0891_ _1071_/Q _0891_/B vssd1 vssd1 vccd1 vccd1 _0891_/X sky130_fd_sc_hd__and2_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0591__C _0591_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1090_ _1143_/CLK _1090_/D vssd1 vssd1 vccd1 vccd1 _1090_/Q sky130_fd_sc_hd__dfxtp_1
X_0943_ _1031_/A _1134_/Q vssd1 vssd1 vccd1 vccd1 _0943_/Y sky130_fd_sc_hd__nor2_1
X_0874_ _1067_/Q _0895_/B vssd1 vssd1 vccd1 vccd1 _0874_/X sky130_fd_sc_hd__or2_1
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0590_ _0654_/A vssd1 vssd1 vccd1 vccd1 _0682_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1142_ _1142_/CLK _1142_/D vssd1 vssd1 vccd1 vccd1 _1142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1073_ _1110_/CLK _1073_/D vssd1 vssd1 vccd1 vccd1 _1073_/Q sky130_fd_sc_hd__dfxtp_1
X_0926_ _0914_/X _0929_/C _0934_/C vssd1 vssd1 vccd1 vccd1 _0926_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0857_ _1158_/Q _0865_/A _0866_/A _1057_/Q _0867_/A vssd1 vssd1 vccd1 vccd1 _0857_/X
+ sky130_fd_sc_hd__a221o_1
X_0788_ _1129_/Q _1092_/Q vssd1 vssd1 vccd1 vccd1 _0788_/X sky130_fd_sc_hd__xor2_1
XANTENNA__1011__C1 _0922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0711_ _0711_/A vssd1 vssd1 vccd1 vccd1 _1080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0573_ _0941_/A vssd1 vssd1 vccd1 vccd1 _0887_/A sky130_fd_sc_hd__buf_2
X_0642_ _0642_/A vssd1 vssd1 vccd1 vccd1 _1061_/D sky130_fd_sc_hd__clkbuf_1
X_1125_ _1156_/CLK _1125_/D vssd1 vssd1 vccd1 vccd1 _1125_/Q sky130_fd_sc_hd__dfxtp_1
X_1171__44 vssd1 vssd1 vccd1 vccd1 _1171__44/HI io_wbs_data_o[19] sky130_fd_sc_hd__conb_1
XFILLER_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1056_ _1105_/CLK _1056_/D vssd1 vssd1 vccd1 vccd1 _1056_/Q sky130_fd_sc_hd__dfxtp_1
X_0909_ _0913_/B _0908_/A _0908_/Y _0843_/X vssd1 vssd1 vccd1 vccd1 _1127_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput28 _1121_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0625_ _1159_/Q vssd1 vssd1 vccd1 vccd1 _0629_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__0736__A_N input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0556_ _0556_/A vssd1 vssd1 vccd1 vccd1 _1103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1039_ input12/X _0821_/A _1042_/S vssd1 vssd1 vccd1 vccd1 _1039_/X sky130_fd_sc_hd__mux2_1
X_1108_ _1110_/CLK _1108_/D vssd1 vssd1 vccd1 vccd1 _1108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0608_ input14/X _1052_/Q _0619_/S vssd1 vssd1 vccd1 vccd1 _0609_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0539_ _0539_/A vssd1 vssd1 vccd1 vccd1 _1098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0890_ _0832_/A _0853_/A _0895_/B _0889_/X vssd1 vssd1 vccd1 vccd1 _0890_/X sky130_fd_sc_hd__o211a_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0698__A0 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0622__A0 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0689__A0 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0942_ _0942_/A vssd1 vssd1 vccd1 vccd1 _1133_/D sky130_fd_sc_hd__clkbuf_1
X_0873_ _0807_/A _0853_/X _0872_/X vssd1 vssd1 vccd1 vccd1 _0873_/X sky130_fd_sc_hd__o21a_1
XANTENNA__0613__A0 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1177__50 vssd1 vssd1 vccd1 vccd1 _1177__50/HI io_wbs_data_o[25] sky130_fd_sc_hd__conb_1
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1072_ _1095_/CLK _1072_/D vssd1 vssd1 vccd1 vccd1 _1072_/Q sky130_fd_sc_hd__dfxtp_1
X_1141_ _1141_/CLK _1141_/D vssd1 vssd1 vccd1 vccd1 _1141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0925_ _0934_/C _0929_/C _1031_/A vssd1 vssd1 vccd1 vccd1 _0925_/X sky130_fd_sc_hd__a21o_1
X_0787_ _0785_/Y _1094_/Q _0758_/Y _1130_/Q _0786_/Y vssd1 vssd1 vccd1 vccd1 _0787_/X
+ sky130_fd_sc_hd__o221a_1
X_0856_ _0682_/A _0682_/B _0856_/C _0861_/D vssd1 vssd1 vccd1 vccd1 _0867_/A sky130_fd_sc_hd__and4bb_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0710_ _0752_/A _0710_/B vssd1 vssd1 vccd1 vccd1 _0711_/A sky130_fd_sc_hd__or2_1
X_0641_ _0647_/A _0641_/B vssd1 vssd1 vccd1 vccd1 _0642_/A sky130_fd_sc_hd__and2_1
X_0572_ _0845_/A vssd1 vssd1 vccd1 vccd1 _0941_/A sky130_fd_sc_hd__clkbuf_2
X_1124_ _1159_/CLK _1124_/D vssd1 vssd1 vccd1 vccd1 _1124_/Q sky130_fd_sc_hd__dfxtp_1
X_1055_ _1106_/CLK _1055_/D vssd1 vssd1 vccd1 vccd1 _1055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0908_ _0908_/A _0908_/B vssd1 vssd1 vccd1 vccd1 _0908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput29 _1122_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[4] sky130_fd_sc_hd__buf_2
X_0839_ _1115_/Q _0846_/C _0839_/C vssd1 vssd1 vccd1 vccd1 _0842_/B sky130_fd_sc_hd__or3_1
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0624_ _0624_/A vssd1 vssd1 vccd1 vccd1 _1056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0555_ _0554_/X _1104_/Q _0558_/S vssd1 vssd1 vccd1 vccd1 _0556_/A sky130_fd_sc_hd__mux2_1
X_1038_ _0948_/B _1027_/Y _1037_/X _1156_/Q vssd1 vssd1 vccd1 vccd1 _1156_/D sky130_fd_sc_hd__a2bb2o_1
X_1107_ _1149_/CLK _1107_/D vssd1 vssd1 vccd1 vccd1 _1107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0607_ _0607_/A vssd1 vssd1 vccd1 vccd1 _1051_/D sky130_fd_sc_hd__clkbuf_1
X_0538_ _0529_/X _1099_/Q _0564_/A vssd1 vssd1 vccd1 vccd1 _0539_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_clock clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _1152_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA_input12_A io_wbs_m2s_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A io_wbs_m2s_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0941_ _0941_/A _0941_/B _0941_/C vssd1 vssd1 vccd1 vccd1 _0942_/A sky130_fd_sc_hd__and3_1
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0872_ _1074_/Q _0865_/A _0866_/A _1059_/Q _0867_/A vssd1 vssd1 vccd1 vccd1 _0872_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1071_ _1095_/CLK _1071_/D vssd1 vssd1 vccd1 vccd1 _1071_/Q sky130_fd_sc_hd__dfxtp_1
X_1140_ _1142_/CLK _1140_/D vssd1 vssd1 vccd1 vccd1 _1140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0924_ _1130_/Q vssd1 vssd1 vccd1 vccd1 _0934_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0598__A0 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0786_ _1127_/Q _0807_/A vssd1 vssd1 vccd1 vccd1 _0786_/Y sky130_fd_sc_hd__xnor2_1
X_0855_ _0682_/A _0682_/B _0855_/C _0861_/D vssd1 vssd1 vccd1 vccd1 _0866_/A sky130_fd_sc_hd__and4bb_1
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0571_ _0611_/A vssd1 vssd1 vccd1 vccd1 _0845_/A sky130_fd_sc_hd__clkbuf_2
X_0640_ _1061_/Q _1139_/Q _0646_/S vssd1 vssd1 vccd1 vccd1 _0641_/B sky130_fd_sc_hd__mux2_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1123_ _1142_/CLK _1123_/D vssd1 vssd1 vccd1 vccd1 _1123_/Q sky130_fd_sc_hd__dfxtp_1
X_1054_ _1105_/CLK _1054_/D vssd1 vssd1 vccd1 vccd1 _1054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0907_ _0913_/B _0902_/A _0906_/Y vssd1 vssd1 vccd1 vccd1 _0908_/B sky130_fd_sc_hd__a21o_1
X_0769_ _0769_/A vssd1 vssd1 vccd1 vccd1 _1096_/D sky130_fd_sc_hd__clkbuf_1
X_0838_ _0846_/C _0839_/C _1115_/Q vssd1 vssd1 vccd1 vccd1 _0838_/Y sky130_fd_sc_hd__o21ai_1
X_1162__35 vssd1 vssd1 vccd1 vccd1 _1162__35/HI io_wbs_data_o[10] sky130_fd_sc_hd__conb_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0554_ _1053_/Q _1103_/Q _0557_/S vssd1 vssd1 vccd1 vccd1 _0554_/X sky130_fd_sc_hd__mux2_1
X_0623_ _0630_/A _0623_/B vssd1 vssd1 vccd1 vccd1 _0624_/A sky130_fd_sc_hd__and2_1
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1106_ _1106_/CLK _1106_/D vssd1 vssd1 vccd1 vccd1 _1106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1037_ _1037_/A _1155_/Q _1037_/C _1037_/D vssd1 vssd1 vccd1 vccd1 _1037_/X sky130_fd_sc_hd__or4_1
Xclkbuf_4_10_0_clock clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _1106_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__0716__A0 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0606_ _0887_/A _0606_/B vssd1 vssd1 vccd1 vccd1 _0607_/A sky130_fd_sc_hd__and2_1
X_0537_ _0569_/B vssd1 vssd1 vccd1 vccd1 _0564_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1041__C1 _0922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0940_ _0940_/A _0940_/B vssd1 vssd1 vccd1 vccd1 _0941_/C sky130_fd_sc_hd__nand2_1
X_0871_ _0869_/X _0870_/X _0804_/X vssd1 vssd1 vccd1 vccd1 _1119_/D sky130_fd_sc_hd__o21a_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1168__41 vssd1 vssd1 vccd1 vccd1 _1168__41/HI io_wbs_data_o[16] sky130_fd_sc_hd__conb_1
XFILLER_45_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1070_ _1095_/CLK _1070_/D vssd1 vssd1 vccd1 vccd1 _1070_/Q sky130_fd_sc_hd__dfxtp_1
X_0923_ _1129_/Q _0908_/A _0921_/Y _0922_/X vssd1 vssd1 vccd1 vccd1 _1129_/D sky130_fd_sc_hd__o211a_1
X_0854_ _0682_/B _0708_/B _0855_/C _0854_/D vssd1 vssd1 vccd1 vccd1 _0865_/A sky130_fd_sc_hd__and4bb_1
X_0785_ _1131_/Q vssd1 vssd1 vccd1 vccd1 _0785_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0570_ _0601_/A vssd1 vssd1 vccd1 vccd1 _0611_/A sky130_fd_sc_hd__inv_2
X_1122_ _1141_/CLK _1122_/D vssd1 vssd1 vccd1 vccd1 _1122_/Q sky130_fd_sc_hd__dfxtp_1
X_1053_ _1105_/CLK _1053_/D vssd1 vssd1 vccd1 vccd1 _1053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0906_ _0913_/B _0902_/A _1037_/A vssd1 vssd1 vccd1 vccd1 _0906_/Y sky130_fd_sc_hd__o21ai_1
X_0837_ _1095_/Q _1006_/C vssd1 vssd1 vccd1 vccd1 _0837_/X sky130_fd_sc_hd__xor2_1
X_0699_ _0699_/A _0699_/B vssd1 vssd1 vccd1 vccd1 _0700_/A sky130_fd_sc_hd__and2_1
X_0768_ _0850_/B _0922_/A vssd1 vssd1 vccd1 vccd1 _0769_/A sky130_fd_sc_hd__and2_1
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0553_ _0553_/A vssd1 vssd1 vccd1 vccd1 _1102_/D sky130_fd_sc_hd__clkbuf_1
X_0622_ input18/X _1056_/Q _0622_/S vssd1 vssd1 vccd1 vccd1 _0623_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1105_ _1105_/CLK _1105_/D vssd1 vssd1 vccd1 vccd1 _1105_/Q sky130_fd_sc_hd__dfxtp_1
X_1036_ _1155_/Q _1027_/Y _1035_/Y _1025_/Y vssd1 vssd1 vccd1 vccd1 _1155_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0605_ input13/X _1051_/Q _0622_/S vssd1 vssd1 vccd1 vccd1 _0606_/B sky130_fd_sc_hd__mux2_1
X_0536_ _0770_/S vssd1 vssd1 vccd1 vccd1 _0569_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_41_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1019_ _1152_/Q _1023_/C _0987_/C _1013_/A _1017_/Y vssd1 vssd1 vccd1 vccd1 _1019_/X
+ sky130_fd_sc_hd__o2111a_1
Xclkbuf_4_8_0_clock clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 _1105_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0616__A0 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0870_ _1066_/Q _0878_/B vssd1 vssd1 vccd1 vccd1 _0870_/X sky130_fd_sc_hd__and2_1
X_0999_ _0999_/A _0999_/B _0999_/C vssd1 vssd1 vccd1 vccd1 _0999_/X sky130_fd_sc_hd__and3_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1183__56 vssd1 vssd1 vccd1 vccd1 _1183__56/HI io_wbs_data_o[31] sky130_fd_sc_hd__conb_1
Xclkbuf_3_5_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0922_ _0922_/A vssd1 vssd1 vccd1 vccd1 _0922_/X sky130_fd_sc_hd__buf_2
X_0853_ _0853_/A vssd1 vssd1 vccd1 vccd1 _0853_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0784_ _0780_/X _0784_/B _0784_/C _0784_/D vssd1 vssd1 vccd1 vccd1 _0784_/X sky130_fd_sc_hd__and4b_1
Xinput1 io_rxd vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1121_ _1121_/CLK _1121_/D vssd1 vssd1 vccd1 vccd1 _1121_/Q sky130_fd_sc_hd__dfxtp_1
X_1052_ _1110_/CLK _1052_/D vssd1 vssd1 vccd1 vccd1 _1052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0905_ _1107_/Q vssd1 vssd1 vccd1 vccd1 _1037_/A sky130_fd_sc_hd__inv_2
X_0767_ _0767_/A vssd1 vssd1 vccd1 vccd1 _1095_/D sky130_fd_sc_hd__clkbuf_1
X_0836_ _0834_/X _0835_/Y _0822_/X vssd1 vssd1 vccd1 vccd1 _1114_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0698_ input16/X _1077_/Q _0702_/S vssd1 vssd1 vccd1 vccd1 _0699_/B sky130_fd_sc_hd__mux2_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0621_ _0621_/A vssd1 vssd1 vccd1 vccd1 _1055_/D sky130_fd_sc_hd__clkbuf_1
X_0552_ _0551_/X _1103_/Q _0558_/S vssd1 vssd1 vccd1 vccd1 _0553_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1035_ _1155_/Q _1037_/D vssd1 vssd1 vccd1 vccd1 _1035_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1104_ _1105_/CLK _1104_/D vssd1 vssd1 vccd1 vccd1 _1104_/Q sky130_fd_sc_hd__dfxtp_1
X_0819_ _0824_/A _0832_/D vssd1 vssd1 vccd1 vccd1 _0820_/B sky130_fd_sc_hd__xnor2_2
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_4_0_clock clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 _1142_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0604_ _0604_/A vssd1 vssd1 vccd1 vccd1 _1050_/D sky130_fd_sc_hd__clkbuf_1
X_0535_ _0802_/C _0833_/B vssd1 vssd1 vccd1 vccd1 _0770_/S sky130_fd_sc_hd__nor2_1
X_1018_ _1013_/A _1023_/B _1017_/Y vssd1 vssd1 vccd1 vccd1 _1018_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A io_wbs_m2s_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_0998_ _1044_/A _0820_/B _0987_/C _0997_/Y vssd1 vssd1 vccd1 vccd1 _0998_/X sky130_fd_sc_hd__o211a_1
XANTENNA_input2_A io_uart_select vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0921_ _1031_/A _0929_/C _0920_/Y _0914_/X vssd1 vssd1 vccd1 vccd1 _0921_/Y sky130_fd_sc_hd__o31ai_1
X_0783_ _1126_/Q _1089_/Q vssd1 vssd1 vccd1 vccd1 _0784_/D sky130_fd_sc_hd__xnor2_1
X_0852_ _0861_/B _0856_/C _0861_/D vssd1 vssd1 vccd1 vccd1 _0853_/A sky130_fd_sc_hd__nand3_1
XANTENNA__0755__A0 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput2 io_uart_select vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1120_ _1159_/CLK _1120_/D vssd1 vssd1 vccd1 vccd1 _1120_/Q sky130_fd_sc_hd__dfxtp_1
X_1051_ _1105_/CLK _1051_/D vssd1 vssd1 vccd1 vccd1 _1051_/Q sky130_fd_sc_hd__dfxtp_1
X_0904_ _1127_/Q vssd1 vssd1 vccd1 vccd1 _0913_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0766_ _0766_/A _0766_/B vssd1 vssd1 vccd1 vccd1 _0767_/A sky130_fd_sc_hd__and2_1
X_0835_ _0846_/C _0839_/C vssd1 vssd1 vccd1 vccd1 _0835_/Y sky130_fd_sc_hd__nand2_1
X_0697_ _0697_/A vssd1 vssd1 vccd1 vccd1 _1076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_clock clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 _1135_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__0719__A0 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0551_ _1052_/Q _1102_/Q _0557_/S vssd1 vssd1 vccd1 vccd1 _0551_/X sky130_fd_sc_hd__mux2_1
X_0620_ _0752_/A _0620_/B vssd1 vssd1 vccd1 vccd1 _0621_/A sky130_fd_sc_hd__or2_1
XFILLER_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1034_ _1037_/A _1044_/A _1037_/D _1033_/X vssd1 vssd1 vccd1 vccd1 _1154_/D sky130_fd_sc_hd__o31ai_1
X_1103_ _1105_/CLK _1103_/D vssd1 vssd1 vccd1 vccd1 _1103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0749_ _0766_/A _0749_/B vssd1 vssd1 vccd1 vccd1 _0750_/A sky130_fd_sc_hd__and2_1
X_0818_ _1112_/Q _0827_/D vssd1 vssd1 vccd1 vccd1 _0821_/B sky130_fd_sc_hd__or2_1
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0603_ _0752_/A _0603_/B vssd1 vssd1 vccd1 vccd1 _0604_/A sky130_fd_sc_hd__or2_1
X_0534_ _1112_/Q _0534_/B _0827_/D _0534_/D vssd1 vssd1 vccd1 vccd1 _0833_/B sky130_fd_sc_hd__or4_2
XFILLER_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1017_ _1151_/Q vssd1 vssd1 vccd1 vccd1 _1017_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0997_ _1147_/Q _1007_/A vssd1 vssd1 vccd1 vccd1 _0997_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0920_ _1129_/Q _0920_/B vssd1 vssd1 vccd1 vccd1 _0920_/Y sky130_fd_sc_hd__nor2_1
X_0782_ _1128_/Q _1091_/Q vssd1 vssd1 vccd1 vccd1 _0784_/C sky130_fd_sc_hd__xnor2_1
X_0851_ _0854_/D vssd1 vssd1 vccd1 vccd1 _0861_/D sky130_fd_sc_hd__clkbuf_1
X_1174__47 vssd1 vssd1 vccd1 vccd1 _1174__47/HI io_wbs_data_o[22] sky130_fd_sc_hd__conb_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 io_wbs_m2s_addr[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1050_ _1105_/CLK _1050_/D vssd1 vssd1 vccd1 vccd1 _1050_/Q sky130_fd_sc_hd__dfxtp_1
X_0903_ _0902_/A _0898_/Y _0902_/Y _0843_/X vssd1 vssd1 vccd1 vccd1 _1126_/D sky130_fd_sc_hd__o211a_1
XFILLER_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0834_ _0846_/C _0839_/C _0833_/X vssd1 vssd1 vccd1 vccd1 _0834_/X sky130_fd_sc_hd__or3b_1
X_0765_ input18/X _1095_/Q _0765_/S vssd1 vssd1 vccd1 vccd1 _0766_/B sky130_fd_sc_hd__mux2_1
X_0696_ _0699_/A _0696_/B vssd1 vssd1 vccd1 vccd1 _0697_/A sky130_fd_sc_hd__and2_1
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0550_ _0550_/A vssd1 vssd1 vccd1 vccd1 _1101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1102_ _1105_/CLK _1102_/D vssd1 vssd1 vccd1 vccd1 _1102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1033_ _0987_/C _1027_/B _1031_/Y _1032_/Y vssd1 vssd1 vccd1 vccd1 _1033_/X sky130_fd_sc_hd__a31o_1
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0817_ _0794_/B _0827_/D _1112_/Q vssd1 vssd1 vccd1 vccd1 _0817_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0679_ input17/X _0657_/A _0678_/X _0674_/X vssd1 vssd1 vccd1 vccd1 _1071_/D sky130_fd_sc_hd__o211a_1
X_0748_ input13/X _0807_/A _0748_/S vssd1 vssd1 vccd1 vccd1 _0749_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0602_ input12/X _1050_/Q _0619_/S vssd1 vssd1 vccd1 vccd1 _0603_/B sky130_fd_sc_hd__mux2_1
X_0533_ _1115_/Q _1114_/Q _1113_/Q vssd1 vssd1 vccd1 vccd1 _0534_/D sky130_fd_sc_hd__or3_1
XANTENNA__0619__A0 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1016_ _1013_/Y _1014_/X _1015_/X vssd1 vssd1 vccd1 vccd1 _1150_/D sky130_fd_sc_hd__a21oi_1
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0996_ _0993_/X _0995_/X _0822_/X vssd1 vssd1 vccd1 vccd1 _1146_/D sky130_fd_sc_hd__a21oi_1
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0850_ _0593_/B _0850_/B vssd1 vssd1 vccd1 vccd1 _0854_/D sky130_fd_sc_hd__and2b_1
X_0781_ _1132_/Q _1095_/Q vssd1 vssd1 vccd1 vccd1 _0784_/B sky130_fd_sc_hd__xnor2_1
Xinput4 io_wbs_m2s_addr[1] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0979_ _1144_/Q _1143_/Q vssd1 vssd1 vccd1 vccd1 _0999_/C sky130_fd_sc_hd__nor2_1
XANTENNA__0903__C1 _0843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0902_ _0902_/A _0908_/A vssd1 vssd1 vccd1 vccd1 _0902_/Y sky130_fd_sc_hd__nand2_1
X_0833_ _0833_/A _0833_/B _1006_/C vssd1 vssd1 vccd1 vccd1 _0833_/X sky130_fd_sc_hd__or3b_1
X_0764_ _0764_/A vssd1 vssd1 vccd1 vccd1 _1094_/D sky130_fd_sc_hd__clkbuf_1
X_0695_ input15/X _1076_/Q _0702_/S vssd1 vssd1 vccd1 vccd1 _0696_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1032_ _1154_/Q vssd1 vssd1 vccd1 vccd1 _1032_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1101_ _1106_/CLK _1101_/D vssd1 vssd1 vccd1 vccd1 _1101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0747_ _1090_/Q vssd1 vssd1 vccd1 vccd1 _0807_/A sky130_fd_sc_hd__clkbuf_2
X_0816_ _0811_/Y _0815_/X _0683_/A vssd1 vssd1 vccd1 vccd1 _1111_/D sky130_fd_sc_hd__a21oi_1
X_0678_ _1071_/Q _0680_/B vssd1 vssd1 vccd1 vccd1 _0678_/X sky130_fd_sc_hd__or2_1
XFILLER_29_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_3_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0601_ _0601_/A vssd1 vssd1 vccd1 vccd1 _0752_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0660__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0532_ _1111_/Q _1110_/Q _1109_/Q _1108_/Q vssd1 vssd1 vccd1 vccd1 _0827_/D sky130_fd_sc_hd__or4_1
X_1015_ _1023_/A _0988_/X _0837_/X _0822_/A vssd1 vssd1 vccd1 vccd1 _1015_/X sky130_fd_sc_hd__a31o_1
XFILLER_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0655__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0995_ _0999_/B _0999_/C _1027_/A _0999_/A vssd1 vssd1 vccd1 vccd1 _0995_/X sky130_fd_sc_hd__a31o_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0780_ input1/X _1134_/Q _1133_/Q vssd1 vssd1 vccd1 vccd1 _0780_/X sky130_fd_sc_hd__or3_1
Xinput5 io_wbs_m2s_addr[2] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0978_ _0988_/A vssd1 vssd1 vccd1 vccd1 _0987_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1165__38 vssd1 vssd1 vccd1 vccd1 _1165__38/HI io_wbs_data_o[13] sky130_fd_sc_hd__conb_1
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0901_ _0940_/A vssd1 vssd1 vccd1 vccd1 _0908_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0763_ _0766_/A _0763_/B vssd1 vssd1 vccd1 vccd1 _0764_/A sky130_fd_sc_hd__and2_1
X_0832_ _0832_/A _1093_/Q _1092_/Q _0832_/D vssd1 vssd1 vccd1 vccd1 _1006_/C sky130_fd_sc_hd__or4_2
X_0694_ _0694_/A vssd1 vssd1 vccd1 vccd1 _1075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1031_ _1031_/A _1153_/Q vssd1 vssd1 vccd1 vccd1 _1031_/Y sky130_fd_sc_hd__nand2_1
X_1100_ _1106_/CLK _1100_/D vssd1 vssd1 vccd1 vccd1 _1100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0746_ _0746_/A vssd1 vssd1 vccd1 vccd1 _1089_/D sky130_fd_sc_hd__clkbuf_1
X_0815_ _0795_/Y _0991_/B _0811_/B _1111_/Q vssd1 vssd1 vccd1 vccd1 _0815_/X sky130_fd_sc_hd__a211o_1
X_0677_ input16/X _0657_/A _0676_/X _0674_/X vssd1 vssd1 vccd1 vccd1 _1070_/D sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_3_7_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input19_A io_wbs_m2s_stb vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0660__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0600_ _0600_/A vssd1 vssd1 vccd1 vccd1 _1049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0531_ _1117_/Q _1116_/Q vssd1 vssd1 vccd1 vccd1 _0534_/B sky130_fd_sc_hd__or2_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1014_ _1012_/B _0988_/X _1150_/Q vssd1 vssd1 vccd1 vccd1 _1014_/X sky130_fd_sc_hd__a21bo_1
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0729_ input17/X _1086_/Q _0732_/S vssd1 vssd1 vccd1 vccd1 _0730_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0655__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0994_ _1146_/Q vssd1 vssd1 vccd1 vccd1 _0999_/A sky130_fd_sc_hd__inv_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput6 io_wbs_m2s_addr[3] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0977_ _1143_/Q _0976_/A _0976_/Y _0922_/X vssd1 vssd1 vccd1 vccd1 _1143_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0900_ _0914_/A vssd1 vssd1 vccd1 vccd1 _0940_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0762_ input17/X _0832_/A _0765_/S vssd1 vssd1 vccd1 vccd1 _0763_/B sky130_fd_sc_hd__mux2_1
X_0831_ _1093_/Q _0824_/A _0832_/D _0832_/A vssd1 vssd1 vccd1 vccd1 _0833_/A sky130_fd_sc_hd__o31a_1
X_0693_ _0699_/A _0693_/B vssd1 vssd1 vccd1 vccd1 _0694_/A sky130_fd_sc_hd__and2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1030_ _1153_/Q _1154_/Q vssd1 vssd1 vccd1 vccd1 _1037_/D sky130_fd_sc_hd__or2_1
Xinput20 io_wbs_m2s_we vssd1 vssd1 vccd1 vccd1 _0593_/B sky130_fd_sc_hd__clkbuf_2
X_0814_ _0832_/D _0814_/B vssd1 vssd1 vccd1 vccd1 _0991_/B sky130_fd_sc_hd__and2_1
X_0676_ _1070_/Q _0680_/B vssd1 vssd1 vccd1 vccd1 _0676_/X sky130_fd_sc_hd__or2_1
X_0745_ _0766_/A _0745_/B vssd1 vssd1 vccd1 vccd1 _0746_/A sky130_fd_sc_hd__and2_1
X_1159_ _1159_/CLK _1159_/D vssd1 vssd1 vccd1 vccd1 _1159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0584__A _0584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0530_ _0827_/C vssd1 vssd1 vccd1 vccd1 _0802_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1013_ _1013_/A _1023_/B vssd1 vssd1 vccd1 vccd1 _1013_/Y sky130_fd_sc_hd__nand2_1
X_0728_ _0728_/A vssd1 vssd1 vccd1 vccd1 _1085_/D sky130_fd_sc_hd__clkbuf_1
X_0659_ _0682_/A _0682_/B vssd1 vssd1 vccd1 vccd1 _0861_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0993_ _0993_/A _1007_/A _1027_/A vssd1 vssd1 vccd1 vccd1 _0993_/X sky130_fd_sc_hd__or3b_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 io_wbs_m2s_addr[4] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
X_0976_ _0976_/A _0976_/B vssd1 vssd1 vccd1 vccd1 _0976_/Y sky130_fd_sc_hd__nand2_1
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0667__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0830_ _1114_/Q vssd1 vssd1 vccd1 vccd1 _0846_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__0960__A _0960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0761_ _1094_/Q vssd1 vssd1 vccd1 vccd1 _0832_/A sky130_fd_sc_hd__clkbuf_2
X_0692_ input14/X _1075_/Q _0702_/S vssd1 vssd1 vccd1 vccd1 _0693_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1170__43 vssd1 vssd1 vccd1 vccd1 _1170__43/HI io_wbs_data_o[18] sky130_fd_sc_hd__conb_1
XFILLER_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0959_ _1139_/Q _1138_/Q _0962_/S vssd1 vssd1 vccd1 vccd1 _0960_/B sky130_fd_sc_hd__mux2_1
XFILLER_46_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0780__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput10 io_wbs_m2s_addr[7] vssd1 vssd1 vccd1 vccd1 _0591_/C sky130_fd_sc_hd__buf_2
X_0813_ _0807_/A _0800_/A _1088_/Q _1091_/Q vssd1 vssd1 vccd1 vccd1 _0814_/B sky130_fd_sc_hd__o31ai_1
Xinput21 reset vssd1 vssd1 vccd1 vccd1 _0601_/A sky130_fd_sc_hd__clkbuf_2
X_0744_ input12/X _0800_/A _0748_/S vssd1 vssd1 vccd1 vccd1 _0745_/B sky130_fd_sc_hd__mux2_1
X_0675_ input15/X _0657_/X _0672_/X _0674_/X vssd1 vssd1 vccd1 vccd1 _1069_/D sky130_fd_sc_hd__o211a_1
XFILLER_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1158_ _1158_/CLK _1158_/D vssd1 vssd1 vccd1 vccd1 _1158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1089_ _1143_/CLK _1089_/D vssd1 vssd1 vccd1 vccd1 _1089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1012_ _1150_/Q _1012_/B vssd1 vssd1 vccd1 vccd1 _1013_/A sky130_fd_sc_hd__and2b_1
XANTENNA__0685__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0727_ _0740_/A _0727_/B vssd1 vssd1 vccd1 vccd1 _0728_/A sky130_fd_sc_hd__and2_1
X_0589_ input6/X input5/X vssd1 vssd1 vccd1 vccd1 _0654_/A sky130_fd_sc_hd__or2_1
X_0658_ _0686_/A vssd1 vssd1 vccd1 vccd1 _0682_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _1149_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0992_ _0992_/A vssd1 vssd1 vccd1 vccd1 _1007_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0592__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 io_wbs_m2s_addr[5] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ _0799_/B _1023_/A _1143_/Q vssd1 vssd1 vccd1 vccd1 _0976_/B sky130_fd_sc_hd__a21o_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0760_ input16/X _0748_/S _0759_/Y vssd1 vssd1 vccd1 vccd1 _1093_/D sky130_fd_sc_hd__o21a_1
X_0691_ _0691_/A vssd1 vssd1 vccd1 vccd1 _1074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0958_ _0958_/A vssd1 vssd1 vccd1 vccd1 _1137_/D sky130_fd_sc_hd__clkbuf_1
X_0889_ _1078_/Q _0865_/X _0866_/X _1063_/Q _0867_/X vssd1 vssd1 vccd1 vccd1 _0889_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0812_ _1091_/Q _1090_/Q _1089_/Q _1088_/Q vssd1 vssd1 vccd1 vccd1 _0832_/D sky130_fd_sc_hd__or4_2
X_0743_ _1089_/Q vssd1 vssd1 vccd1 vccd1 _0800_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 io_wbs_m2s_data[0] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_2
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0674_ _0972_/A vssd1 vssd1 vccd1 vccd1 _0674_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1157_ _1158_/CLK _1157_/D vssd1 vssd1 vccd1 vccd1 _1157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1088_ _1143_/CLK _1088_/D vssd1 vssd1 vccd1 vccd1 _1088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1011_ _1149_/Q _0976_/A _1010_/Y _0922_/X vssd1 vssd1 vccd1 vccd1 _1149_/D sky130_fd_sc_hd__o211a_1
XANTENNA__0685__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0726_ input16/X _1085_/Q _0726_/S vssd1 vssd1 vccd1 vccd1 _0727_/B sky130_fd_sc_hd__mux2_1
X_0657_ _0657_/A vssd1 vssd1 vccd1 vccd1 _0657_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0588_ _0563_/S _0585_/Y _0683_/A vssd1 vssd1 vccd1 vccd1 _1048_/D sky130_fd_sc_hd__a21oi_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input17_A io_wbs_m2s_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0709_ input11/X _1080_/Q _0732_/S vssd1 vssd1 vccd1 vccd1 _0710_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input9_A io_wbs_m2s_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0991_ _1006_/B _0991_/B vssd1 vssd1 vccd1 vccd1 _0993_/A sky130_fd_sc_hd__and2_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0592__C input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 io_wbs_m2s_addr[6] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0974_ _1006_/B vssd1 vssd1 vccd1 vccd1 _1023_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0690_ _0699_/A _0690_/B vssd1 vssd1 vccd1 vccd1 _0691_/A sky130_fd_sc_hd__and2_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0888_ _0885_/X _0886_/X _0887_/X vssd1 vssd1 vccd1 vccd1 _1123_/D sky130_fd_sc_hd__o21a_1
X_0957_ _0960_/A _0957_/B vssd1 vssd1 vccd1 vccd1 _0958_/A sky130_fd_sc_hd__and2_1
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1161__34 vssd1 vssd1 vccd1 vccd1 _1161__34/HI io_wbs_data_o[9] sky130_fd_sc_hd__conb_1
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput12 io_wbs_m2s_data[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_4
X_0742_ _0845_/A vssd1 vssd1 vccd1 vccd1 _0766_/A sky130_fd_sc_hd__clkbuf_1
X_0673_ _0845_/A vssd1 vssd1 vccd1 vccd1 _0972_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0811_ _1111_/Q _0811_/B vssd1 vssd1 vccd1 vccd1 _0811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1156_ _1156_/CLK _1156_/D vssd1 vssd1 vccd1 vccd1 _1156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1087_ _1121_/CLK _1087_/D vssd1 vssd1 vccd1 vccd1 _1087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1010_ _1006_/X _1009_/Y _0976_/A vssd1 vssd1 vccd1 vccd1 _1010_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0945__C1 _0922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0725_ _0725_/A vssd1 vssd1 vccd1 vccd1 _1084_/D sky130_fd_sc_hd__clkbuf_1
X_0656_ _0858_/A _0737_/A _0858_/B _0858_/C vssd1 vssd1 vccd1 vccd1 _0657_/A sky130_fd_sc_hd__or4_2
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0587_ _0822_/A vssd1 vssd1 vccd1 vccd1 _0683_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1139_ _1141_/CLK _1139_/D vssd1 vssd1 vccd1 vccd1 _1139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0927__C1 _0584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0708_ _0708_/A _0708_/B vssd1 vssd1 vccd1 vccd1 _0732_/S sky130_fd_sc_hd__or2_2
X_0639_ _0639_/A vssd1 vssd1 vccd1 vccd1 _1060_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_7_0_clock clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 _1159_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__0909__C1 _0843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0990_ _0987_/Y _0989_/X _0822_/X vssd1 vssd1 vccd1 vccd1 _1145_/D sky130_fd_sc_hd__a21oi_1
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0679__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1167__40 vssd1 vssd1 vccd1 vccd1 _1167__40/HI io_wbs_data_o[15] sky130_fd_sc_hd__conb_1
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0973_ _0973_/A vssd1 vssd1 vccd1 vccd1 _1142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__0751__A0 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0956_ _1138_/Q _1137_/Q _0962_/S vssd1 vssd1 vccd1 vccd1 _0957_/B sky130_fd_sc_hd__mux2_1
X_0887_ _0887_/A vssd1 vssd1 vccd1 vccd1 _0887_/X sky130_fd_sc_hd__buf_2
XFILLER_46_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput13 io_wbs_m2s_data[2] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_4
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0810_ _0806_/Y _0809_/X _0683_/A vssd1 vssd1 vccd1 vccd1 _1110_/D sky130_fd_sc_hd__a21oi_1
X_0672_ _1069_/Q _0672_/B vssd1 vssd1 vccd1 vccd1 _0672_/X sky130_fd_sc_hd__or2_1
X_0741_ _0741_/A vssd1 vssd1 vccd1 vccd1 _1088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1155_ _1156_/CLK _1155_/D vssd1 vssd1 vccd1 vccd1 _1155_/Q sky130_fd_sc_hd__dfxtp_1
X_1086_ _1121_/CLK _1086_/D vssd1 vssd1 vccd1 vccd1 _1086_/Q sky130_fd_sc_hd__dfxtp_1
X_0939_ _1133_/Q _0934_/X _1026_/A vssd1 vssd1 vccd1 vccd1 _0940_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0724_ _0740_/A _0724_/B vssd1 vssd1 vccd1 vccd1 _0725_/A sky130_fd_sc_hd__and2_1
X_0586_ _0601_/A vssd1 vssd1 vccd1 vccd1 _0822_/A sky130_fd_sc_hd__clkbuf_2
X_0655_ input2/X input4/X vssd1 vssd1 vccd1 vccd1 _0858_/C sky130_fd_sc_hd__nand2_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1069_ _1142_/CLK _1069_/D vssd1 vssd1 vccd1 vccd1 _1069_/Q sky130_fd_sc_hd__dfxtp_1
X_1138_ _1142_/CLK _1138_/D vssd1 vssd1 vccd1 vccd1 _1138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_clock clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 _1158_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0707_ _0707_/A vssd1 vssd1 vccd1 vccd1 _1079_/D sky130_fd_sc_hd__clkbuf_1
X_0569_ _1045_/Q _0569_/B _0563_/S vssd1 vssd1 vccd1 vccd1 _0569_/X sky130_fd_sc_hd__or3b_1
X_0638_ _0647_/A _0638_/B vssd1 vssd1 vccd1 vccd1 _0639_/A sky130_fd_sc_hd__and2_1
XFILLER_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1119__D _1119_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1182__55 vssd1 vssd1 vccd1 vccd1 _1182__55/HI io_wbs_data_o[30] sky130_fd_sc_hd__conb_1
Xclkbuf_3_0_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0972_ _0972_/A _0972_/B vssd1 vssd1 vccd1 vccd1 _0973_/A sky130_fd_sc_hd__and2_1
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0760__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0886_ _1070_/Q _0891_/B vssd1 vssd1 vccd1 vccd1 _0886_/X sky130_fd_sc_hd__and2_1
X_0955_ _0955_/A vssd1 vssd1 vccd1 vccd1 _1136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 io_wbs_m2s_data[3] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_2
X_0740_ _0740_/A _0740_/B vssd1 vssd1 vccd1 vccd1 _0741_/A sky130_fd_sc_hd__and2_1
X_0671_ input14/X _0657_/X _0670_/X _0664_/X vssd1 vssd1 vccd1 vccd1 _1068_/D sky130_fd_sc_hd__o211a_1
X_1154_ _1156_/CLK _1154_/D vssd1 vssd1 vccd1 vccd1 _1154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1085_ _1105_/CLK _1085_/D vssd1 vssd1 vccd1 vccd1 _1085_/Q sky130_fd_sc_hd__dfxtp_1
X_0938_ _0940_/A _0934_/X _1133_/Q vssd1 vssd1 vccd1 vccd1 _0941_/B sky130_fd_sc_hd__a21o_1
X_0869_ _0800_/A _0853_/X _0859_/X _0868_/X vssd1 vssd1 vccd1 vccd1 _0869_/X sky130_fd_sc_hd__o211a_1
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0723_ input15/X _1084_/Q _0726_/S vssd1 vssd1 vccd1 vccd1 _0724_/B sky130_fd_sc_hd__mux2_1
X_0654_ _0654_/A _0686_/A vssd1 vssd1 vccd1 vccd1 _0858_/B sky130_fd_sc_hd__or2_1
X_0585_ _1047_/Q _0583_/B _1048_/Q vssd1 vssd1 vccd1 vccd1 _0585_/Y sky130_fd_sc_hd__o21ai_1
X_1137_ _1137_/CLK _1137_/D vssd1 vssd1 vccd1 vccd1 _1137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1068_ _1141_/CLK _1068_/D vssd1 vssd1 vccd1 vccd1 _1068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0706_ _0720_/A _0706_/B vssd1 vssd1 vccd1 vccd1 _0707_/A sky130_fd_sc_hd__and2_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0568_ _0833_/B vssd1 vssd1 vccd1 vccd1 _0820_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0637_ _1060_/Q _1138_/Q _0646_/S vssd1 vssd1 vccd1 vccd1 _0638_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input15_A io_wbs_m2s_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0898__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A io_wbs_m2s_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ input1/X _1142_/Q _0971_/S vssd1 vssd1 vccd1 vccd1 _0972_/B sky130_fd_sc_hd__mux2_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0885_ _1093_/Q _0853_/A _0859_/X _0884_/X vssd1 vssd1 vccd1 vccd1 _0885_/X sky130_fd_sc_hd__o211a_1
X_0954_ _0960_/A _0954_/B vssd1 vssd1 vccd1 vccd1 _0955_/A sky130_fd_sc_hd__and2_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 io_wbs_m2s_data[4] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_2
X_0670_ _1068_/Q _0672_/B vssd1 vssd1 vccd1 vccd1 _0670_/X sky130_fd_sc_hd__or2_1
X_1153_ _1156_/CLK _1153_/D vssd1 vssd1 vccd1 vccd1 _1153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1084_ _1121_/CLK _1084_/D vssd1 vssd1 vccd1 vccd1 _1084_/Q sky130_fd_sc_hd__dfxtp_1
X_0937_ _0937_/A vssd1 vssd1 vccd1 vccd1 _1132_/D sky130_fd_sc_hd__clkbuf_1
X_0799_ _0800_/A _0799_/B vssd1 vssd1 vccd1 vccd1 _0807_/B sky130_fd_sc_hd__nor2_1
X_0868_ _1157_/Q _0865_/X _0866_/X _1058_/Q _0867_/X vssd1 vssd1 vccd1 vccd1 _0868_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0722_ _0722_/A vssd1 vssd1 vccd1 vccd1 _0740_/A sky130_fd_sc_hd__clkbuf_2
X_0653_ input3/X vssd1 vssd1 vccd1 vccd1 _0858_/A sky130_fd_sc_hd__inv_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0584_ _0584_/A _0794_/B _0584_/C vssd1 vssd1 vccd1 vccd1 _1047_/D sky130_fd_sc_hd__nor3_1
X_1067_ _1142_/CLK _1067_/D vssd1 vssd1 vccd1 vccd1 _1067_/Q sky130_fd_sc_hd__dfxtp_1
X_1136_ _1137_/CLK _1136_/D vssd1 vssd1 vccd1 vccd1 _1136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0705_ input18/X _1079_/Q _0705_/S vssd1 vssd1 vccd1 vccd1 _0706_/B sky130_fd_sc_hd__mux2_1
X_0636_ _0636_/A vssd1 vssd1 vccd1 vccd1 _1059_/D sky130_fd_sc_hd__clkbuf_1
X_0567_ _0802_/C vssd1 vssd1 vccd1 vccd1 _0794_/B sky130_fd_sc_hd__clkbuf_2
X_1119_ _1156_/CLK _1119_/D vssd1 vssd1 vccd1 vccd1 _1119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0619_ input17/X _1055_/Q _0619_/S vssd1 vssd1 vccd1 vccd1 _0620_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0970_ _0970_/A vssd1 vssd1 vccd1 vccd1 _1141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1173__46 vssd1 vssd1 vccd1 vccd1 _1173__46/HI io_wbs_data_o[21] sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_0_clock_A clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_2_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0953_ _1137_/Q _1136_/Q _0962_/S vssd1 vssd1 vccd1 vccd1 _0954_/B sky130_fd_sc_hd__mux2_1
X_0884_ _1077_/Q _0865_/X _0866_/X _1062_/Q _0867_/X vssd1 vssd1 vccd1 vccd1 _0884_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput16 io_wbs_m2s_data[5] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_4
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0709__A0 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1152_ _1152_/CLK _1152_/D vssd1 vssd1 vccd1 vccd1 _1152_/Q sky130_fd_sc_hd__dfxtp_1
X_1083_ _1121_/CLK _1083_/D vssd1 vssd1 vccd1 vccd1 _1083_/Q sky130_fd_sc_hd__dfxtp_1
X_0936_ _0941_/A _0936_/B _0936_/C vssd1 vssd1 vccd1 vccd1 _0937_/A sky130_fd_sc_hd__and3_1
X_0867_ _0867_/A vssd1 vssd1 vccd1 vccd1 _0867_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0798_ _1108_/Q _0794_/B _1109_/Q vssd1 vssd1 vccd1 vccd1 _0798_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0875__C1 _0843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0721_ _0721_/A vssd1 vssd1 vccd1 vccd1 _1083_/D sky130_fd_sc_hd__clkbuf_1
X_0583_ _1047_/Q _0583_/B vssd1 vssd1 vccd1 vccd1 _0584_/C sky130_fd_sc_hd__xor2_1
X_0652_ _0652_/A vssd1 vssd1 vccd1 vccd1 _1064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1066_ _1095_/CLK _1066_/D vssd1 vssd1 vccd1 vccd1 _1066_/Q sky130_fd_sc_hd__dfxtp_1
X_1135_ _1135_/CLK _1135_/D vssd1 vssd1 vccd1 vccd1 _1135_/Q sky130_fd_sc_hd__dfxtp_1
X_0919_ _0934_/D vssd1 vssd1 vccd1 vccd1 _0929_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0704_ _0704_/A vssd1 vssd1 vccd1 vccd1 _1078_/D sky130_fd_sc_hd__clkbuf_1
X_0566_ _1045_/Q vssd1 vssd1 vccd1 vccd1 _0566_/Y sky130_fd_sc_hd__inv_2
X_0635_ _0647_/A _0635_/B vssd1 vssd1 vccd1 vccd1 _0636_/A sky130_fd_sc_hd__and2_1
X_1118_ _1159_/CLK _1118_/D vssd1 vssd1 vccd1 vccd1 _1118_/Q sky130_fd_sc_hd__dfxtp_1
X_1049_ _1106_/CLK _1049_/D vssd1 vssd1 vccd1 vccd1 _1049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1179__52 vssd1 vssd1 vccd1 vccd1 _1179__52/HI io_wbs_data_o[27] sky130_fd_sc_hd__conb_1
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0549_ _0548_/X _1102_/Q _0558_/S vssd1 vssd1 vccd1 vccd1 _0550_/A sky130_fd_sc_hd__mux2_1
X_0618_ _0618_/A vssd1 vssd1 vccd1 vccd1 _1054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input20_A io_wbs_m2s_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_6_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0952_ _0952_/A vssd1 vssd1 vccd1 vccd1 _1135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0883_ _0881_/X _0882_/X _0804_/X vssd1 vssd1 vccd1 vccd1 _1122_/D sky130_fd_sc_hd__o21a_1
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 io_wbs_m2s_data[6] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1151_ _1152_/CLK _1151_/D vssd1 vssd1 vccd1 vccd1 _1151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1082_ _1121_/CLK _1082_/D vssd1 vssd1 vccd1 vccd1 _1082_/Q sky130_fd_sc_hd__dfxtp_1
X_0935_ _1026_/A _0934_/X _0940_/A vssd1 vssd1 vccd1 vccd1 _0936_/C sky130_fd_sc_hd__o21ai_1
X_0866_ _0866_/A vssd1 vssd1 vccd1 vccd1 _0866_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0797_ _0794_/Y _0796_/X _0683_/A vssd1 vssd1 vccd1 vccd1 _1108_/D sky130_fd_sc_hd__a21oi_1
XFILLER_22_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0720_ _0720_/A _0720_/B vssd1 vssd1 vccd1 vccd1 _0721_/A sky130_fd_sc_hd__and2_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0582_ _1045_/Q _1046_/Q _0833_/B vssd1 vssd1 vccd1 vccd1 _0583_/B sky130_fd_sc_hd__or3_1
X_0651_ _0699_/A _0651_/B vssd1 vssd1 vccd1 vccd1 _0652_/A sky130_fd_sc_hd__and2_1
X_1134_ _1156_/CLK _1134_/D vssd1 vssd1 vccd1 vccd1 _1134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1065_ _1141_/CLK _1065_/D vssd1 vssd1 vccd1 vccd1 _1065_/Q sky130_fd_sc_hd__dfxtp_1
X_0918_ _1129_/Q _1128_/Q _1127_/Q _1126_/Q vssd1 vssd1 vccd1 vccd1 _0934_/D sky130_fd_sc_hd__and4_1
X_0849_ _0849_/A vssd1 vssd1 vccd1 vccd1 _1117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0703_ _0720_/A _0703_/B vssd1 vssd1 vccd1 vccd1 _0704_/A sky130_fd_sc_hd__and2_1
X_0565_ _0565_/A vssd1 vssd1 vccd1 vccd1 _1106_/D sky130_fd_sc_hd__clkbuf_1
X_0634_ _1059_/Q _1137_/Q _0646_/S vssd1 vssd1 vccd1 vccd1 _0635_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1117_ _1117_/CLK _1117_/D vssd1 vssd1 vccd1 vccd1 _1117_/Q sky130_fd_sc_hd__dfxtp_1
X_1048_ _1117_/CLK _1048_/D vssd1 vssd1 vccd1 vccd1 _1048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0548_ _1051_/Q _1101_/Q _0557_/S vssd1 vssd1 vccd1 vccd1 _0548_/X sky130_fd_sc_hd__mux2_1
X_0617_ _0630_/A _0617_/B vssd1 vssd1 vccd1 vccd1 _0618_/A sky130_fd_sc_hd__and2_1
XFILLER_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input13_A io_wbs_m2s_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1164__37 vssd1 vssd1 vccd1 vccd1 _1164__37/HI io_wbs_data_o[12] sky130_fd_sc_hd__conb_1
XANTENNA_input5_A io_wbs_m2s_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0681__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0882_ _1069_/Q _0891_/B vssd1 vssd1 vccd1 vccd1 _0882_/X sky130_fd_sc_hd__and2_1
X_0951_ _0960_/A _0951_/B vssd1 vssd1 vccd1 vccd1 _0952_/A sky130_fd_sc_hd__and2_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 io_wbs_m2s_data[7] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_4
X_1150_ _1152_/CLK _1150_/D vssd1 vssd1 vccd1 vccd1 _1150_/Q sky130_fd_sc_hd__dfxtp_1
X_1081_ _1110_/CLK _1081_/D vssd1 vssd1 vccd1 vccd1 _1081_/Q sky130_fd_sc_hd__dfxtp_1
X_0934_ _1132_/Q _1131_/Q _0934_/C _0934_/D vssd1 vssd1 vccd1 vccd1 _0934_/X sky130_fd_sc_hd__and4_1
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0865_ _0865_/A vssd1 vssd1 vccd1 vccd1 _0865_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0796_ _0799_/B _0795_/Y _0821_/A _1108_/Q vssd1 vssd1 vccd1 vccd1 _0796_/X sky130_fd_sc_hd__a211o_1
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0650_ _1064_/Q _1142_/Q _1159_/Q vssd1 vssd1 vccd1 vccd1 _0651_/B sky130_fd_sc_hd__mux2_1
X_0581_ _0601_/A vssd1 vssd1 vccd1 vccd1 _0584_/A sky130_fd_sc_hd__buf_2
X_1133_ _1156_/CLK _1133_/D vssd1 vssd1 vccd1 vccd1 _1133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1064_ _1137_/CLK _1064_/D vssd1 vssd1 vccd1 vccd1 _1064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0917_ _0917_/A vssd1 vssd1 vccd1 vccd1 _1128_/D sky130_fd_sc_hd__clkbuf_1
X_0779_ _1107_/Q _0947_/B vssd1 vssd1 vccd1 vccd1 _1044_/B sky130_fd_sc_hd__nand2_1
X_0848_ _0960_/A _0848_/B vssd1 vssd1 vccd1 vccd1 _0849_/A sky130_fd_sc_hd__and2_1
XFILLER_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0702_ input17/X _1078_/Q _0702_/S vssd1 vssd1 vccd1 vccd1 _0703_/B sky130_fd_sc_hd__mux2_1
X_0633_ _1159_/Q vssd1 vssd1 vccd1 vccd1 _0646_/S sky130_fd_sc_hd__clkbuf_2
X_0564_ _0564_/A _0564_/B vssd1 vssd1 vccd1 vccd1 _0565_/A sky130_fd_sc_hd__or2_1
XFILLER_0_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1047_ _1117_/CLK _1047_/D vssd1 vssd1 vccd1 vccd1 _1047_/Q sky130_fd_sc_hd__dfxtp_1
X_1116_ _1117_/CLK _1116_/D vssd1 vssd1 vccd1 vccd1 _1116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0616_ input16/X _1054_/Q _0622_/S vssd1 vssd1 vccd1 vccd1 _0617_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0547_ _0547_/A vssd1 vssd1 vccd1 vccd1 _1100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0748__A0 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0739__A0 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0881_ _0824_/A _0853_/A _0859_/X _0880_/X vssd1 vssd1 vccd1 vccd1 _0881_/X sky130_fd_sc_hd__o211a_1
X_0950_ _1136_/Q _1135_/Q _0962_/S vssd1 vssd1 vccd1 vccd1 _0951_/B sky130_fd_sc_hd__mux2_1
XANTENNA__0653__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0896__C1 _0843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 io_wbs_m2s_stb vssd1 vssd1 vccd1 vccd1 _0850_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1080_ _1110_/CLK _1080_/D vssd1 vssd1 vccd1 vccd1 _1080_/Q sky130_fd_sc_hd__dfxtp_1
X_0933_ _0940_/A _0929_/X _1132_/Q vssd1 vssd1 vccd1 vccd1 _0936_/B sky130_fd_sc_hd__a21o_1
X_0864_ _0860_/X _0863_/X _0804_/X vssd1 vssd1 vccd1 vccd1 _1118_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0795_ _0820_/A vssd1 vssd1 vccd1 vccd1 _0795_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0580_ _0580_/A vssd1 vssd1 vccd1 vccd1 _1046_/D sky130_fd_sc_hd__clkbuf_1
X_1132_ _1149_/CLK _1132_/D vssd1 vssd1 vccd1 vccd1 _1132_/Q sky130_fd_sc_hd__dfxtp_1
X_1063_ _1141_/CLK _1063_/D vssd1 vssd1 vccd1 vccd1 _1063_/Q sky130_fd_sc_hd__dfxtp_1
X_0916_ _0941_/A _0916_/B _0916_/C vssd1 vssd1 vccd1 vccd1 _0917_/A sky130_fd_sc_hd__and3_1
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0778_ _1153_/Q _1154_/Q _1156_/Q _1155_/Q vssd1 vssd1 vccd1 vccd1 _0947_/B sky130_fd_sc_hd__nor4_1
X_0847_ _0569_/B _1023_/C _0846_/X _1117_/Q vssd1 vssd1 vccd1 vccd1 _0848_/B sky130_fd_sc_hd__a22o_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0563_ _1056_/Q _1106_/Q _0563_/S vssd1 vssd1 vccd1 vccd1 _0564_/B sky130_fd_sc_hd__mux2_1
X_0701_ _0722_/A vssd1 vssd1 vccd1 vccd1 _0720_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0632_ _0722_/A vssd1 vssd1 vccd1 vccd1 _0647_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1046_ _1117_/CLK _1046_/D vssd1 vssd1 vccd1 vccd1 _1046_/Q sky130_fd_sc_hd__dfxtp_1
X_1115_ _1152_/CLK _1115_/D vssd1 vssd1 vccd1 vccd1 _1115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0615_ _0615_/A vssd1 vssd1 vccd1 vccd1 _1053_/D sky130_fd_sc_hd__clkbuf_1
X_0546_ _0544_/X _1101_/Q _0558_/S vssd1 vssd1 vccd1 vccd1 _0547_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1029_ _1029_/A vssd1 vssd1 vccd1 vccd1 _1153_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_12_0_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _1143_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0529_ _1098_/Q _0563_/S vssd1 vssd1 vccd1 vccd1 _0529_/X sky130_fd_sc_hd__and2_1
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0880_ _1076_/Q _0865_/X _0866_/X _1061_/Q _0867_/X vssd1 vssd1 vccd1 vccd1 _0880_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0932_ _0932_/A vssd1 vssd1 vccd1 vccd1 _1131_/D sky130_fd_sc_hd__clkbuf_1
X_0863_ _1065_/Q _0878_/B vssd1 vssd1 vccd1 vccd1 _0863_/X sky130_fd_sc_hd__and2_1
X_0794_ _1108_/Q _0794_/B vssd1 vssd1 vccd1 vccd1 _0794_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1131_ _1149_/CLK _1131_/D vssd1 vssd1 vccd1 vccd1 _1131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1062_ _1141_/CLK _1062_/D vssd1 vssd1 vccd1 vccd1 _1062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0915_ _1031_/A _0920_/B _0914_/X vssd1 vssd1 vccd1 vccd1 _0916_/C sky130_fd_sc_hd__o21ai_1
X_0777_ _1037_/C vssd1 vssd1 vccd1 vccd1 _1044_/A sky130_fd_sc_hd__clkbuf_2
X_0846_ _1116_/Q _1115_/Q _0846_/C _0846_/D vssd1 vssd1 vccd1 vccd1 _0846_/X sky130_fd_sc_hd__or4_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0700_ _0700_/A vssd1 vssd1 vccd1 vccd1 _1077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0562_ _0562_/A vssd1 vssd1 vccd1 vccd1 _1105_/D sky130_fd_sc_hd__clkbuf_1
X_0631_ _0631_/A vssd1 vssd1 vccd1 vccd1 _1058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1114_ _1152_/CLK _1114_/D vssd1 vssd1 vccd1 vccd1 _1114_/Q sky130_fd_sc_hd__dfxtp_1
X_1045_ _1106_/CLK _1045_/D vssd1 vssd1 vccd1 vccd1 _1045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0829_ _0564_/A _0825_/Y _0826_/Y _0839_/C _0584_/A vssd1 vssd1 vccd1 vccd1 _1113_/D
+ sky130_fd_sc_hd__a221oi_1
XFILLER_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0923__C1 _0922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0614_ _0630_/A _0614_/B vssd1 vssd1 vccd1 vccd1 _0615_/A sky130_fd_sc_hd__and2_1
X_0545_ _0569_/B vssd1 vssd1 vccd1 vccd1 _0558_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1028_ _1025_/Y _1027_/Y _1153_/Q vssd1 vssd1 vccd1 vccd1 _1029_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0675__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0528_ _0560_/S vssd1 vssd1 vccd1 vccd1 _0563_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input11_A io_wbs_m2s_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_A io_wbs_m2s_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0931_ _0941_/A _0931_/B _0931_/C vssd1 vssd1 vccd1 vccd1 _0932_/A sky130_fd_sc_hd__and3_1
X_0862_ _0891_/B vssd1 vssd1 vccd1 vccd1 _0878_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0793_ _1044_/A _1044_/B _0976_/A _0674_/X vssd1 vssd1 vccd1 vccd1 _1107_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1130_ _1149_/CLK _1130_/D vssd1 vssd1 vccd1 vccd1 _1130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1061_ _1141_/CLK _1061_/D vssd1 vssd1 vccd1 vccd1 _1061_/Q sky130_fd_sc_hd__dfxtp_1
X_0914_ _0914_/A vssd1 vssd1 vccd1 vccd1 _0914_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0845_ _0845_/A vssd1 vssd1 vccd1 vccd1 _0960_/A sky130_fd_sc_hd__buf_2
X_0776_ _0992_/A _1007_/B _0946_/C vssd1 vssd1 vccd1 vccd1 _1037_/C sky130_fd_sc_hd__or3_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0702__A0 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0561_ _0560_/X _1106_/Q _0569_/B vssd1 vssd1 vccd1 vccd1 _0562_/A sky130_fd_sc_hd__mux2_1
X_0630_ _0630_/A _0630_/B vssd1 vssd1 vccd1 vccd1 _0631_/A sky130_fd_sc_hd__and2_1
X_1044_ _1044_/A _1044_/B vssd1 vssd1 vccd1 vccd1 _1159_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1113_ _1117_/CLK _1113_/D vssd1 vssd1 vccd1 vccd1 _1113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0759_ _0758_/Y _0748_/S _0584_/A vssd1 vssd1 vccd1 vccd1 _0759_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0828_ _0846_/D vssd1 vssd1 vccd1 vccd1 _0839_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0613_ input15/X _1053_/Q _0622_/S vssd1 vssd1 vccd1 vccd1 _0614_/B sky130_fd_sc_hd__mux2_1
X_1176__49 vssd1 vssd1 vccd1 vccd1 _1176__49/HI io_wbs_data_o[24] sky130_fd_sc_hd__conb_1
X_0544_ _1050_/Q _1100_/Q _0557_/S vssd1 vssd1 vccd1 vccd1 _0544_/X sky130_fd_sc_hd__mux2_1
X_1027_ _1027_/A _1027_/B vssd1 vssd1 vccd1 vccd1 _1027_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_6_0_clock clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 _1095_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_29_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0527_ _1073_/Q _0827_/C vssd1 vssd1 vccd1 vccd1 _0560_/S sky130_fd_sc_hd__nand2_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0593__A _0850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0768__A _0850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1160__33 vssd1 vssd1 vccd1 vccd1 _1160__33/HI io_wbs_data_o[8] sky130_fd_sc_hd__conb_1
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_3_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_0930_ _1026_/A _0929_/X _0914_/X vssd1 vssd1 vccd1 vccd1 _0931_/C sky130_fd_sc_hd__o21ai_1
X_0792_ _1027_/A vssd1 vssd1 vccd1 vccd1 _0976_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0861_ input3/X _0861_/B _0861_/C _0861_/D vssd1 vssd1 vccd1 vccd1 _0891_/B sky130_fd_sc_hd__and4_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1060_ _1137_/CLK _1060_/D vssd1 vssd1 vccd1 vccd1 _1060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0913_ _1128_/Q _0913_/B _1126_/Q vssd1 vssd1 vccd1 vccd1 _0920_/B sky130_fd_sc_hd__and3_1
X_0775_ _1152_/Q _1151_/Q _1150_/Q vssd1 vssd1 vccd1 vccd1 _0946_/C sky130_fd_sc_hd__or3_1
X_0844_ _0534_/B _1023_/C _0842_/Y _0843_/X vssd1 vssd1 vccd1 vccd1 _1116_/D sky130_fd_sc_hd__o211a_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0560_ _1055_/Q _1105_/Q _0560_/S vssd1 vssd1 vccd1 vccd1 _0560_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1043_ _0629_/S _1042_/X _0664_/X vssd1 vssd1 vccd1 vccd1 _1158_/D sky130_fd_sc_hd__o21a_1
X_1112_ _1117_/CLK _1112_/D vssd1 vssd1 vccd1 vccd1 _1112_/Q sky130_fd_sc_hd__dfxtp_1
X_0758_ _1093_/Q vssd1 vssd1 vccd1 vccd1 _0758_/Y sky130_fd_sc_hd__inv_2
X_0827_ _1113_/Q _1112_/Q _0827_/C _0827_/D vssd1 vssd1 vccd1 vccd1 _0846_/D sky130_fd_sc_hd__or4_1
XFILLER_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0689_ input13/X _1074_/Q _0702_/S vssd1 vssd1 vccd1 vccd1 _0690_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_2_0_clock clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 _1121_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0612_ _0722_/A vssd1 vssd1 vccd1 vccd1 _0630_/A sky130_fd_sc_hd__clkbuf_2
X_0543_ _0560_/S vssd1 vssd1 vccd1 vccd1 _0557_/S sky130_fd_sc_hd__clkbuf_2
X_1026_ _1026_/A _1037_/C vssd1 vssd1 vccd1 vccd1 _1027_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0602__A0 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0526_ _1045_/Q _1046_/Q _1048_/Q _1047_/Q vssd1 vssd1 vccd1 vccd1 _0827_/C sky130_fd_sc_hd__nor4_1
X_1009_ _1012_/B _1009_/B vssd1 vssd1 vccd1 vccd1 _1009_/Y sky130_fd_sc_hd__nor2_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0593__B _0593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0791_ _0988_/A vssd1 vssd1 vccd1 vccd1 _1027_/A sky130_fd_sc_hd__clkbuf_2
X_0860_ _0799_/B _0853_/X _0857_/X _0859_/X vssd1 vssd1 vccd1 vccd1 _0860_/X sky130_fd_sc_hd__o211a_1
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0989_ _0999_/C _0988_/X _0999_/B vssd1 vssd1 vccd1 vccd1 _0989_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0912_ _1026_/A vssd1 vssd1 vccd1 vccd1 _1031_/A sky130_fd_sc_hd__clkbuf_2
X_0774_ _1149_/Q _1148_/Q _1147_/Q vssd1 vssd1 vccd1 vccd1 _1007_/B sky130_fd_sc_hd__or3_1
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0843_ _0922_/A vssd1 vssd1 vccd1 vccd1 _0843_/X sky130_fd_sc_hd__buf_2
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1042_ input11/X _1158_/Q _1042_/S vssd1 vssd1 vccd1 vccd1 _1042_/X sky130_fd_sc_hd__mux2_1
X_1111_ _1152_/CLK _1111_/D vssd1 vssd1 vccd1 vccd1 _1111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0757_ _0757_/A vssd1 vssd1 vccd1 vccd1 _1092_/D sky130_fd_sc_hd__clkbuf_1
X_0688_ _0705_/S vssd1 vssd1 vccd1 vccd1 _0702_/S sky130_fd_sc_hd__clkbuf_2
X_0826_ _0821_/A _0821_/B _1113_/Q vssd1 vssd1 vccd1 vccd1 _0826_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0542_ _0542_/A vssd1 vssd1 vccd1 vccd1 _1099_/D sky130_fd_sc_hd__clkbuf_1
X_0611_ _0611_/A vssd1 vssd1 vccd1 vccd1 _0722_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1025_ _1037_/A _1037_/C vssd1 vssd1 vccd1 vccd1 _1025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0809_ _0795_/Y _0986_/B _0811_/B vssd1 vssd1 vccd1 vccd1 _0809_/X sky130_fd_sc_hd__a21o_1
XANTENNA__0669__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1181__54 vssd1 vssd1 vccd1 vccd1 _1181__54/HI io_wbs_data_o[29] sky130_fd_sc_hd__conb_1
XFILLER_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0525_ _1157_/Q _1081_/Q _1074_/Q _1082_/Q _0524_/X vssd1 vssd1 vccd1 vccd1 _0525_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1008_ _1148_/Q _1147_/Q _1007_/A _1149_/Q vssd1 vssd1 vccd1 vccd1 _1009_/B sky130_fd_sc_hd__o31a_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0592__A_N input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0732__A0 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0790_ _0784_/X _0787_/X _0789_/Y _1107_/Q vssd1 vssd1 vccd1 vccd1 _0988_/A sky130_fd_sc_hd__a31o_1
XANTENNA__0971__A0 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0723__A0 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0988_ _0988_/A vssd1 vssd1 vccd1 vccd1 _0988_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input1_A io_rxd vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0705__A0 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0911_ _1107_/Q vssd1 vssd1 vccd1 vccd1 _1026_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0842_ _1116_/Q _0842_/B vssd1 vssd1 vccd1 vccd1 _0842_/Y sky130_fd_sc_hd__xnor2_1
X_0773_ _1146_/Q _1145_/Q _1144_/Q _1143_/Q vssd1 vssd1 vccd1 vccd1 _0992_/A sky130_fd_sc_hd__or4_1
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ _1110_/CLK _1110_/D vssd1 vssd1 vccd1 vccd1 _1110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1041_ _0629_/S _1039_/X _1040_/X _0922_/X vssd1 vssd1 vccd1 vccd1 _1157_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0825_ _1093_/Q _0825_/B vssd1 vssd1 vccd1 vccd1 _0825_/Y sky130_fd_sc_hd__xnor2_1
X_0756_ _0766_/A _0756_/B vssd1 vssd1 vccd1 vccd1 _0757_/A sky130_fd_sc_hd__and2_1
X_0687_ _1159_/Q _1042_/S vssd1 vssd1 vccd1 vccd1 _0705_/S sky130_fd_sc_hd__or2_1
XFILLER_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0844__C1 _0843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0541_ _0540_/X _1100_/Q _0564_/A vssd1 vssd1 vccd1 vccd1 _0542_/A sky130_fd_sc_hd__mux2_1
X_0610_ _0610_/A vssd1 vssd1 vccd1 vccd1 _1052_/D sky130_fd_sc_hd__clkbuf_1
X_1024_ _1022_/X _1023_/Y _0822_/X vssd1 vssd1 vccd1 vccd1 _1152_/D sky130_fd_sc_hd__a21oi_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_1_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0808_ _1110_/Q _0808_/B vssd1 vssd1 vccd1 vccd1 _0811_/B sky130_fd_sc_hd__or2_1
X_0739_ input11/X _0799_/B _0748_/S vssd1 vssd1 vccd1 vccd1 _0740_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0524_ _1158_/Q _1080_/Q _1075_/Q _1083_/Q _0523_/X vssd1 vssd1 vccd1 vccd1 _0524_/X
+ sky130_fd_sc_hd__a221o_1
X_1007_ _1007_/A _1007_/B vssd1 vssd1 vccd1 vccd1 _1012_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0987_ _0999_/B _0999_/C _0987_/C _0987_/D vssd1 vssd1 vccd1 vccd1 _0987_/Y sky130_fd_sc_hd__nand4_1
XFILLER_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0910_ _0913_/B _0902_/A _0914_/A _1128_/Q vssd1 vssd1 vccd1 vccd1 _0916_/B sky130_fd_sc_hd__a31o_1
X_0841_ _1095_/Q _1006_/C vssd1 vssd1 vccd1 vccd1 _1023_/C sky130_fd_sc_hd__nor2_2
X_0772_ _0772_/A vssd1 vssd1 vccd1 vccd1 _1097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1040_ _1157_/Q _0629_/S vssd1 vssd1 vccd1 vccd1 _1040_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0755_ input15/X _0824_/A _0765_/S vssd1 vssd1 vccd1 vccd1 _0756_/B sky130_fd_sc_hd__mux2_1
X_0824_ _0824_/A _0832_/D vssd1 vssd1 vccd1 vccd1 _0825_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0686_ _0686_/A _0686_/B _0708_/B _0855_/C vssd1 vssd1 vccd1 vccd1 _1042_/S sky130_fd_sc_hd__or4b_2
XANTENNA__0605__A0 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0540_ _1049_/Q _1099_/Q _0563_/S vssd1 vssd1 vccd1 vccd1 _0540_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1023_ _1023_/A _1023_/B _1023_/C vssd1 vssd1 vccd1 vccd1 _1023_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_3_5_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0807_ _0807_/A _0807_/B vssd1 vssd1 vccd1 vccd1 _0986_/B sky130_fd_sc_hd__xnor2_1
X_0738_ _0765_/S vssd1 vssd1 vccd1 vccd1 _0748_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0669_ input13/X _0657_/X _0668_/X _0664_/X vssd1 vssd1 vccd1 vccd1 _1067_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1125__D _1125_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1172__45 vssd1 vssd1 vccd1 vccd1 _1172__45/HI io_wbs_data_o[20] sky130_fd_sc_hd__conb_1
X_0523_ _1085_/Q _1077_/Q _1076_/Q _1084_/Q _0522_/X vssd1 vssd1 vccd1 vccd1 _0523_/X
+ sky130_fd_sc_hd__a221o_1
X_1006_ _0833_/A _1006_/B _1006_/C vssd1 vssd1 vccd1 vccd1 _1006_/X sky130_fd_sc_hd__and3b_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0986_ _1023_/A _0986_/B vssd1 vssd1 vccd1 vccd1 _0987_/D sky130_fd_sc_hd__nand2_1
XFILLER_27_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0771_ _0822_/A _0771_/B vssd1 vssd1 vccd1 vccd1 _0772_/A sky130_fd_sc_hd__or2_1
X_0840_ _0564_/A _0837_/X _0838_/Y _0842_/B _0584_/A vssd1 vssd1 vccd1 vccd1 _1115_/D
+ sky130_fd_sc_hd__a221oi_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0969_ _0972_/A _0969_/B vssd1 vssd1 vccd1 vccd1 _0970_/A sky130_fd_sc_hd__and2_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0754_ _1092_/Q vssd1 vssd1 vccd1 vccd1 _0824_/A sky130_fd_sc_hd__clkbuf_2
X_0685_ input4/X input3/X input2/X vssd1 vssd1 vccd1 vccd1 _0855_/C sky130_fd_sc_hd__nor3b_1
X_0823_ _0817_/Y _0821_/X _0822_/X vssd1 vssd1 vccd1 vccd1 _1112_/D sky130_fd_sc_hd__a21oi_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1099_ _1106_/CLK _1099_/D vssd1 vssd1 vccd1 vccd1 _1099_/Q sky130_fd_sc_hd__dfxtp_1
X_1178__51 vssd1 vssd1 vccd1 vccd1 _1178__51/HI io_wbs_data_o[26] sky130_fd_sc_hd__conb_1
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1022_ _1017_/Y _1013_/A _1027_/A _1021_/Y vssd1 vssd1 vccd1 vccd1 _1022_/X sky130_fd_sc_hd__a31o_1
XFILLER_39_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0668_ _1067_/Q _0672_/B vssd1 vssd1 vccd1 vccd1 _0668_/X sky130_fd_sc_hd__or2_1
X_0737_ _0737_/A _0858_/B _0856_/C vssd1 vssd1 vccd1 vccd1 _0765_/S sky130_fd_sc_hd__or3b_4
X_0806_ _1110_/Q _0808_/B vssd1 vssd1 vccd1 vccd1 _0806_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0599_ _0887_/A _0599_/B vssd1 vssd1 vccd1 vccd1 _0600_/A sky130_fd_sc_hd__and2_1
XANTENNA__0762__A0 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0522_ _1087_/Q _1079_/Q _1078_/Q _1086_/Q vssd1 vssd1 vccd1 vccd1 _0522_/X sky130_fd_sc_hd__a22o_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1005_ _1002_/X _1003_/X _1004_/X vssd1 vssd1 vccd1 vccd1 _1148_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__0744__A0 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput30 _1123_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0726__A0 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

