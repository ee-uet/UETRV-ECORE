* NGSPICE file created from Core.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

.subckt Core clock io_dbus_addr[0] io_dbus_addr[10] io_dbus_addr[11] io_dbus_addr[12]
+ io_dbus_addr[13] io_dbus_addr[14] io_dbus_addr[15] io_dbus_addr[16] io_dbus_addr[17]
+ io_dbus_addr[18] io_dbus_addr[19] io_dbus_addr[1] io_dbus_addr[20] io_dbus_addr[21]
+ io_dbus_addr[22] io_dbus_addr[23] io_dbus_addr[24] io_dbus_addr[25] io_dbus_addr[26]
+ io_dbus_addr[27] io_dbus_addr[28] io_dbus_addr[29] io_dbus_addr[2] io_dbus_addr[30]
+ io_dbus_addr[31] io_dbus_addr[3] io_dbus_addr[4] io_dbus_addr[5] io_dbus_addr[6]
+ io_dbus_addr[7] io_dbus_addr[8] io_dbus_addr[9] io_dbus_ld_type[0] io_dbus_ld_type[1]
+ io_dbus_ld_type[2] io_dbus_rd_en io_dbus_rdata[0] io_dbus_rdata[10] io_dbus_rdata[11]
+ io_dbus_rdata[12] io_dbus_rdata[13] io_dbus_rdata[14] io_dbus_rdata[15] io_dbus_rdata[16]
+ io_dbus_rdata[17] io_dbus_rdata[18] io_dbus_rdata[19] io_dbus_rdata[1] io_dbus_rdata[20]
+ io_dbus_rdata[21] io_dbus_rdata[22] io_dbus_rdata[23] io_dbus_rdata[24] io_dbus_rdata[25]
+ io_dbus_rdata[26] io_dbus_rdata[27] io_dbus_rdata[28] io_dbus_rdata[29] io_dbus_rdata[2]
+ io_dbus_rdata[30] io_dbus_rdata[31] io_dbus_rdata[3] io_dbus_rdata[4] io_dbus_rdata[5]
+ io_dbus_rdata[6] io_dbus_rdata[7] io_dbus_rdata[8] io_dbus_rdata[9] io_dbus_st_type[0]
+ io_dbus_st_type[1] io_dbus_valid io_dbus_wdata[0] io_dbus_wdata[10] io_dbus_wdata[11]
+ io_dbus_wdata[12] io_dbus_wdata[13] io_dbus_wdata[14] io_dbus_wdata[15] io_dbus_wdata[16]
+ io_dbus_wdata[17] io_dbus_wdata[18] io_dbus_wdata[19] io_dbus_wdata[1] io_dbus_wdata[20]
+ io_dbus_wdata[21] io_dbus_wdata[22] io_dbus_wdata[23] io_dbus_wdata[24] io_dbus_wdata[25]
+ io_dbus_wdata[26] io_dbus_wdata[27] io_dbus_wdata[28] io_dbus_wdata[29] io_dbus_wdata[2]
+ io_dbus_wdata[30] io_dbus_wdata[31] io_dbus_wdata[3] io_dbus_wdata[4] io_dbus_wdata[5]
+ io_dbus_wdata[6] io_dbus_wdata[7] io_dbus_wdata[8] io_dbus_wdata[9] io_dbus_wr_en
+ io_ibus_addr[0] io_ibus_addr[10] io_ibus_addr[11] io_ibus_addr[12] io_ibus_addr[13]
+ io_ibus_addr[14] io_ibus_addr[15] io_ibus_addr[16] io_ibus_addr[17] io_ibus_addr[18]
+ io_ibus_addr[19] io_ibus_addr[1] io_ibus_addr[20] io_ibus_addr[21] io_ibus_addr[22]
+ io_ibus_addr[23] io_ibus_addr[24] io_ibus_addr[25] io_ibus_addr[26] io_ibus_addr[27]
+ io_ibus_addr[28] io_ibus_addr[29] io_ibus_addr[2] io_ibus_addr[30] io_ibus_addr[31]
+ io_ibus_addr[3] io_ibus_addr[4] io_ibus_addr[5] io_ibus_addr[6] io_ibus_addr[7]
+ io_ibus_addr[8] io_ibus_addr[9] io_ibus_inst[0] io_ibus_inst[10] io_ibus_inst[11]
+ io_ibus_inst[12] io_ibus_inst[13] io_ibus_inst[14] io_ibus_inst[15] io_ibus_inst[16]
+ io_ibus_inst[17] io_ibus_inst[18] io_ibus_inst[19] io_ibus_inst[1] io_ibus_inst[20]
+ io_ibus_inst[21] io_ibus_inst[22] io_ibus_inst[23] io_ibus_inst[24] io_ibus_inst[25]
+ io_ibus_inst[26] io_ibus_inst[27] io_ibus_inst[28] io_ibus_inst[29] io_ibus_inst[2]
+ io_ibus_inst[30] io_ibus_inst[31] io_ibus_inst[3] io_ibus_inst[4] io_ibus_inst[5]
+ io_ibus_inst[6] io_ibus_inst[7] io_ibus_inst[8] io_ibus_inst[9] io_ibus_valid io_irq_motor_irq
+ io_irq_spi_irq io_irq_uart_irq reset vccd1 vssd1
XFILLER_79_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09671_ _10254_/A vssd1 vssd1 vccd1 vccd1 _09920_/S sky130_fd_sc_hd__buf_4
X_18869_ _19001_/CLK _18869_/D vssd1 vssd1 vccd1 vccd1 _18869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13083__A2 _13081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10841__A1 _09547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15780__A1 _14750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12346__A1 _12338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14181__A _14189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10452__S0 _10180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09938_ _10277_/S vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__buf_2
XANTENNA__16600__S _16602_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17037__A1 _17036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15724__B _15732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09869_ _20038_/Q _19876_/Q _19285_/Q _19055_/Q _09635_/X _09639_/X vssd1 vssd1 vccd1
+ vccd1 _09869_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _18713_/Q _17096_/B _11887_/Y _11899_/X vssd1 vssd1 vccd1 vccd1 _11900_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _13048_/B vssd1 vssd1 vccd1 vccd1 _12880_/X sky130_fd_sc_hd__buf_2
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11831_/A vssd1 vssd1 vccd1 vccd1 _11831_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10507__S1 _10492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16836__A _16836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11045__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _13519_/B _14547_/X _14507_/X vssd1 vssd1 vccd1 vccd1 _14550_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11897_/A _19012_/Q vssd1 vssd1 vccd1 vccd1 _11762_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _17735_/A vssd1 vssd1 vccd1 vccd1 _13501_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11180__S1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10713_ _09624_/A _10711_/X _10712_/X vssd1 vssd1 vccd1 vccd1 _10713_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _14514_/A _14485_/C vssd1 vssd1 vccd1 vccd1 _14481_/Y sky130_fd_sc_hd__nor2_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16047__S _16053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _18662_/Q _13081_/A _12890_/A _14493_/B vssd1 vssd1 vccd1 vccd1 _11693_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16220_ _16220_/A vssd1 vssd1 vccd1 vccd1 _19126_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12034__A0 _18971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13432_ _18482_/Q _12943_/X _12944_/X _18706_/Q _13431_/X vssd1 vssd1 vccd1 vccd1
+ _13432_/X sky130_fd_sc_hd__a221o_1
X_10644_ _19144_/Q _19405_/Q _19304_/Q _19639_/Q _09726_/A _10626_/X vssd1 vssd1 vccd1
+ vccd1 _10644_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12585__A1 _18539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16151_ _17426_/A _18280_/B vssd1 vssd1 vccd1 vccd1 _16208_/A sky130_fd_sc_hd__or2_4
XFILLER_166_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10575_ _10690_/A _10574_/X _10149_/A vssd1 vssd1 vccd1 vccd1 _10575_/X sky130_fd_sc_hd__a21o_1
X_13363_ _13005_/X _13359_/X _13361_/X _13362_/X vssd1 vssd1 vccd1 vccd1 _17071_/A
+ sky130_fd_sc_hd__o31a_4
XANTENNA__16571__A _16617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_23_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15102_ _15102_/A vssd1 vssd1 vccd1 vccd1 _15102_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_154_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12314_ _14812_/B _12587_/A vssd1 vssd1 vccd1 vccd1 _12428_/A sky130_fd_sc_hd__or2_2
XFILLER_170_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16082_ _16082_/A vssd1 vssd1 vccd1 vccd1 _19064_/D sky130_fd_sc_hd__clkbuf_1
X_13294_ _18666_/Q _13081_/X _13082_/X _18734_/Q vssd1 vssd1 vccd1 vccd1 _13294_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15033_ _14887_/X _14862_/X _15039_/S vssd1 vssd1 vccd1 vccd1 _15033_/X sky130_fd_sc_hd__mux2_1
X_19910_ _19910_/CLK _19910_/D vssd1 vssd1 vccd1 vccd1 _19910_/Q sky130_fd_sc_hd__dfxtp_1
X_12245_ _12220_/A _12220_/B _12244_/X vssd1 vssd1 vccd1 vccd1 _12246_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10348__B1 _09823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12888__A2 _11732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19841_ _19942_/CLK _19841_/D vssd1 vssd1 vccd1 vccd1 _19841_/Q sky130_fd_sc_hd__dfxtp_1
X_12176_ _12658_/A _12831_/B _12260_/C _09263_/A vssd1 vssd1 vccd1 vccd1 _15219_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_122_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17606__S _17606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _19661_/Q _19427_/Q _18492_/Q _19757_/Q _11258_/S _10983_/X vssd1 vssd1 vccd1
+ vccd1 _11127_/X sky130_fd_sc_hd__mux4_1
X_19772_ _19868_/CLK _19772_/D vssd1 vssd1 vccd1 vccd1 _19772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16984_ _16390_/X _19449_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16985_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17028__A1 _17026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09913__A _09913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ _11058_/A vssd1 vssd1 vccd1 vccd1 _11058_/X sky130_fd_sc_hd__buf_2
XANTENNA__11848__B1 _11772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18723_ _18724_/CLK _18723_/D vssd1 vssd1 vccd1 vccd1 _18723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15935_ _19004_/Q _15927_/X _15928_/X _15934_/Y vssd1 vssd1 vccd1 vccd1 _19004_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10009_ _10009_/A vssd1 vssd1 vccd1 vccd1 _10010_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18654_ _18724_/CLK _18654_/D vssd1 vssd1 vccd1 vccd1 _18654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15866_ _15866_/A vssd1 vssd1 vccd1 vccd1 _18982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17605_ _17605_/A vssd1 vssd1 vccd1 vccd1 _19705_/D sky130_fd_sc_hd__clkbuf_1
X_14817_ _14869_/A vssd1 vssd1 vccd1 vccd1 _14956_/S sky130_fd_sc_hd__buf_2
XFILLER_91_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18585_ _18719_/CLK _18585_/D vssd1 vssd1 vccd1 vccd1 _18585_/Q sky130_fd_sc_hd__dfxtp_1
X_15797_ _15797_/A vssd1 vssd1 vccd1 vccd1 _18962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17536_ _19674_/Q vssd1 vssd1 vccd1 vccd1 _17537_/A sky130_fd_sc_hd__clkbuf_1
X_14748_ _15762_/A vssd1 vssd1 vccd1 vccd1 _14748_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17467_ _17467_/A vssd1 vssd1 vccd1 vccd1 _19640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14679_ _18792_/Q _13508_/B _14683_/S vssd1 vssd1 vccd1 vccd1 _14680_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19206_ _19959_/CLK _19206_/D vssd1 vssd1 vccd1 vccd1 _19206_/Q sky130_fd_sc_hd__dfxtp_1
X_16418_ _19198_/Q _13778_/X _16424_/S vssd1 vssd1 vccd1 vccd1 _16419_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17398_ _19610_/Q _17055_/X _17398_/S vssd1 vssd1 vccd1 vccd1 _17399_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19137_ _19986_/CLK _19137_/D vssd1 vssd1 vccd1 vccd1 _19137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16349_ _16381_/A vssd1 vssd1 vccd1 vccd1 _16362_/S sky130_fd_sc_hd__buf_4
XANTENNA__18172__S _18180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19068_ _20013_/CLK _19068_/D vssd1 vssd1 vccd1 vccd1 _19068_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15514__A1 _12717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18019_ _18019_/A vssd1 vssd1 vccd1 vccd1 _19875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12514__A _12514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16420__S _16424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09723_ _10906_/S vssd1 vssd1 vccd1 vccd1 _10859_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__09823__A _09823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11564__S _11566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09654_ _10449_/S vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ _10980_/A vssd1 vssd1 vccd1 vccd1 _09586_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11162__S1 _11015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12567__A1 _09468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10360_ _10365_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10360_/X sky130_fd_sc_hd__or2_1
XFILLER_136_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_197_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10291_ _19215_/Q _19806_/Q _19968_/Q _19183_/Q _10279_/X _10283_/X vssd1 vssd1 vccd1
+ vccd1 _10292_/B sky130_fd_sc_hd__mux4_2
X_12030_ _12078_/A _14865_/A _15094_/A vssd1 vssd1 vccd1 vccd1 _12031_/B sky130_fd_sc_hd__or3_2
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15735__A _15735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16330__S _16330_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13981_ _18567_/Q _13982_/C _18568_/Q vssd1 vssd1 vccd1 vccd1 _13983_/B sky130_fd_sc_hd__a21oi_1
XFILLER_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15720_ _15773_/B vssd1 vssd1 vccd1 vccd1 _15720_/X sky130_fd_sc_hd__clkbuf_2
X_12932_ _18647_/Q _12889_/X _12890_/X _14450_/B vssd1 vssd1 vccd1 vccd1 _12932_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _18904_/Q _18525_/Q _15655_/S vssd1 vssd1 vccd1 vccd1 _15652_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _12863_/A _12863_/B vssd1 vssd1 vccd1 vccd1 _12863_/Y sky130_fd_sc_hd__nor2_4
XFILLER_2_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18257__S _18263_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17161__S _17161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14602_ _12349_/A _11860_/D _14615_/S vssd1 vssd1 vccd1 vccd1 _14603_/B sky130_fd_sc_hd__mux2_1
XANTENNA__15470__A _15474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _17659_/X _20016_/Q _18374_/S vssd1 vssd1 vccd1 vccd1 _18371_/A sky130_fd_sc_hd__mux2_1
X_11814_ _18657_/Q vssd1 vssd1 vccd1 vccd1 _14280_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15582_/A vssd1 vssd1 vccd1 vccd1 _18873_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12448_/S _12792_/X _12813_/B _12154_/X vssd1 vssd1 vccd1 vccd1 _12794_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17321_ _17321_/A vssd1 vssd1 vccd1 vccd1 _19575_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14533_ _18746_/Q _13650_/A _11860_/C _14548_/A vssd1 vssd1 vccd1 vccd1 _14533_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _18567_/Q _13054_/B _11744_/X vssd1 vssd1 vccd1 vccd1 _11745_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17157_/X _19545_/Q _17254_/S vssd1 vssd1 vccd1 vccd1 _17253_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15744__A1 _09522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14464_ _18720_/Q _14461_/B _14463_/Y vssd1 vssd1 vccd1 vccd1 _18720_/D sky130_fd_sc_hd__o21a_1
X_11676_ _12060_/A _11700_/B vssd1 vssd1 vccd1 vccd1 _11677_/B sky130_fd_sc_hd__nor2_1
X_16203_ _16203_/A vssd1 vssd1 vccd1 vccd1 _19118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12558__A1 _18474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13415_ _18817_/Q _13269_/X _12879_/X _18784_/Q _13414_/X vssd1 vssd1 vccd1 vccd1
+ _13415_/X sky130_fd_sc_hd__a221o_1
X_10627_ _20025_/Q _19863_/Q _19272_/Q _19042_/Q _10691_/S _10626_/X vssd1 vssd1 vccd1
+ vccd1 _10628_/B sky130_fd_sc_hd__mux4_1
X_17183_ _17720_/A vssd1 vssd1 vccd1 vccd1 _17183_/X sky130_fd_sc_hd__clkbuf_1
X_14395_ _14398_/B _14398_/C _14366_/X vssd1 vssd1 vccd1 vccd1 _14395_/Y sky130_fd_sc_hd__a21oi_1
X_16134_ _16134_/A vssd1 vssd1 vccd1 vccd1 _19088_/D sky130_fd_sc_hd__clkbuf_1
X_13346_ _13346_/A vssd1 vssd1 vccd1 vccd1 _18446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09908__A _11574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10558_ _20026_/Q _19864_/Q _19273_/Q _19043_/Q _10125_/S _10492_/A vssd1 vssd1 vccd1
+ vccd1 _10558_/X sky130_fd_sc_hd__mux4_1
XFILLER_142_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16065_ _16065_/A vssd1 vssd1 vccd1 vccd1 _19059_/D sky130_fd_sc_hd__clkbuf_1
X_13277_ _18569_/Q _13070_/X _13272_/X _13274_/X _13276_/X vssd1 vssd1 vccd1 vccd1
+ _13657_/B sky130_fd_sc_hd__a2111o_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10489_ _09884_/A _10478_/X _10487_/X _09913_/A _10488_/Y vssd1 vssd1 vccd1 vccd1
+ _12850_/B sky130_fd_sc_hd__o32a_4
X_15016_ _15016_/A vssd1 vssd1 vccd1 vccd1 _15198_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__10416__S0 _10319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12228_ _12770_/S _12221_/A _12227_/X _12556_/A vssd1 vssd1 vccd1 vccd1 _12228_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19824_ _19824_/CLK _19824_/D vssd1 vssd1 vccd1 vccd1 _19824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12159_ _18460_/Q _12556_/A _12557_/A vssd1 vssd1 vccd1 vccd1 _12159_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10741__B1 _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19755_ _19755_/CLK _19755_/D vssd1 vssd1 vccd1 vccd1 _19755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16967_ _16364_/X _19441_/Q _16975_/S vssd1 vssd1 vccd1 vccd1 _16968_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18706_ _18744_/CLK _18706_/D vssd1 vssd1 vccd1 vccd1 _18706_/Q sky130_fd_sc_hd__dfxtp_1
X_15918_ _18999_/Q _15942_/A vssd1 vssd1 vccd1 vccd1 _15918_/X sky130_fd_sc_hd__and2_1
X_16898_ _16898_/A vssd1 vssd1 vccd1 vccd1 _19410_/D sky130_fd_sc_hd__clkbuf_1
X_19686_ _19842_/CLK _19686_/D vssd1 vssd1 vccd1 vccd1 _19686_/Q sky130_fd_sc_hd__dfxtp_1
X_15849_ _15871_/A _17203_/B vssd1 vssd1 vccd1 vccd1 _18977_/D sky130_fd_sc_hd__nor2_1
X_18637_ _18655_/CLK _18637_/D vssd1 vssd1 vccd1 vccd1 _18637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18167__S _18169_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09370_ _15773_/A _11680_/B _09378_/A vssd1 vssd1 vccd1 vccd1 _09394_/A sky130_fd_sc_hd__or3_2
X_18568_ _20005_/CLK _18568_/D vssd1 vssd1 vccd1 vccd1 _18568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15983__A1 _19025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09330__B_N _18940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11144__S1 _11015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17519_ _17519_/A vssd1 vssd1 vccd1 vccd1 _19665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18499_ _20022_/CLK _18499_/D vssd1 vssd1 vccd1 vccd1 _18499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17100__A _17199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__A _11166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17246__S _17254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09553__A _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__A _18848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09706_ _11145_/A vssd1 vssd1 vccd1 vccd1 _10952_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10496__C1 _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09637_ _09637_/A vssd1 vssd1 vccd1 vccd1 _10057_/A sky130_fd_sc_hd__buf_4
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13803__A _17039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _09568_/A vssd1 vssd1 vccd1 vccd1 _09568_/X sky130_fd_sc_hd__buf_2
XFILLER_71_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09499_ _09502_/A _09499_/B vssd1 vssd1 vccd1 vccd1 _11948_/A sky130_fd_sc_hd__nor2_1
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13014__S _13215_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ _11581_/A _11582_/B _11580_/C vssd1 vssd1 vccd1 vccd1 _11530_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10894__S0 _10892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11461_ _11606_/A _11606_/B _11606_/C vssd1 vssd1 vccd1 vccd1 _11462_/C sky130_fd_sc_hd__a21o_2
XFILLER_139_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13200_ _13005_/X _13186_/Y _13198_/X _13199_/X vssd1 vssd1 vccd1 vccd1 _17039_/A
+ sky130_fd_sc_hd__o31a_4
X_10412_ _18444_/Q _19473_/Q _19510_/Q _19084_/Q _10319_/X _10320_/X vssd1 vssd1 vccd1
+ vccd1 _10412_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17010__A _17010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14180_ _18632_/Q _18631_/Q _14180_/C vssd1 vssd1 vccd1 vccd1 _14182_/B sky130_fd_sc_hd__and3_1
X_11392_ _11388_/X _11390_/X _11391_/X _11435_/A vssd1 vssd1 vccd1 vccd1 _11392_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15449__B _15449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13131_ _18874_/Q _18875_/Q _13131_/C vssd1 vssd1 vccd1 vccd1 _13143_/B sky130_fd_sc_hd__and3_1
X_10343_ _19935_/Q _19549_/Q _19999_/Q _19118_/Q _10005_/A _10207_/A vssd1 vssd1 vccd1
+ vccd1 _10344_/B sky130_fd_sc_hd__mux4_1
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10274_ _09849_/X _10264_/X _10273_/X _09540_/X _18856_/Q vssd1 vssd1 vccd1 vccd1
+ _15966_/C sky130_fd_sc_hd__a32o_4
XANTENNA_input55_A io_ibus_inst[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ _13047_/Y _13061_/X _13350_/S vssd1 vssd1 vccd1 vccd1 _13062_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12013_ _12188_/A vssd1 vssd1 vccd1 vccd1 _13700_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17870_ _19809_/Q _17078_/X _17876_/S vssd1 vssd1 vccd1 vccd1 _17871_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11071__S0 _11049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16821_ _16821_/A vssd1 vssd1 vccd1 vccd1 _16830_/S sky130_fd_sc_hd__buf_4
XFILLER_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19540_ _19990_/CLK _19540_/D vssd1 vssd1 vccd1 vccd1 _19540_/Q sky130_fd_sc_hd__dfxtp_1
X_16752_ _19346_/Q _13842_/X _16758_/S vssd1 vssd1 vccd1 vccd1 _16753_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13964_ _18562_/Q _18561_/Q _13964_/C vssd1 vssd1 vccd1 vccd1 _13966_/B sky130_fd_sc_hd__and3_1
XFILLER_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15703_ _18928_/Q _18549_/Q _15703_/S vssd1 vssd1 vccd1 vccd1 _15704_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10487__C1 _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ _15735_/A _16691_/B _16150_/B vssd1 vssd1 vccd1 vccd1 _16993_/A sky130_fd_sc_hd__nand3_2
XFILLER_111_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19471_ _19865_/CLK _19471_/D vssd1 vssd1 vccd1 vccd1 _19471_/Q sky130_fd_sc_hd__dfxtp_1
X_16683_ _16390_/X _19316_/Q _16685_/S vssd1 vssd1 vccd1 vccd1 _16684_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13895_ _18537_/Q _13893_/X _12528_/X _12533_/Y _13890_/X vssd1 vssd1 vccd1 vccd1
+ _18537_/D sky130_fd_sc_hd__o221a_1
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18422_ _17735_/X _20040_/Q _18422_/S vssd1 vssd1 vccd1 vccd1 _18423_/A sky130_fd_sc_hd__mux2_1
X_15634_ _15690_/A vssd1 vssd1 vccd1 vccd1 _15703_/S sky130_fd_sc_hd__buf_4
XFILLER_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12846_ _12863_/A vssd1 vssd1 vccd1 vccd1 _12851_/A sky130_fd_sc_hd__buf_8
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_196_clock clkbuf_opt_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19978_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__A1 _14993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18353_ _18409_/A vssd1 vssd1 vccd1 vccd1 _18422_/S sky130_fd_sc_hd__buf_6
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15565_ _18866_/Q _18898_/Q _15567_/S vssd1 vssd1 vccd1 vccd1 _15566_/A sky130_fd_sc_hd__mux2_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ _12260_/A _12657_/X _12864_/C _11945_/A vssd1 vssd1 vccd1 vccd1 _12778_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17128_/X _19568_/Q _17304_/S vssd1 vssd1 vccd1 vccd1 _17305_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14518_/A _14518_/C _14507_/X vssd1 vssd1 vccd1 vccd1 _14516_/Y sky130_fd_sc_hd__a21oi_1
X_11728_ _18749_/Q _15715_/B _11728_/C vssd1 vssd1 vccd1 vccd1 _11728_/X sky130_fd_sc_hd__or3_1
X_18284_ _18284_/A vssd1 vssd1 vccd1 vccd1 _19977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10885__S0 _10704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15496_ _15101_/X _15498_/B _14994_/X _15495_/X vssd1 vssd1 vccd1 vccd1 _15496_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ _17131_/X _19537_/Q _17243_/S vssd1 vssd1 vccd1 vccd1 _17236_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14447_ _14450_/A _14447_/B vssd1 vssd1 vccd1 vccd1 _18714_/D sky130_fd_sc_hd__nor2_1
XFILLER_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ _14755_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _14812_/A sky130_fd_sc_hd__nor2_1
XANTENNA__14544__A input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17166_ _17166_/A vssd1 vssd1 vccd1 vccd1 _19510_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09638__A _10057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14378_ _18689_/Q _14378_/B _14378_/C vssd1 vssd1 vccd1 vccd1 _14384_/C sky130_fd_sc_hd__and3_1
XFILLER_171_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16117_ _16117_/A vssd1 vssd1 vccd1 vccd1 _19080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13329_ _18736_/Q vssd1 vssd1 vccd1 vccd1 _14510_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17097_ _17634_/A vssd1 vssd1 vccd1 vccd1 _17097_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_134_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18819_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16048_ _16048_/A vssd1 vssd1 vccd1 vccd1 _19052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17066__S _17072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19807_ _20034_/CLK _19807_/D vssd1 vssd1 vccd1 vccd1 _19807_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_149_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _18688_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15653__A0 _18905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17999_ _17999_/A vssd1 vssd1 vccd1 vccd1 _19866_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19738_ _19996_/CLK _19738_/D vssd1 vssd1 vccd1 vccd1 _19738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_145_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10478__C1 _09806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11365__S1 _11077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19669_ _20023_/CLK _19669_/D vssd1 vssd1 vccd1 vccd1 _19669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09422_ _11716_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09422_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09353_ _18828_/Q vssd1 vssd1 vccd1 vccd1 _09354_/A sky130_fd_sc_hd__inv_2
XFILLER_127_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10876__S0 _10776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09284_ _09284_/A _11919_/B _09284_/C vssd1 vssd1 vccd1 vccd1 _09287_/C sky130_fd_sc_hd__or3_1
XANTENNA__13769__S _13772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10982__A _11258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14454__A _14472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__A _19526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11745__A2 _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12155__C1 _12154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10921__S _10921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15644__A0 _18901_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10222__A _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15732__B _15732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10961_ _11295_/S vssd1 vssd1 vccd1 vccd1 _11023_/S sky130_fd_sc_hd__buf_2
XFILLER_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12700_ _18783_/Q _12700_/B vssd1 vssd1 vccd1 vccd1 _12750_/C sky130_fd_sc_hd__and2_1
XFILLER_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13680_ _18887_/Q _13681_/B vssd1 vssd1 vccd1 vccd1 _13693_/C sky130_fd_sc_hd__or2_2
X_10892_ _10892_/A vssd1 vssd1 vccd1 vccd1 _10892_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17149__A0 _17147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ _18541_/Q _12553_/X _12627_/X _12630_/Y vssd1 vssd1 vccd1 vccd1 _12631_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_54_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15350_ _15355_/A _15355_/B vssd1 vssd1 vccd1 vccd1 _15350_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12562_ _12562_/A _12582_/C vssd1 vssd1 vccd1 vccd1 _12562_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14301_ _18666_/Q _14306_/D _14792_/A vssd1 vssd1 vccd1 vccd1 _14302_/B sky130_fd_sc_hd__o21ai_1
X_11513_ _15947_/C _12844_/A vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__and2_1
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15281_ _15136_/X _15280_/X _15331_/S vssd1 vssd1 vccd1 vccd1 _15281_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16055__S _16057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12493_ _12493_/A _12519_/A vssd1 vssd1 vccd1 vccd1 _12497_/A sky130_fd_sc_hd__xor2_4
X_17020_ _17020_/A vssd1 vssd1 vccd1 vccd1 _17020_/X sky130_fd_sc_hd__clkbuf_1
X_14232_ _14232_/A vssd1 vssd1 vccd1 vccd1 _18646_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09458__A _09458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_51_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19829_/CLK sky130_fd_sc_hd__clkbuf_16
X_11444_ _11086_/A _11441_/X _11443_/X vssd1 vssd1 vccd1 vccd1 _11444_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12394__C1 _12012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11736__A2 _11815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17675__A _17675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ _18625_/Q _14164_/C _18626_/Q vssd1 vssd1 vccd1 vccd1 _14165_/B sky130_fd_sc_hd__a21oi_1
XFILLER_164_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18270__S _18274_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11375_ _11058_/A _11366_/Y _11370_/Y _11374_/Y _09872_/A vssd1 vssd1 vccd1 vccd1
+ _11375_/X sky130_fd_sc_hd__o311a_1
XFILLER_124_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13114_ _17023_/A vssd1 vssd1 vccd1 vccd1 _17665_/A sky130_fd_sc_hd__clkbuf_2
X_10326_ _18855_/Q _09540_/A _09547_/X _10325_/X vssd1 vssd1 vccd1 vccd1 _15964_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_125_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18971_ _19485_/CLK _18971_/D vssd1 vssd1 vccd1 vccd1 _18971_/Q sky130_fd_sc_hd__dfxtp_2
X_14094_ _14094_/A vssd1 vssd1 vccd1 vccd1 _14143_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14686__A1 _13546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output161_A _12728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_66_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19976_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _19832_/Q _17049_/X _17926_/S vssd1 vssd1 vccd1 vccd1 _17923_/A sky130_fd_sc_hd__mux2_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13046_/A _13046_/C _18872_/Q vssd1 vssd1 vccd1 vccd1 _13047_/A sky130_fd_sc_hd__a21oi_1
X_10257_ _10252_/Y _10255_/X _10256_/X _10365_/A vssd1 vssd1 vccd1 vccd1 _10257_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10188_ _10449_/S vssd1 vssd1 vccd1 vccd1 _10354_/S sky130_fd_sc_hd__buf_4
X_17853_ _17853_/A vssd1 vssd1 vccd1 vccd1 _19801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16804_ _16355_/X _19369_/Q _16808_/S vssd1 vssd1 vccd1 vccd1 _16805_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15923__A _15940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17784_ _17795_/A vssd1 vssd1 vccd1 vccd1 _17793_/S sky130_fd_sc_hd__buf_6
X_14996_ _15286_/A _14996_/B vssd1 vssd1 vccd1 vccd1 _14996_/X sky130_fd_sc_hd__or2_1
XFILLER_75_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19523_ _19523_/CLK _19523_/D vssd1 vssd1 vccd1 vccd1 _19523_/Q sky130_fd_sc_hd__dfxtp_1
X_16735_ _16735_/A vssd1 vssd1 vccd1 vccd1 _19338_/D sky130_fd_sc_hd__clkbuf_1
X_13947_ _18557_/Q _18556_/Q _18555_/Q _13947_/D vssd1 vssd1 vccd1 vccd1 _13958_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14539__A _16836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16666_ _16364_/X _19308_/Q _16674_/S vssd1 vssd1 vccd1 vccd1 _16667_/A sky130_fd_sc_hd__mux2_1
X_19454_ _19816_/CLK _19454_/D vssd1 vssd1 vccd1 vccd1 _19454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13878_ _12258_/A _12258_/B _13870_/X vssd1 vssd1 vccd1 vccd1 _18527_/D sky130_fd_sc_hd__a21o_1
XFILLER_62_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14258__B _14264_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18405_ _17710_/X _20032_/Q _18407_/S vssd1 vssd1 vccd1 vccd1 _18406_/A sky130_fd_sc_hd__mux2_1
X_15617_ _15617_/A vssd1 vssd1 vccd1 vccd1 _18889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10880__C1 _09874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ _12829_/A vssd1 vssd1 vccd1 vccd1 _12829_/X sky130_fd_sc_hd__clkbuf_1
X_16597_ _16597_/A vssd1 vssd1 vccd1 vccd1 _19277_/D sky130_fd_sc_hd__clkbuf_1
X_19385_ _19526_/CLK _19385_/D vssd1 vssd1 vccd1 vccd1 _19385_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18336_ _18336_/A vssd1 vssd1 vccd1 vccd1 _20001_/D sky130_fd_sc_hd__clkbuf_1
X_15548_ _15624_/A vssd1 vssd1 vccd1 vccd1 _15602_/A sky130_fd_sc_hd__buf_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18267_ _18267_/A vssd1 vssd1 vccd1 vccd1 _19970_/D sky130_fd_sc_hd__clkbuf_1
X_15479_ _15405_/X _15477_/X _15478_/X _14826_/A _12645_/X vssd1 vssd1 vccd1 vccd1
+ _15479_/X sky130_fd_sc_hd__a32o_1
XFILLER_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13177__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clock _18998_/CLK vssd1 vssd1 vccd1 vccd1 _19821_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14374__B1 _14366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17218_ _17218_/A vssd1 vssd1 vccd1 vccd1 _19529_/D sky130_fd_sc_hd__clkbuf_1
X_18198_ _17723_/X _19940_/Q _18202_/S vssd1 vssd1 vccd1 vccd1 _18199_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17149_ _17147_/X _19505_/Q _17161_/S vssd1 vssd1 vccd1 vccd1 _17150_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_71_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18180__S _18180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09971_ _09973_/A _09970_/X _09566_/A vssd1 vssd1 vccd1 vccd1 _09971_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14677__A1 _14562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12688__A0 _15972_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12522__A _12522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11783__D _15758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15833__A _15833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13101__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09831__A _10690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11112__B1 _11227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13652__A2 _13517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13353__A _17068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18040__A1 _18836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16051__A0 _13443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09405_ _09405_/A _09405_/B vssd1 vssd1 vccd1 vccd1 _09410_/C sky130_fd_sc_hd__nor2_1
XFILLER_81_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18355__S _18363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09336_ _09697_/C _09698_/A _09698_/B vssd1 vssd1 vccd1 vccd1 _09337_/C sky130_fd_sc_hd__and3_1
XFILLER_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09267_ _09434_/A _09436_/B _09435_/A _09267_/D vssd1 vssd1 vccd1 vccd1 _09275_/A
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__15157__A2 _15160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ _09198_/A vssd1 vssd1 vccd1 vccd1 _12003_/C sky130_fd_sc_hd__buf_2
XFILLER_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12416__B _12416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10217__A _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11160_ _19661_/Q _19427_/Q _18492_/Q _19757_/Q _09721_/A _11015_/X vssd1 vssd1 vccd1
+ vccd1 _11160_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10111_ _10411_/A _10111_/B vssd1 vssd1 vccd1 vccd1 _10111_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11091_ _11309_/A vssd1 vssd1 vccd1 vccd1 _11242_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13528__A _13656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10042_ _19345_/Q _19616_/Q _19840_/Q _19584_/Q _10275_/A _09747_/A vssd1 vssd1 vccd1
+ vccd1 _10042_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14850_ _15353_/A vssd1 vssd1 vccd1 vccd1 _15268_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13801_ _18499_/Q _13800_/X _13804_/S vssd1 vssd1 vccd1 vccd1 _13802_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11329__S1 _11322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input18_A io_dbus_rdata[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14781_ _14781_/A vssd1 vssd1 vccd1 vccd1 _18826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12578__S _12770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11993_ _11993_/A _11993_/B vssd1 vssd1 vccd1 vccd1 _11994_/A sky130_fd_sc_hd__xnor2_4
XFILLER_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14359__A _14407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ _16520_/A vssd1 vssd1 vccd1 vccd1 _19243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13732_ _13732_/A _19023_/Q vssd1 vssd1 vccd1 vccd1 _13732_/Y sky130_fd_sc_hd__nand2_1
X_10944_ _18433_/Q _19462_/Q _19499_/Q _19073_/Q _10892_/X _10893_/X vssd1 vssd1 vccd1
+ vccd1 _10944_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16451_ _19213_/Q _13826_/X _16457_/S vssd1 vssd1 vccd1 vccd1 _16452_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13663_ _18473_/Q _13517_/X _13655_/Y _13662_/X vssd1 vssd1 vccd1 vccd1 _18473_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10875_ _09664_/A _10872_/X _10874_/X vssd1 vssd1 vccd1 vccd1 _10875_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15402_ _15329_/X _15315_/X _15401_/X _15342_/X vssd1 vssd1 vccd1 vccd1 _15402_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ _19957_/CLK _19170_/D vssd1 vssd1 vccd1 vccd1 _19170_/Q sky130_fd_sc_hd__dfxtp_1
X_12614_ _15966_/C _18920_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12641_/A sky130_fd_sc_hd__mux2_2
XANTENNA__11406__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16382_ _16380_/X _19185_/Q _16394_/S vssd1 vssd1 vccd1 vccd1 _16383_/A sky130_fd_sc_hd__mux2_1
X_13594_ _13603_/C _13594_/B vssd1 vssd1 vccd1 vccd1 _13594_/Y sky130_fd_sc_hd__nand2_1
X_18121_ _18860_/Q _13719_/X _18130_/S vssd1 vssd1 vccd1 vccd1 _18121_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11501__S1 _10788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15333_ _15544_/A vssd1 vssd1 vccd1 vccd1 _15399_/A sky130_fd_sc_hd__clkbuf_1
X_12545_ _12545_/A _12545_/B vssd1 vssd1 vccd1 vccd1 _12550_/A sky130_fd_sc_hd__and2_2
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14094__A _14094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18052_ _18052_/A vssd1 vssd1 vccd1 vccd1 _19887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15264_ _14978_/X _15170_/X _15097_/X vssd1 vssd1 vccd1 vccd1 _15440_/B sky130_fd_sc_hd__o21a_1
XFILLER_157_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12476_ _18531_/Q _18532_/Q _12476_/C _12476_/D vssd1 vssd1 vccd1 vccd1 _12477_/D
+ sky130_fd_sc_hd__and4_1
X_17003_ _17003_/A vssd1 vssd1 vccd1 vccd1 _19455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14215_ _18644_/Q _14215_/B vssd1 vssd1 vccd1 vccd1 _14216_/B sky130_fd_sc_hd__and2_1
XANTENNA__17609__S _17617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11427_ _11414_/A _11426_/X _09681_/A vssd1 vssd1 vccd1 vccd1 _11427_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__15918__A _18999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16513__S _16519_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10068__S1 _09646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _15093_/X _15187_/X _15194_/X _15048_/X _12150_/Y vssd1 vssd1 vccd1 vccd1
+ _15195_/X sky130_fd_sc_hd__a32o_1
XANTENNA__14822__A _15368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output86_A _12621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09916__A _15978_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ _14146_/A _14153_/C vssd1 vssd1 vccd1 vccd1 _14146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11358_ _19322_/Q _19593_/Q _19817_/Q _19561_/Q _11356_/X _11357_/X vssd1 vssd1 vccd1
+ vccd1 _11359_/B sky130_fd_sc_hd__mux4_1
XANTENNA__14659__A1 _13733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10309_ _10305_/A _10308_/X _10107_/X vssd1 vssd1 vccd1 vccd1 _10309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_140_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14077_ _14078_/A _14078_/C _14076_/Y vssd1 vssd1 vccd1 vccd1 _18601_/D sky130_fd_sc_hd__o21a_1
X_18954_ _18956_/CLK _18954_/D vssd1 vssd1 vccd1 vccd1 _18954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11289_ _11278_/A _11288_/X _09682_/A vssd1 vssd1 vccd1 vccd1 _11289_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_112_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11568__S1 _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17905_ _17905_/A vssd1 vssd1 vccd1 vccd1 _19824_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _13046_/A _13046_/C vssd1 vssd1 vccd1 vccd1 _13028_/X sky130_fd_sc_hd__xor2_1
X_18885_ _19055_/CLK _18885_/D vssd1 vssd1 vccd1 vccd1 _18885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17344__S _17348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17836_ _17836_/A vssd1 vssd1 vccd1 vccd1 _19793_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11893__A1 _18606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09651__A _10655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10797__A _10953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17767_ _17675_/X _19763_/Q _17771_/S vssd1 vssd1 vccd1 vccd1 _17768_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_18_clock_A _18998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14831__A1 _12807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ _14993_/A _15201_/B vssd1 vssd1 vccd1 vccd1 _14979_/X sky130_fd_sc_hd__and2_1
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19506_ _20026_/CLK _19506_/D vssd1 vssd1 vccd1 vccd1 _19506_/Q sky130_fd_sc_hd__dfxtp_1
X_16718_ _16718_/A vssd1 vssd1 vccd1 vccd1 _19330_/D sky130_fd_sc_hd__clkbuf_1
X_17698_ _17697_/X _19738_/Q _17698_/S vssd1 vssd1 vccd1 vccd1 _17699_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19437_ _19767_/CLK _19437_/D vssd1 vssd1 vccd1 vccd1 _19437_/Q sky130_fd_sc_hd__dfxtp_1
X_16649_ _16649_/A vssd1 vssd1 vccd1 vccd1 _19300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19368_ _19960_/CLK _19368_/D vssd1 vssd1 vccd1 vccd1 _19368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18319_ _18319_/A vssd1 vssd1 vccd1 vccd1 _19993_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12070__A1 _12020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19299_ _20020_/CLK _19299_/D vssd1 vssd1 vccd1 vccd1 _19299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11256__S0 _11212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11030__C1 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09954_ _19683_/Q _19449_/Q _18514_/Q _19779_/Q _09939_/X _09940_/X vssd1 vssd1 vccd1
+ vccd1 _09954_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09885_ _09957_/A vssd1 vssd1 vccd1 vccd1 _11572_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14878__S _14948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13782__S _13788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17254__S _17254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09561__A _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14907__A _14907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13389__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ _10656_/X _10658_/X _10659_/X _10670_/A _09563_/A vssd1 vssd1 vccd1 vccd1
+ _10668_/B sky130_fd_sc_hd__o221a_1
XFILLER_167_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09319_ _09319_/A vssd1 vssd1 vccd1 vccd1 _11903_/A sky130_fd_sc_hd__buf_2
X_10591_ _10670_/A _10590_/X _09562_/A vssd1 vssd1 vccd1 vccd1 _10591_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_167_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12330_ _12330_/A vssd1 vssd1 vccd1 vccd1 _12334_/A sky130_fd_sc_hd__clkinv_2
X_12261_ _11904_/A _12837_/B _12260_/X vssd1 vssd1 vccd1 vccd1 _12323_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11247__S0 _11273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14000_ _14044_/A _14000_/B _14001_/B vssd1 vssd1 vccd1 vccd1 _18574_/D sky130_fd_sc_hd__nor3_1
X_11212_ _11212_/A vssd1 vssd1 vccd1 vccd1 _11212_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12192_ _12192_/A _12277_/D vssd1 vssd1 vccd1 vccd1 _12192_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11143_ _09848_/A _11133_/X _11142_/X _09537_/A _18839_/Q vssd1 vssd1 vccd1 vccd1
+ _15923_/C sky130_fd_sc_hd__a32o_4
XFILLER_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput75 _12364_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[13] sky130_fd_sc_hd__buf_2
XFILLER_110_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput86 _12621_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[23] sky130_fd_sc_hd__buf_2
XFILLER_95_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput97 _12094_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[4] sky130_fd_sc_hd__buf_2
X_11074_ _20016_/Q _19854_/Q _19263_/Q _19033_/Q _11063_/X _11073_/X vssd1 vssd1 vccd1
+ vccd1 _11075_/B sky130_fd_sc_hd__mux4_1
X_15951_ _15951_/A vssd1 vssd1 vccd1 vccd1 _15951_/X sky130_fd_sc_hd__buf_2
XFILLER_0_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10025_ _10037_/S vssd1 vssd1 vccd1 vccd1 _10095_/S sky130_fd_sc_hd__buf_2
X_14902_ _14996_/B _12783_/A _14933_/S vssd1 vssd1 vccd1 vccd1 _14902_/X sky130_fd_sc_hd__mux2_1
X_18670_ _18688_/CLK _18670_/D vssd1 vssd1 vccd1 vccd1 _18670_/Q sky130_fd_sc_hd__dfxtp_2
X_15882_ _15882_/A vssd1 vssd1 vccd1 vccd1 _18987_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16263__A0 _13238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17621_ _17621_/A vssd1 vssd1 vccd1 vccd1 _19712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ _14990_/A _15201_/B vssd1 vssd1 vccd1 vccd1 _14983_/B sky130_fd_sc_hd__nand2_2
XANTENNA_output124_A _12855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17552_ _19682_/Q vssd1 vssd1 vccd1 vccd1 _17553_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14764_ _14764_/A _14764_/B _14814_/A _14764_/D vssd1 vssd1 vccd1 vccd1 _14765_/D
+ sky130_fd_sc_hd__or4_1
X_11976_ _12193_/A _11999_/A _12001_/A vssd1 vssd1 vccd1 vccd1 _12050_/A sky130_fd_sc_hd__or3_1
X_16503_ _16503_/A vssd1 vssd1 vccd1 vccd1 _19235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13715_ _13714_/A _13714_/C _13714_/B vssd1 vssd1 vccd1 vccd1 _13715_/Y sky130_fd_sc_hd__o21ai_1
X_17483_ _17483_/A vssd1 vssd1 vccd1 vccd1 _17492_/S sky130_fd_sc_hd__buf_4
X_10927_ _10934_/A _10927_/B vssd1 vssd1 vccd1 vccd1 _10927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14695_ _14695_/A vssd1 vssd1 vccd1 vccd1 _18799_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16508__S _16508_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19222_ _19877_/CLK _19222_/D vssd1 vssd1 vccd1 vccd1 _19222_/Q sky130_fd_sc_hd__dfxtp_1
X_16434_ _16434_/A vssd1 vssd1 vccd1 vccd1 _19205_/D sky130_fd_sc_hd__clkbuf_1
X_13646_ _18882_/Q _18883_/Q _13646_/C vssd1 vssd1 vccd1 vccd1 _13654_/B sky130_fd_sc_hd__or3_2
XFILLER_158_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10858_ _10858_/A _10858_/B vssd1 vssd1 vccd1 vccd1 _10858_/X sky130_fd_sc_hd__or2_1
XFILLER_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _16381_/A vssd1 vssd1 vccd1 vccd1 _16378_/S sky130_fd_sc_hd__buf_6
X_19153_ _20002_/CLK _19153_/D vssd1 vssd1 vccd1 vccd1 _19153_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16318__A1 _19165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10289__S1 _10283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13577_ _19003_/Q _13577_/B vssd1 vssd1 vccd1 vccd1 _13577_/X sky130_fd_sc_hd__or2_1
X_10789_ _19204_/Q _19795_/Q _19957_/Q _19172_/Q _10787_/X _10788_/X vssd1 vssd1 vccd1
+ vccd1 _10790_/B sky130_fd_sc_hd__mux4_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18104_ _18104_/A vssd1 vssd1 vccd1 vccd1 _18118_/S sky130_fd_sc_hd__clkbuf_2
X_15316_ _15321_/A _15321_/B vssd1 vssd1 vccd1 vccd1 _15316_/Y sky130_fd_sc_hd__nand2_1
X_12528_ _12522_/X _12526_/X _12527_/X _12480_/X vssd1 vssd1 vccd1 vccd1 _12528_/X
+ sky130_fd_sc_hd__o211a_1
X_19084_ _19581_/CLK _19084_/D vssd1 vssd1 vccd1 vccd1 _19084_/Q sky130_fd_sc_hd__dfxtp_1
X_16296_ _16296_/A vssd1 vssd1 vccd1 vccd1 _19159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18035_ _18034_/X _19882_/Q _18044_/S vssd1 vssd1 vccd1 vccd1 _18036_/A sky130_fd_sc_hd__mux2_1
X_15247_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15247_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16243__S _16247_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ _12459_/A vssd1 vssd1 vccd1 vccd1 _12515_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14552__A _14552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09646__A _09646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15178_ _15517_/A _15178_/B vssd1 vssd1 vccd1 vccd1 _15178_/X sky130_fd_sc_hd__or2_1
XFILLER_153_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14129_ _18615_/Q _14125_/C _14128_/Y vssd1 vssd1 vccd1 vccd1 _18615_/D sky130_fd_sc_hd__o21a_1
XFILLER_114_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10461__S1 _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19986_ _19986_/CLK _19986_/D vssd1 vssd1 vccd1 vccd1 _19986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18937_ _18975_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _18937_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_67_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09670_ _10251_/S vssd1 vssd1 vccd1 vccd1 _10254_/A sky130_fd_sc_hd__buf_2
X_18868_ _18868_/CLK _18868_/D vssd1 vssd1 vccd1 vccd1 _18868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17819_ _19786_/Q _17004_/X _17821_/S vssd1 vssd1 vccd1 vccd1 _17820_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18799_ _19888_/CLK _18799_/D vssd1 vssd1 vccd1 vccd1 _18799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17802__S _17804_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10320__A _10492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16418__S _16424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10841__A2 _10830_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_clock clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_15_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10990__A _11212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10357__A1 _10054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15992__S _15998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17773__A _17795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10452__S1 _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15296__A1 _12301_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09937_ _09849_/X _09927_/X _09936_/X _09540_/X _18861_/Q vssd1 vssd1 vccd1 vccd1
+ _15976_/C sky130_fd_sc_hd__a32o_4
XFILLER_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11306__B1 _11181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13806__A _17042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09868_ _09868_/A _09868_/B vssd1 vssd1 vccd1 vccd1 _09868_/X sky130_fd_sc_hd__or2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09799_/A vssd1 vssd1 vccd1 vccd1 _09809_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _13726_/A _19005_/Q vssd1 vssd1 vccd1 vccd1 _11830_/Y sky130_fd_sc_hd__nand2_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15740__B _15740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _19012_/Q _13257_/A _11760_/Y vssd1 vssd1 vccd1 vccd1 _11761_/X sky130_fd_sc_hd__or3b_1
XFILLER_14_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13500_ _17093_/A vssd1 vssd1 vccd1 vccd1 _17735_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10712_/A vssd1 vssd1 vccd1 vccd1 _10712_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14485_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _18730_/Q vssd1 vssd1 vccd1 vccd1 _14493_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13431_ _19909_/Q _13431_/B vssd1 vssd1 vccd1 vccd1 _13431_/X sky130_fd_sc_hd__and2_1
X_10643_ _10643_/A _10643_/B vssd1 vssd1 vccd1 vccd1 _10643_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16150_ _16474_/B _16150_/B _15735_/A vssd1 vssd1 vccd1 vccd1 _18280_/B sky130_fd_sc_hd__or3b_2
XANTENNA__13782__A1 _13781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13362_ input17/X _13340_/X _13319_/X vssd1 vssd1 vccd1 vccd1 _13362_/X sky130_fd_sc_hd__a21o_1
X_10574_ _19241_/Q _19736_/Q _10574_/S vssd1 vssd1 vccd1 vccd1 _10574_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15101_ _15368_/A vssd1 vssd1 vccd1 vccd1 _15101_/X sky130_fd_sc_hd__clkbuf_2
X_12313_ _12313_/A vssd1 vssd1 vccd1 vccd1 _12313_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11996__A _12583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16081_ _12909_/X _19064_/Q _16089_/S vssd1 vssd1 vccd1 vccd1 _16082_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13293_ _18602_/Q _11683_/X _11733_/X _18634_/Q vssd1 vssd1 vccd1 vccd1 _13293_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15032_ _14881_/X _14884_/X _15032_/S vssd1 vssd1 vccd1 vccd1 _15032_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09466__A _09466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ _12213_/A _14871_/A vssd1 vssd1 vccd1 vccd1 _12244_/X sky130_fd_sc_hd__and2b_1
XFILLER_174_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19840_ _20033_/CLK _19840_/D vssd1 vssd1 vccd1 vccd1 _19840_/Q sky130_fd_sc_hd__dfxtp_1
X_12175_ _12175_/A vssd1 vssd1 vccd1 vccd1 _12260_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11126_ _10996_/X _11125_/X _11140_/A vssd1 vssd1 vccd1 vccd1 _11126_/X sky130_fd_sc_hd__a21o_1
X_19771_ _19771_/CLK _19771_/D vssd1 vssd1 vccd1 vccd1 _19771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16983_ _16983_/A vssd1 vssd1 vccd1 vccd1 _19448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18722_ _18724_/CLK _18722_/D vssd1 vssd1 vccd1 vccd1 _18722_/Q sky130_fd_sc_hd__dfxtp_1
X_11057_ _19525_/Q vssd1 vssd1 vccd1 vccd1 _11058_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15934_ _15936_/A _15934_/B vssd1 vssd1 vccd1 vccd1 _15934_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10008_ _11487_/A vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__clkbuf_2
X_18653_ _18653_/CLK _18653_/D vssd1 vssd1 vccd1 vccd1 _18653_/Q sky130_fd_sc_hd__dfxtp_1
X_15865_ _15881_/A _16839_/B vssd1 vssd1 vccd1 vccd1 _15866_/A sky130_fd_sc_hd__and2_1
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17604_ _17157_/X _19705_/Q _17606_/S vssd1 vssd1 vccd1 vccd1 _17605_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17622__S _17628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14816_ _14927_/A vssd1 vssd1 vccd1 vccd1 _14869_/A sky130_fd_sc_hd__clkbuf_2
X_18584_ _18719_/CLK _18584_/D vssd1 vssd1 vccd1 vccd1 _18584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15796_ _15807_/A _15796_/B vssd1 vssd1 vccd1 vccd1 _15797_/A sky130_fd_sc_hd__or2_1
XFILLER_52_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17535_ _17535_/A vssd1 vssd1 vccd1 vccd1 _19673_/D sky130_fd_sc_hd__clkbuf_1
X_14747_ _18822_/Q _11865_/A _15732_/B _12393_/A _14780_/A vssd1 vssd1 vccd1 vccd1
+ _18822_/D sky130_fd_sc_hd__o221a_1
XFILLER_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11959_ _14931_/A _11959_/B vssd1 vssd1 vccd1 vccd1 _11964_/A sky130_fd_sc_hd__xnor2_2
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13470__B1 _11852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17466_ _17154_/X _19640_/Q _17470_/S vssd1 vssd1 vccd1 vccd1 _17467_/A sky130_fd_sc_hd__mux2_1
X_14678_ _14678_/A vssd1 vssd1 vccd1 vccd1 _18791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19205_ _19764_/CLK _19205_/D vssd1 vssd1 vccd1 vccd1 _19205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16417_ _16417_/A vssd1 vssd1 vccd1 vccd1 _19197_/D sky130_fd_sc_hd__clkbuf_1
X_13629_ _13587_/X _13627_/X _13628_/Y _13590_/X _19009_/Q vssd1 vssd1 vccd1 vccd1
+ _13629_/X sky130_fd_sc_hd__a32o_2
XFILLER_158_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17397_ _17397_/A vssd1 vssd1 vccd1 vccd1 _19609_/D sky130_fd_sc_hd__clkbuf_1
X_19136_ _20015_/CLK _19136_/D vssd1 vssd1 vccd1 vccd1 _19136_/Q sky130_fd_sc_hd__dfxtp_1
X_16348_ _17684_/A vssd1 vssd1 vccd1 vccd1 _16348_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17069__S _17072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16279_ _16279_/A vssd1 vssd1 vccd1 vccd1 _19151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19067_ _19980_/CLK _19067_/D vssd1 vssd1 vccd1 vccd1 _19067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18018_ _19875_/Q _17084_/X _18020_/S vssd1 vssd1 vccd1 vccd1 _18019_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16701__S _16703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19969_ _20034_/CLK _19969_/D vssd1 vssd1 vccd1 vccd1 _19969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09722_ _10954_/S vssd1 vssd1 vccd1 vccd1 _10906_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__11839__A1 _12060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__B _12835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09653_ _09653_/A vssd1 vssd1 vccd1 vccd1 _10449_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_103_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15841__A _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10050__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09584_ _19522_/Q vssd1 vssd1 vccd1 vccd1 _10980_/A sky130_fd_sc_hd__buf_2
XFILLER_43_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16148__S _16148_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10370__S0 _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12016__A1 _18753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13213__B1 _11855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18363__S _18363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09985__S _10254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12567__A2 _12587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10290_ _10290_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _10290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10650__A2_N _09843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16611__S _16613_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14920__A _15103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13980_ _18567_/Q _13982_/C _13979_/Y vssd1 vssd1 vccd1 vccd1 _18567_/D sky130_fd_sc_hd__o21a_1
XFILLER_58_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10189__S0 _10354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ _18715_/Q vssd1 vssd1 vccd1 vccd1 _14450_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11056__A _11131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _12863_/A _12862_/B vssd1 vssd1 vccd1 vccd1 _12862_/Y sky130_fd_sc_hd__nor2_2
X_15650_ _15650_/A vssd1 vssd1 vccd1 vccd1 _18903_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14601_ _14601_/A vssd1 vssd1 vccd1 vccd1 _14615_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_61_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15441__B2 _12574_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11813_ _13656_/A vssd1 vssd1 vccd1 vccd1 _11813_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15470__B _15474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15581_ _13580_/A _18905_/Q _15589_/S vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _18548_/Q _12793_/B vssd1 vssd1 vccd1 vccd1 _12813_/B sky130_fd_sc_hd__nand2_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17151_/X _19575_/Q _17326_/S vssd1 vssd1 vccd1 vccd1 _17321_/A sky130_fd_sc_hd__mux2_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14124_/B _14529_/B _14531_/Y vssd1 vssd1 vccd1 vccd1 _18745_/D sky130_fd_sc_hd__o21a_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _18695_/Q _11698_/Y _11743_/X _11712_/Y vssd1 vssd1 vccd1 vccd1 _11744_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _17251_/A vssd1 vssd1 vccd1 vccd1 _19544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14463_ _14472_/A _14468_/C vssd1 vssd1 vccd1 vccd1 _14463_/Y sky130_fd_sc_hd__nor2_1
X_11675_ _18949_/Q vssd1 vssd1 vccd1 vccd1 _12060_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16202_ _13344_/X _19118_/Q _16206_/S vssd1 vssd1 vccd1 vccd1 _16203_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09959__B1 _09809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13414_ _18481_/Q _12943_/X _12944_/X _18705_/Q _13413_/X vssd1 vssd1 vccd1 vccd1
+ _13414_/X sky130_fd_sc_hd__a221o_1
XANTENNA__14952__A0 _12807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10626_ _10626_/A vssd1 vssd1 vccd1 vccd1 _10626_/X sky130_fd_sc_hd__buf_2
X_17182_ _17182_/A vssd1 vssd1 vccd1 vccd1 _19515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14394_ _18693_/Q _14390_/Y _14393_/Y vssd1 vssd1 vccd1 vccd1 _18693_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10569__A1 _10572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10113__S0 _09595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16133_ _13365_/X _19088_/Q _16133_/S vssd1 vssd1 vccd1 vccd1 _16134_/A sky130_fd_sc_hd__mux2_1
X_13345_ _13344_/X _18446_/Q _13366_/S vssd1 vssd1 vccd1 vccd1 _13346_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10557_ _10557_/A _10557_/B vssd1 vssd1 vccd1 vccd1 _10557_/X sky130_fd_sc_hd__or2_1
XFILLER_143_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16064_ _19059_/Q _16063_/X _16073_/S vssd1 vssd1 vccd1 vccd1 _16065_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13507__B2 _18996_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ _18665_/Q _11815_/X _12890_/X _14501_/A vssd1 vssd1 vccd1 vccd1 _13276_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10488_ _18852_/Q vssd1 vssd1 vccd1 vccd1 _10488_/Y sky130_fd_sc_hd__inv_2
X_15015_ _15013_/X _15014_/X _15113_/S vssd1 vssd1 vccd1 vccd1 _15015_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17617__S _17617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15835__A1_N input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12227_ _12393_/A _12393_/B _12393_/C _12227_/D vssd1 vssd1 vccd1 vccd1 _12227_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__10416__S1 _10320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10135__A _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09924__A _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19823_ _19853_/CLK _19823_/D vssd1 vssd1 vccd1 vccd1 _19823_/Q sky130_fd_sc_hd__dfxtp_1
X_12158_ _18104_/A vssd1 vssd1 vccd1 vccd1 _12557_/A sky130_fd_sc_hd__buf_2
XFILLER_69_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11109_ _09721_/A _11104_/Y _11105_/Y _11108_/X vssd1 vssd1 vccd1 vccd1 _11109_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_111_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19754_ _20013_/CLK _19754_/D vssd1 vssd1 vccd1 vccd1 _19754_/Q sky130_fd_sc_hd__dfxtp_1
X_16966_ _16977_/A vssd1 vssd1 vccd1 vccd1 _16975_/S sky130_fd_sc_hd__buf_6
XANTENNA__16209__A0 _13385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12089_ _11223_/X _18901_/Q _12179_/S vssd1 vssd1 vccd1 vccd1 _14914_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15680__A1 _12554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18705_ _18819_/CLK _18705_/D vssd1 vssd1 vccd1 vccd1 _18705_/Q sky130_fd_sc_hd__dfxtp_1
X_15917_ _15978_/B vssd1 vssd1 vccd1 vccd1 _15928_/A sky130_fd_sc_hd__clkbuf_2
X_19685_ _20039_/CLK _19685_/D vssd1 vssd1 vccd1 vccd1 _19685_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13691__A0 _18477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16897_ _16368_/X _19410_/Q _16903_/S vssd1 vssd1 vccd1 vccd1 _16898_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17352__S _17352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18636_ _18731_/CLK _18636_/D vssd1 vssd1 vccd1 vccd1 _18636_/Q sky130_fd_sc_hd__dfxtp_1
X_15848_ input41/X _15834_/X _15789_/X _15847_/Y vssd1 vssd1 vccd1 vccd1 _17203_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18567_ _19973_/CLK _18567_/D vssd1 vssd1 vccd1 vccd1 _18567_/Q sky130_fd_sc_hd__dfxtp_1
X_15779_ _15779_/A _15783_/B vssd1 vssd1 vccd1 vccd1 _15779_/X sky130_fd_sc_hd__or2_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17518_ _19665_/Q vssd1 vssd1 vccd1 vccd1 _17519_/A sky130_fd_sc_hd__clkbuf_1
X_18498_ _19731_/CLK _18498_/D vssd1 vssd1 vccd1 vccd1 _18498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15196__A0 _18839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17449_ _17449_/A vssd1 vssd1 vccd1 vccd1 _19632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18183__S _18191_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14943__A0 _12713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11757__B1 _14672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19119_ _19936_/CLK _19119_/D vssd1 vssd1 vccd1 vccd1 _19119_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_141_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16431__S _16435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__A _18858_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12260__A _12260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15671__A1 _12446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ _11164_/A vssd1 vssd1 vccd1 vccd1 _11145_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12485__A1 _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12485__B2 _12484_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09350__A1 _09425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _09636_/A vssd1 vssd1 vccd1 vccd1 _09637_/A sky130_fd_sc_hd__buf_2
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_66_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09567_ _09567_/A vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10919__S _10919_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13091__A _13091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _14782_/A _14782_/C vssd1 vssd1 vccd1 vccd1 _09498_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10343__S0 _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14934__A0 _12618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13198__C1 _13289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11460_ _11462_/B _11460_/B vssd1 vssd1 vccd1 vccd1 _11606_/C sky130_fd_sc_hd__nand2_1
XFILLER_109_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10411_ _10411_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10411_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11391_ _19656_/Q _19422_/Q _18487_/Q _19752_/Q _10960_/A _11388_/A vssd1 vssd1 vccd1
+ vccd1 _11391_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10420__B1 _10078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13130_ _13110_/A _13131_/C _18875_/Q vssd1 vssd1 vccd1 vccd1 _13132_/B sky130_fd_sc_hd__a21oi_1
X_10342_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10342_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ _18840_/Q _13560_/B _13215_/S vssd1 vssd1 vccd1 vccd1 _13061_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10273_ _10266_/X _10268_/X _10270_/X _10272_/X _09876_/X vssd1 vssd1 vccd1 vccd1
+ _10273_/X sky130_fd_sc_hd__a221o_2
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12012_ _15633_/B vssd1 vssd1 vccd1 vccd1 _12012_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09744__A _10473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input48_A io_ibus_inst[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11071__S1 _10973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16820_ _16820_/A vssd1 vssd1 vccd1 vccd1 _19376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16751_ _16751_/A vssd1 vssd1 vccd1 vccd1 _19345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13963_ _18561_/Q _13964_/C _18562_/Q vssd1 vssd1 vccd1 vccd1 _13965_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__18268__S _18274_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09877__C1 _09876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15702_ _15702_/A vssd1 vssd1 vccd1 vccd1 _18927_/D sky130_fd_sc_hd__clkbuf_1
X_19470_ _20040_/CLK _19470_/D vssd1 vssd1 vccd1 vccd1 _19470_/Q sky130_fd_sc_hd__dfxtp_1
X_12914_ _18938_/Q vssd1 vssd1 vccd1 vccd1 _16150_/B sky130_fd_sc_hd__buf_4
X_16682_ _16682_/A vssd1 vssd1 vccd1 vccd1 _19315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13894_ _12501_/B _13893_/X _12506_/Y _12509_/X _13890_/X vssd1 vssd1 vccd1 vccd1
+ _18536_/D sky130_fd_sc_hd__o221a_1
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18421_ _18421_/A vssd1 vssd1 vccd1 vccd1 _20039_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15633_ _15633_/A _15633_/B _15633_/C _15633_/D vssd1 vssd1 vccd1 vccd1 _15690_/A
+ sky130_fd_sc_hd__and4_4
X_12845_ _12845_/A vssd1 vssd1 vccd1 vccd1 _12863_/A sky130_fd_sc_hd__buf_12
XANTENNA__12228__A1 _12770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14097__A _14143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17900__S _17904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18352_ _18352_/A _18352_/B _18352_/C vssd1 vssd1 vccd1 vccd1 _18409_/A sky130_fd_sc_hd__or3_4
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _15564_/A vssd1 vssd1 vccd1 vccd1 _18865_/D sky130_fd_sc_hd__clkbuf_1
X_12776_ _18547_/Q _12673_/X _12772_/Y _12775_/Y vssd1 vssd1 vccd1 vccd1 _12776_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10334__S0 _10152_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17303_/A vssd1 vssd1 vccd1 vccd1 _19567_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11727_/A vssd1 vssd1 vccd1 vccd1 _11728_/C sky130_fd_sc_hd__inv_2
X_14515_ _18738_/Q _14512_/B _14514_/Y vssd1 vssd1 vccd1 vccd1 _18738_/D sky130_fd_sc_hd__o21a_1
X_18283_ _17634_/X _19977_/Q _18291_/S vssd1 vssd1 vccd1 vccd1 _18284_/A sky130_fd_sc_hd__mux2_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _15506_/A _15498_/A vssd1 vssd1 vccd1 vccd1 _15495_/X sky130_fd_sc_hd__or2_1
XANTENNA__10885__S1 _10048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13728__A1 _12422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17234_ _17280_/S vssd1 vssd1 vccd1 vccd1 _17243_/S sky130_fd_sc_hd__buf_2
XANTENNA__09919__A _11533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11658_ _11667_/A vssd1 vssd1 vccd1 vccd1 _11660_/A sky130_fd_sc_hd__clkbuf_2
X_14446_ _18714_/Q vssd1 vssd1 vccd1 vccd1 _14450_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11739__B1 _13451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10609_ _19929_/Q _19543_/Q _19993_/Q _19112_/Q _10657_/S _10050_/A vssd1 vssd1 vccd1
+ vccd1 _10610_/B sky130_fd_sc_hd__mux4_1
XFILLER_31_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17165_ _17163_/X _19510_/Q _17177_/S vssd1 vssd1 vccd1 vccd1 _17166_/A sky130_fd_sc_hd__mux2_1
X_14377_ _14377_/A vssd1 vssd1 vccd1 vccd1 _14379_/B sky130_fd_sc_hd__inv_2
XFILLER_156_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11589_ _11589_/A _11626_/A _11589_/C vssd1 vssd1 vccd1 vccd1 _11591_/A sky130_fd_sc_hd__and3_1
X_16116_ _13238_/X _19080_/Q _16122_/S vssd1 vssd1 vccd1 vccd1 _16117_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13328_ _13357_/C _13359_/B _13328_/C vssd1 vssd1 vccd1 vccd1 _13328_/X sky130_fd_sc_hd__and3b_1
XFILLER_155_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17096_ _17203_/A _17096_/B vssd1 vssd1 vccd1 vccd1 _19489_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16047_ _13406_/X _19052_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16048_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13259_ _12956_/A _11760_/Y _13257_/Y _13258_/Y _13307_/A vssd1 vssd1 vccd1 vccd1
+ _13259_/X sky130_fd_sc_hd__a311o_1
XFILLER_130_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09654__A _10449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13361__C1 _13289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19806_ _20030_/CLK _19806_/D vssd1 vssd1 vccd1 vccd1 _19806_/Q sky130_fd_sc_hd__dfxtp_1
X_17998_ _19866_/Q _17055_/X _17998_/S vssd1 vssd1 vccd1 vccd1 _17999_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15653__A1 _12234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19737_ _19995_/CLK _19737_/D vssd1 vssd1 vccd1 vccd1 _19737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16949_ _16339_/X _19433_/Q _16953_/S vssd1 vssd1 vccd1 vccd1 _16950_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18178__S _18180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17082__S _17088_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13904__A _13910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19668_ _19764_/CLK _19668_/D vssd1 vssd1 vccd1 vccd1 _19668_/Q sky130_fd_sc_hd__dfxtp_1
X_09421_ _18826_/Q vssd1 vssd1 vccd1 vccd1 _11716_/A sky130_fd_sc_hd__inv_2
XFILLER_25_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18619_ _18653_/CLK _18619_/D vssd1 vssd1 vccd1 vccd1 _18619_/Q sky130_fd_sc_hd__dfxtp_1
X_19599_ _19853_/CLK _19599_/D vssd1 vssd1 vccd1 vccd1 _19599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09352_ _18830_/Q _14789_/A _18828_/Q vssd1 vssd1 vccd1 vccd1 _09352_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09283_ _09283_/A _09283_/B _09285_/C _09283_/D vssd1 vssd1 vccd1 vccd1 _09284_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10650__B1 _09883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09829__A _11237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13195__A2 _13120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10402__B1 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17257__S _17265_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13785__S _13788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14470__A _14495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09564__A _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10960_ _10960_/A vssd1 vssd1 vccd1 vccd1 _11295_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_141_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10564__S0 _10529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09619_ _11206_/A vssd1 vssd1 vccd1 vccd1 _11140_/A sky130_fd_sc_hd__clkbuf_2
X_10891_ _09546_/A _10880_/X _10889_/X _10078_/A _10890_/Y vssd1 vssd1 vccd1 vccd1
+ _15934_/B sky130_fd_sc_hd__o32a_4
XFILLER_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13025__S _13116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ _12679_/C _12629_/Y _12425_/X vssd1 vssd1 vccd1 vccd1 _12630_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12561_ _12562_/A _12582_/C vssd1 vssd1 vccd1 vccd1 _12561_/X sky130_fd_sc_hd__or2_1
XFILLER_157_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11512_ _11617_/A _11617_/B _11617_/C _11510_/X _11511_/Y vssd1 vssd1 vccd1 vccd1
+ _11616_/B sky130_fd_sc_hd__a41o_1
X_14300_ _18666_/Q _18665_/Q _18664_/Q _14300_/D vssd1 vssd1 vccd1 vccd1 _14312_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__09739__A _10624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15280_ _15115_/X _15119_/X _15280_/S vssd1 vssd1 vccd1 vccd1 _15280_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12492_ _10539_/A _18915_/Q _12687_/A vssd1 vssd1 vccd1 vccd1 _12519_/A sky130_fd_sc_hd__mux2_4
XANTENNA__11988__B _15094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14231_ _14385_/A _14231_/B _14234_/B vssd1 vssd1 vccd1 vccd1 _14232_/A sky130_fd_sc_hd__and3_1
X_11443_ _09828_/A _11442_/X _11401_/A vssd1 vssd1 vccd1 vccd1 _11443_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17956__A _18024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__B hold4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12165__A _12165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14162_ _18625_/Q _14164_/C _14161_/Y vssd1 vssd1 vccd1 vccd1 _18625_/D sky130_fd_sc_hd__o21a_1
X_11374_ _11421_/A _11371_/X _11373_/X vssd1 vssd1 vccd1 vccd1 _11374_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13113_ _13113_/A _13113_/B vssd1 vssd1 vccd1 vccd1 _17023_/A sky130_fd_sc_hd__and2_4
X_10325_ _10194_/A _10310_/X _10324_/X vssd1 vssd1 vccd1 vccd1 _10325_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18970_ _19524_/CLK _18970_/D vssd1 vssd1 vccd1 vccd1 _18970_/Q sky130_fd_sc_hd__dfxtp_2
X_14093_ _14095_/A _14095_/C _14092_/Y vssd1 vssd1 vccd1 vccd1 _18607_/D sky130_fd_sc_hd__o21a_1
XFILLER_98_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14380__A _18690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _17921_/A vssd1 vssd1 vccd1 vccd1 _19831_/D sky130_fd_sc_hd__clkbuf_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13044_/A vssd1 vssd1 vccd1 vccd1 _18430_/D sky130_fd_sc_hd__clkbuf_1
X_10256_ _19678_/Q _19444_/Q _18509_/Q _19774_/Q _09967_/X _09612_/A vssd1 vssd1 vccd1
+ vccd1 _10256_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output154_A _12564_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11509__A _15940_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17852_ _19801_/Q _17052_/X _17854_/S vssd1 vssd1 vccd1 vccd1 _17853_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10187_ _10181_/X _10184_/X _10186_/X _10312_/A _10107_/X vssd1 vssd1 vccd1 vccd1
+ _10194_/B sky130_fd_sc_hd__o221a_1
X_16803_ _16803_/A vssd1 vssd1 vccd1 vccd1 _19368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12449__A1 _18470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17783_ _17783_/A vssd1 vssd1 vccd1 vccd1 _19770_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15923__B _15955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14995_ _15368_/A vssd1 vssd1 vccd1 vccd1 _15286_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19522_ _19523_/CLK _19522_/D vssd1 vssd1 vccd1 vccd1 _19522_/Q sky130_fd_sc_hd__dfxtp_1
X_16734_ _19338_/Q _13816_/X _16736_/S vssd1 vssd1 vccd1 vccd1 _16735_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13946_ _13946_/A _13946_/B _13946_/C vssd1 vssd1 vccd1 vccd1 _18556_/D sky130_fd_sc_hd__nor3_1
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19453_ _19816_/CLK _19453_/D vssd1 vssd1 vccd1 vccd1 _19453_/Q sky130_fd_sc_hd__dfxtp_1
X_16665_ _16676_/A vssd1 vssd1 vccd1 vccd1 _16674_/S sky130_fd_sc_hd__buf_6
X_13877_ _12790_/X _12233_/X _12234_/X _13946_/A vssd1 vssd1 vccd1 vccd1 _18526_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18404_ _18404_/A vssd1 vssd1 vccd1 vccd1 _20031_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17630__S _17632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15616_ _18889_/Q _18921_/Q _15622_/S vssd1 vssd1 vccd1 vccd1 _15617_/A sky130_fd_sc_hd__mux2_1
X_19384_ _19526_/CLK _19384_/D vssd1 vssd1 vccd1 vccd1 _19384_/Q sky130_fd_sc_hd__dfxtp_1
X_12828_ _15899_/A _12828_/B vssd1 vssd1 vccd1 vccd1 _12829_/A sky130_fd_sc_hd__and2_2
X_16596_ _19277_/Q _13826_/X _16602_/S vssd1 vssd1 vccd1 vccd1 _16597_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18335_ _17713_/X _20001_/Q _18335_/S vssd1 vssd1 vccd1 vccd1 _18336_/A sky130_fd_sc_hd__mux2_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _15405_/X _15545_/X _15546_/X _14826_/A _12791_/B vssd1 vssd1 vccd1 vccd1
+ _15547_/X sky130_fd_sc_hd__a32o_2
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14555__A _14672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _15978_/C _18926_/Q _12782_/S vssd1 vssd1 vccd1 vccd1 _12760_/A sky130_fd_sc_hd__mux2_4
XFILLER_91_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09649__A _10872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18266_ _19970_/Q _17716_/A _18274_/S vssd1 vssd1 vccd1 vccd1 _18267_/A sky130_fd_sc_hd__mux2_1
X_15478_ _15478_/A _15478_/B vssd1 vssd1 vccd1 vccd1 _15478_/X sky130_fd_sc_hd__or2_1
X_17217_ _17106_/X _19529_/Q _17221_/S vssd1 vssd1 vccd1 vccd1 _17218_/A sky130_fd_sc_hd__mux2_1
X_14429_ _14433_/C _14431_/C _14428_/Y vssd1 vssd1 vccd1 vccd1 _18703_/D sky130_fd_sc_hd__o21a_1
X_18197_ _18197_/A vssd1 vssd1 vccd1 vccd1 _19939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11188__A1 _11237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_14_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17148_ _17180_/A vssd1 vssd1 vccd1 vccd1 _17161_/S sky130_fd_sc_hd__buf_2
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09970_ _18449_/Q _19478_/Q _19515_/Q _19089_/Q _09657_/A _09637_/A vssd1 vssd1 vccd1
+ vccd1 _09970_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17079_ _19479_/Q _17078_/X _17088_/S vssd1 vssd1 vccd1 vccd1 _17080_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09384__A _18950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11035__S1 _10893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10794__S0 _10787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13101__A2 _13091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17379__A1 _17026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11112__A1 _10854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10469__S _10469_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09404_ _14227_/B _11869_/B vssd1 vssd1 vccd1 vccd1 _09405_/B sky130_fd_sc_hd__nor2_4
XFILLER_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11154__A _11154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ _17098_/B _18981_/Q vssd1 vssd1 vccd1 vccd1 _09698_/B sky130_fd_sc_hd__or2b_1
XFILLER_139_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16156__S _16162_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09266_ _11919_/A _09313_/A vssd1 vssd1 vccd1 vccd1 _09267_/D sky130_fd_sc_hd__nor2_1
XANTENNA__09559__A _09559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_180_clock _18998_/CLK vssd1 vssd1 vccd1 vccd1 _18972_/CLK sky130_fd_sc_hd__clkbuf_16
X_09197_ _11667_/A _09197_/B vssd1 vssd1 vccd1 vccd1 _09198_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12416__C _12416_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10110_ _20036_/Q _19874_/Q _19283_/Q _19053_/Q _10314_/S _10109_/X vssd1 vssd1 vccd1
+ vccd1 _10111_/B sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_195_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _20010_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11090_ _11440_/A vssd1 vssd1 vccd1 vccd1 _11309_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_161_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10041_ _10093_/A _10041_/B vssd1 vssd1 vccd1 vccd1 _10041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11351__A1 _10854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16839__B _16839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13800_ _17036_/A vssd1 vssd1 vccd1 vccd1 _13800_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14780_ _14780_/A _14780_/B vssd1 vssd1 vccd1 vccd1 _14781_/A sky130_fd_sc_hd__and2_1
X_11992_ _11971_/A _12871_/A _11991_/X vssd1 vssd1 vccd1 vccd1 _11993_/B sky130_fd_sc_hd__a21oi_2
XFILLER_57_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10943_ _10952_/A _10943_/B vssd1 vssd1 vccd1 vccd1 _10943_/X sky130_fd_sc_hd__or2_1
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13731_ _19023_/Q _13731_/B vssd1 vssd1 vccd1 vccd1 _13731_/X sky130_fd_sc_hd__or2_1
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_133_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19900_/CLK sky130_fd_sc_hd__clkbuf_16
X_16450_ _16450_/A vssd1 vssd1 vccd1 vccd1 _19212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10874_ _10664_/A _10873_/X _10929_/A vssd1 vssd1 vccd1 vccd1 _10874_/X sky130_fd_sc_hd__a21o_1
X_13662_ _13650_/X _13661_/X _13517_/A vssd1 vssd1 vccd1 vccd1 _13662_/X sky130_fd_sc_hd__a21bo_1
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15401_ _15365_/X _15314_/X _15399_/X _15400_/X vssd1 vssd1 vccd1 vccd1 _15401_/X
+ sky130_fd_sc_hd__a211o_1
X_12613_ _12613_/A _15463_/A vssd1 vssd1 vccd1 vccd1 _12642_/A sky130_fd_sc_hd__xnor2_2
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16381_ _16381_/A vssd1 vssd1 vccd1 vccd1 _16394_/S sky130_fd_sc_hd__buf_4
XANTENNA__16066__S _16066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12603__A1 _18476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13593_ _18875_/Q _13593_/B vssd1 vssd1 vccd1 vccd1 _13594_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18120_ _18120_/A vssd1 vssd1 vccd1 vccd1 _19907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09469__A _18989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15332_ _15247_/X _15044_/X _14986_/X vssd1 vssd1 vccd1 vccd1 _15332_/X sky130_fd_sc_hd__o21a_1
X_12544_ _12544_/A _14860_/A vssd1 vssd1 vccd1 vccd1 _12545_/B sky130_fd_sc_hd__or2_1
XFILLER_157_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_148_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _18653_/CLK sky130_fd_sc_hd__clkbuf_16
X_18051_ _18050_/X _19887_/Q _18061_/S vssd1 vssd1 vccd1 vccd1 _18052_/A sky130_fd_sc_hd__mux2_1
X_12475_ _18524_/Q _18525_/Q _18528_/Q _18529_/Q vssd1 vssd1 vccd1 vccd1 _12476_/D
+ sky130_fd_sc_hd__and4_1
X_15263_ _15152_/X _15262_/X _15348_/S vssd1 vssd1 vccd1 vccd1 _15263_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ _19455_/Q _17001_/X _17008_/S vssd1 vssd1 vccd1 vccd1 _17003_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11426_ _20009_/Q _19847_/Q _19256_/Q _19026_/Q _11124_/A _11073_/A vssd1 vssd1 vccd1
+ vccd1 _11426_/X sky130_fd_sc_hd__mux4_1
X_14214_ _18643_/Q _14210_/B _14213_/Y vssd1 vssd1 vccd1 vccd1 _18643_/D sky130_fd_sc_hd__o21a_1
X_15194_ _15478_/A _15194_/B vssd1 vssd1 vccd1 vccd1 _15194_/X sky130_fd_sc_hd__or2_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_188_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15918__B _15942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14145_ _14156_/D vssd1 vssd1 vccd1 vccd1 _14153_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11357_ _19385_/Q vssd1 vssd1 vccd1 vccd1 _11357_/X sky130_fd_sc_hd__buf_2
XANTENNA__09916__B _12863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12119__A0 _12118_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ _18446_/Q _19475_/Q _19512_/Q _19086_/Q _09655_/A _10185_/X vssd1 vssd1 vccd1
+ vccd1 _10308_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output79_A _12470_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14076_ _14078_/A _14078_/C _14059_/X vssd1 vssd1 vccd1 vccd1 _14076_/Y sky130_fd_sc_hd__a21oi_1
X_18953_ _18956_/CLK _18953_/D vssd1 vssd1 vccd1 vccd1 _18953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11288_ _20012_/Q _19850_/Q _19259_/Q _19029_/Q _11125_/S _11077_/X vssd1 vssd1 vccd1
+ vccd1 _11288_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17904_ _19824_/Q _17023_/X _17904_/S vssd1 vssd1 vccd1 vccd1 _17905_/A sky130_fd_sc_hd__mux2_1
X_13027_ _18871_/Q vssd1 vssd1 vccd1 vccd1 _13046_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10239_ _18859_/Q vssd1 vssd1 vccd1 vccd1 _10239_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13331__A2 _13373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18884_ _19350_/CLK _18884_/D vssd1 vssd1 vccd1 vccd1 _18884_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11342__A1 _11344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17835_ _19793_/Q _17026_/X _17843_/S vssd1 vssd1 vccd1 vccd1 _17836_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17766_ _17766_/A vssd1 vssd1 vccd1 vccd1 _19762_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13095__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14978_ _15068_/A vssd1 vssd1 vccd1 vccd1 _14978_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19505_ _20026_/CLK _19505_/D vssd1 vssd1 vccd1 vccd1 _19505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16717_ _19330_/Q _13790_/X _16725_/S vssd1 vssd1 vccd1 vccd1 _16718_/A sky130_fd_sc_hd__mux2_1
X_13929_ _18551_/Q _18550_/Q _18613_/Q _13929_/D vssd1 vssd1 vccd1 vccd1 _13938_/D
+ sky130_fd_sc_hd__and4_1
X_17697_ _17697_/A vssd1 vssd1 vccd1 vccd1 _17697_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19436_ _19767_/CLK _19436_/D vssd1 vssd1 vccd1 vccd1 _19436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16648_ _16339_/X _19300_/Q _16652_/S vssd1 vssd1 vccd1 vccd1 _16649_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15241__C1 _15951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19367_ _19993_/CLK _19367_/D vssd1 vssd1 vccd1 vccd1 _19367_/Q sky130_fd_sc_hd__dfxtp_1
X_16579_ _16579_/A vssd1 vssd1 vccd1 vccd1 _19269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18318_ _17688_/X _19993_/Q _18324_/S vssd1 vssd1 vccd1 vccd1 _18319_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09379__A _15760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19298_ _19633_/CLK _19298_/D vssd1 vssd1 vccd1 vccd1 _19298_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14347__A1 _14350_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18249_ _18249_/A vssd1 vssd1 vccd1 vccd1 _19962_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18969__CLK _18998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18191__S _18191_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12358__A0 _15940_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10908__A1 _09830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11256__S1 _11208_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09953_ _09833_/X _09950_/X _09952_/X vssd1 vssd1 vccd1 vccd1 _09953_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10053__A _10260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ _09884_/A vssd1 vssd1 vccd1 vccd1 _09884_/X sky130_fd_sc_hd__clkbuf_4
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_11_0_clock clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09842__A _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10988__A _11278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13364__A _17071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_50_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19732_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17221__A0 _17112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18366__S _18374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17270__S _17276_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_65_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _20025_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14195__A _14407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09318_ _14765_/A _14782_/B _11980_/D vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__or3b_1
XFILLER_51_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10590_ _19671_/Q _19437_/Q _18502_/Q _19767_/Q _10657_/S _09607_/A vssd1 vssd1 vccd1
+ vccd1 _10590_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09249_ _09256_/A _09273_/A _09276_/C vssd1 vssd1 vccd1 vccd1 _09290_/A sky130_fd_sc_hd__or3_1
XFILLER_154_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _12260_/A _12658_/A _12260_/C vssd1 vssd1 vccd1 vccd1 _12260_/X sky130_fd_sc_hd__and3_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15738__B _15738_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11211_ _11003_/X _11203_/X _11205_/X _11210_/X _11133_/A vssd1 vssd1 vccd1 vccd1
+ _11211_/X sky130_fd_sc_hd__a221o_1
XFILLER_147_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12191_ _12191_/A _18525_/Q _12477_/C vssd1 vssd1 vccd1 vccd1 _12277_/D sky130_fd_sc_hd__and3_1
XANTENNA__12443__A _12443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11142_ _09560_/A _11135_/X _11137_/X _11141_/X _09873_/A vssd1 vssd1 vccd1 vccd1
+ _11142_/X sky130_fd_sc_hd__a311o_1
XANTENNA__13258__B _18851_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput76 _12390_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[14] sky130_fd_sc_hd__buf_2
XFILLER_122_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput87 _12645_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[24] sky130_fd_sc_hd__buf_2
XFILLER_122_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13313__A2 _13081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11073_ _11073_/A vssd1 vssd1 vccd1 vccd1 _11073_/X sky130_fd_sc_hd__buf_2
X_15950_ _19010_/Q _15927_/X _15928_/X _15949_/Y vssd1 vssd1 vccd1 vccd1 _19010_/D
+ sky130_fd_sc_hd__a22o_1
Xoutput98 _12124_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input30_A io_dbus_rdata[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _10328_/S vssd1 vssd1 vccd1 vccd1 _10037_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14901_ _14901_/A vssd1 vssd1 vccd1 vccd1 _14996_/B sky130_fd_sc_hd__buf_2
X_15881_ _15881_/A _15881_/B vssd1 vssd1 vccd1 vccd1 _15882_/A sky130_fd_sc_hd__and2_1
XANTENNA__11875__A2 _12890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17620_ _17179_/X _19712_/Q _17628_/S vssd1 vssd1 vccd1 vccd1 _17621_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14832_ _14832_/A vssd1 vssd1 vccd1 vccd1 _15201_/B sky130_fd_sc_hd__buf_2
XFILLER_48_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clock _18998_/CLK vssd1 vssd1 vccd1 vccd1 _19324_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17551_ _17551_/A vssd1 vssd1 vccd1 vccd1 _19681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14763_ _14782_/A _15553_/A _14763_/C _14763_/D vssd1 vssd1 vccd1 vccd1 _14764_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18276__S _18278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11975_ _11975_/A _11975_/B _11975_/C _11975_/D vssd1 vssd1 vccd1 vccd1 _12001_/A
+ sky130_fd_sc_hd__nor4_1
XANTENNA_output117_A _12848_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16502_ _19235_/Q _13794_/X _16508_/S vssd1 vssd1 vccd1 vccd1 _16503_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09898__S _09898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13714_ _13714_/A _13714_/B _13714_/C vssd1 vssd1 vccd1 vccd1 _13723_/B sky130_fd_sc_hd__or3_1
X_17482_ _17482_/A vssd1 vssd1 vccd1 vccd1 _19647_/D sky130_fd_sc_hd__clkbuf_1
X_10926_ _19137_/Q _19398_/Q _19297_/Q _19632_/Q _10776_/A _10662_/A vssd1 vssd1 vccd1
+ vccd1 _10927_/B sky130_fd_sc_hd__mux4_1
X_14694_ _18799_/Q _13579_/X _14694_/S vssd1 vssd1 vccd1 vccd1 _14695_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19221_ _19876_/CLK _19221_/D vssd1 vssd1 vccd1 vccd1 _19221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16433_ _19205_/Q _13800_/X _16435_/S vssd1 vssd1 vccd1 vccd1 _16434_/A sky130_fd_sc_hd__mux2_1
X_10857_ _19666_/Q _19432_/Q _18497_/Q _19762_/Q _11488_/S _10856_/X vssd1 vssd1 vccd1
+ vccd1 _10858_/B sky130_fd_sc_hd__mux4_1
X_13645_ _13645_/A vssd1 vssd1 vccd1 vccd1 _18471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12618__A _12618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19152_ _20035_/CLK _19152_/D vssd1 vssd1 vccd1 vccd1 _19152_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _17700_/A vssd1 vssd1 vccd1 vccd1 _16364_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _10793_/A vssd1 vssd1 vccd1 vccd1 _10788_/X sky130_fd_sc_hd__clkbuf_4
X_13576_ _13576_/A vssd1 vssd1 vccd1 vccd1 _18462_/D sky130_fd_sc_hd__clkbuf_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18103_ _18103_/A vssd1 vssd1 vccd1 vccd1 _19902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11260__B1 _11425_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15315_ _15247_/X _15067_/X _14986_/X vssd1 vssd1 vccd1 vccd1 _15315_/X sky130_fd_sc_hd__o21a_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19083_ _20028_/CLK _19083_/D vssd1 vssd1 vccd1 vccd1 _19083_/Q sky130_fd_sc_hd__dfxtp_1
X_12527_ _18473_/Q _12556_/A vssd1 vssd1 vccd1 vccd1 _12527_/X sky130_fd_sc_hd__or2_1
XANTENNA__15929__A _15942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16524__S _16530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16295_ _13501_/X _19159_/Q _16295_/S vssd1 vssd1 vccd1 vccd1 _16296_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18034_ _09425_/B _14562_/X _18050_/S vssd1 vssd1 vccd1 vccd1 _18034_/X sky130_fd_sc_hd__mux2_1
X_15246_ _15244_/Y _15245_/X _15331_/S vssd1 vssd1 vccd1 vccd1 _15246_/X sky130_fd_sc_hd__mux2_1
X_12458_ _12458_/A vssd1 vssd1 vccd1 vccd1 _12458_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11012__B1 _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11409_ _19224_/Q _19719_/Q _11409_/S vssd1 vssd1 vccd1 vccd1 _11409_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15177_ _15178_/B _15177_/B vssd1 vssd1 vccd1 vccd1 _15181_/B sky130_fd_sc_hd__nand2_1
X_12389_ _12389_/A _12389_/B vssd1 vssd1 vccd1 vccd1 _12390_/A sky130_fd_sc_hd__xnor2_4
XFILLER_141_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14128_ _14146_/A _14133_/C vssd1 vssd1 vccd1 vccd1 _14128_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19985_ _19985_/CLK _19985_/D vssd1 vssd1 vccd1 vccd1 _19985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14059_ _14102_/A vssd1 vssd1 vccd1 vccd1 _14059_/X sky130_fd_sc_hd__clkbuf_2
X_18936_ _19524_/CLK _18936_/D vssd1 vssd1 vccd1 vccd1 _18936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09662__A _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18867_ _18867_/CLK _18867_/D vssd1 vssd1 vccd1 vccd1 _18867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17818_ _17818_/A vssd1 vssd1 vccd1 vccd1 _19785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18798_ _19888_/CLK _18798_/D vssd1 vssd1 vccd1 vccd1 _18798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11079__B1 _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17749_ _17649_/X _19755_/Q _17749_/S vssd1 vssd1 vccd1 vccd1 _17750_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15603__S _15611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19419_ _20007_/CLK _19419_/D vssd1 vssd1 vccd1 vccd1 _19419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10841__A3 _10839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10048__A _10048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09837__A _09837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14740__A1 _13742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17265__S _17265_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16493__A1 _13781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09936_ _09929_/X _09931_/X _09933_/X _09935_/X _09876_/X vssd1 vssd1 vccd1 vccd1
+ _09936_/X sky130_fd_sc_hd__a221o_1
XFILLER_104_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11306__A1 _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09867_ _19221_/Q _19812_/Q _19974_/Q _19189_/Q _09598_/X _09851_/A vssd1 vssd1 vccd1
+ vccd1 _09868_/B sky130_fd_sc_hd__mux4_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09798_ _09798_/A vssd1 vssd1 vccd1 vccd1 _09799_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_136_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16609__S _16613_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14918__A _15016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13822__A _17058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _18568_/Q _13054_/B _11759_/X vssd1 vssd1 vccd1 vccd1 _11760_/Y sky130_fd_sc_hd__o21ai_2
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _18438_/Q _19467_/Q _19504_/Q _19078_/Q _10708_/X _10710_/X vssd1 vssd1 vccd1
+ vccd1 _10711_/X sky130_fd_sc_hd__mux4_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10657__S _10657_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ _13082_/A vssd1 vssd1 vccd1 vccd1 _12890_/A sky130_fd_sc_hd__buf_2
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _19671_/Q _19437_/Q _18502_/Q _19767_/Q _09726_/A _10626_/X vssd1 vssd1 vccd1
+ vccd1 _10643_/B sky130_fd_sc_hd__mux4_1
X_13430_ _13188_/A _18861_/Q _12957_/X vssd1 vssd1 vccd1 vccd1 _13430_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_167_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13361_ _13188_/X _11896_/B _13360_/X _13289_/A vssd1 vssd1 vccd1 vccd1 _13361_/X
+ sky130_fd_sc_hd__o211a_1
X_10573_ _19369_/Q _19704_/Q _10573_/S vssd1 vssd1 vccd1 vccd1 _10573_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15100_ _15100_/A _15100_/B vssd1 vssd1 vccd1 vccd1 _15107_/B sky130_fd_sc_hd__nand2_1
X_12312_ _12312_/A _12312_/B vssd1 vssd1 vccd1 vccd1 _12313_/A sky130_fd_sc_hd__and2_4
X_16080_ _16148_/S vssd1 vssd1 vccd1 vccd1 _16089_/S sky130_fd_sc_hd__buf_4
X_13292_ _18810_/Q _13071_/X _12984_/X _12562_/A _13291_/X vssd1 vssd1 vccd1 vccd1
+ _13292_/X sky130_fd_sc_hd__a221o_2
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11488__S _11488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15031_ _15028_/X _15030_/X _15117_/S vssd1 vssd1 vccd1 vccd1 _15031_/X sky130_fd_sc_hd__mux2_1
X_12243_ _12241_/X _12243_/B vssd1 vssd1 vccd1 vccd1 _12246_/A sky130_fd_sc_hd__and2b_2
XFILLER_135_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12174_ _12174_/A vssd1 vssd1 vccd1 vccd1 _12658_/A sky130_fd_sc_hd__buf_2
XFILLER_111_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15484__A _15553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ _19358_/Q _19693_/Q _11125_/S vssd1 vssd1 vccd1 vccd1 _11125_/X sky130_fd_sc_hd__mux2_1
X_19770_ _19996_/CLK _19770_/D vssd1 vssd1 vccd1 vccd1 _19770_/Q sky130_fd_sc_hd__dfxtp_1
X_16982_ _16387_/X _19448_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16983_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13298__A1 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18721_ _18724_/CLK _18721_/D vssd1 vssd1 vccd1 vccd1 _18721_/Q sky130_fd_sc_hd__dfxtp_1
X_15933_ _15053_/X _15928_/A _12239_/Y _15932_/X vssd1 vssd1 vccd1 vccd1 _19003_/D
+ sky130_fd_sc_hd__a31o_1
X_11056_ _11131_/A _11056_/B vssd1 vssd1 vccd1 vccd1 _11056_/X sky130_fd_sc_hd__or2_1
XANTENNA__11848__A2 _12943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10007_ _10007_/A _10007_/B vssd1 vssd1 vccd1 vccd1 _10007_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11517__A _15958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18652_ _18688_/CLK _18652_/D vssd1 vssd1 vccd1 vccd1 _18652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10421__A _15960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15864_ _14749_/B _15856_/X _15788_/X input47/X vssd1 vssd1 vccd1 vccd1 _16839_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17603_ _17603_/A vssd1 vssd1 vccd1 vccd1 _19704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14815_ _14815_/A _14815_/B _14815_/C _14815_/D vssd1 vssd1 vccd1 vccd1 _14927_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_18_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18583_ _18719_/CLK _18583_/D vssd1 vssd1 vccd1 vccd1 _18583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16519__S _16519_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15795_ _15793_/Y _15834_/A _15789_/A _09481_/C vssd1 vssd1 vccd1 vccd1 _15796_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_45_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17534_ _19673_/Q vssd1 vssd1 vccd1 vccd1 _17535_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14746_ _14800_/A vssd1 vssd1 vccd1 vccd1 _14780_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11958_ _11945_/A _11943_/X _11945_/Y _12029_/A vssd1 vssd1 vccd1 vccd1 _11959_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13470__A1 _18676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14547__B _15762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13451__B _13451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17465_ _17465_/A vssd1 vssd1 vccd1 vccd1 _19639_/D sky130_fd_sc_hd__clkbuf_1
X_10909_ _10788_/X _10906_/X _10908_/X vssd1 vssd1 vccd1 vccd1 _10909_/X sky130_fd_sc_hd__a21o_1
XFILLER_149_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14677_ _18791_/Q _14562_/X _14683_/S vssd1 vssd1 vccd1 vccd1 _14678_/A sky130_fd_sc_hd__mux2_1
X_11889_ _12889_/A vssd1 vssd1 vccd1 vccd1 _11889_/X sky130_fd_sc_hd__clkbuf_2
X_19204_ _19957_/CLK _19204_/D vssd1 vssd1 vccd1 vccd1 _19204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16416_ _19197_/Q _13774_/X _16424_/S vssd1 vssd1 vccd1 vccd1 _16417_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13628_ _13709_/A _19009_/Q vssd1 vssd1 vccd1 vccd1 _13628_/Y sky130_fd_sc_hd__nand2_1
X_17396_ _19609_/Q _17052_/X _17398_/S vssd1 vssd1 vccd1 vccd1 _17397_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19135_ _19726_/CLK _19135_/D vssd1 vssd1 vccd1 vccd1 _19135_/Q sky130_fd_sc_hd__dfxtp_1
X_16347_ _16347_/A vssd1 vssd1 vccd1 vccd1 _19174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16254__S _16258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13559_ _13559_/A vssd1 vssd1 vccd1 vccd1 _18460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14563__A _14601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09657__A _09657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19066_ _19979_/CLK _19066_/D vssd1 vssd1 vccd1 vccd1 _19066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16278_ _13354_/X _19151_/Q _16280_/S vssd1 vssd1 vccd1 vccd1 _16279_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18017_ _18017_/A vssd1 vssd1 vccd1 vccd1 _19874_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13179__A _17036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15229_ _14858_/X _15203_/X _15074_/X vssd1 vssd1 vccd1 vccd1 _15229_/X sky130_fd_sc_hd__o21a_1
XFILLER_172_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12514__C _15397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17085__S _17088_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19968_ _20030_/CLK _19968_/D vssd1 vssd1 vccd1 vccd1 _19968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09721_ _09721_/A vssd1 vssd1 vccd1 vccd1 _10954_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18919_ _18924_/CLK _18919_/D vssd1 vssd1 vccd1 vccd1 _18919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19899_ _19899_/CLK _19899_/D vssd1 vssd1 vccd1 vccd1 _19899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17813__S _17821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _09652_/A vssd1 vssd1 vccd1 vccd1 _09653_/A sky130_fd_sc_hd__buf_4
XFILLER_94_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09583_ _09929_/A vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__buf_2
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16429__S _16435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13461__A1 _12967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10370__S1 _10054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13788__S _13788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15569__A _15602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17784__A _17795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15910__A0 _12032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09919_ _11533_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09919_/X sky130_fd_sc_hd__and2_1
XFILLER_59_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10189__S1 _10185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20039_ _20039_/CLK _20039_/D vssd1 vssd1 vccd1 vccd1 _20039_/Q sky130_fd_sc_hd__dfxtp_1
X_12930_ _14026_/B _11732_/X _11733_/X _18615_/Q vssd1 vssd1 vccd1 vccd1 _12930_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10241__A _15972_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12861_/A vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14648__A _14648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14600_/A vssd1 vssd1 vccd1 vccd1 _18768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _12188_/A _11812_/B vssd1 vssd1 vccd1 vccd1 _11860_/C sky130_fd_sc_hd__nand2_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _15602_/A vssd1 vssd1 vccd1 vccd1 _15589_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12792_ _18548_/Q _12793_/B vssd1 vssd1 vccd1 vccd1 _12792_/X sky130_fd_sc_hd__or2_1
XFILLER_57_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13452__A1 _18483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14531_ _14124_/B _14529_/B _14507_/X vssd1 vssd1 vccd1 vccd1 _14531_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11743_/A _11743_/B _11743_/C vssd1 vssd1 vccd1 vccd1 _11743_/X sky130_fd_sc_hd__or3_1
XFILLER_15_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _17154_/X _19544_/Q _17254_/S vssd1 vssd1 vccd1 vccd1 _17251_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14462_ _14462_/A vssd1 vssd1 vccd1 vccd1 _14468_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _15719_/A _13510_/B vssd1 vssd1 vccd1 vccd1 _14672_/B sky130_fd_sc_hd__nor2_2
XFILLER_14_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16201_ _16201_/A vssd1 vssd1 vccd1 vccd1 _19117_/D sky130_fd_sc_hd__clkbuf_1
X_13413_ _19908_/Q _13431_/B vssd1 vssd1 vccd1 vccd1 _13413_/X sky130_fd_sc_hd__and2_1
XFILLER_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ _10625_/A vssd1 vssd1 vccd1 vccd1 _10626_/A sky130_fd_sc_hd__buf_2
X_17181_ _17179_/X _19515_/Q _17193_/S vssd1 vssd1 vccd1 vccd1 _17182_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14952__A1 _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14393_ _14413_/A _14398_/C vssd1 vssd1 vccd1 vccd1 _14393_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11310__S0 _11230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16132_ _16132_/A vssd1 vssd1 vccd1 vccd1 _19087_/D sky130_fd_sc_hd__clkbuf_1
X_13344_ _17707_/A vssd1 vssd1 vccd1 vccd1 _13344_/X sky130_fd_sc_hd__clkbuf_1
X_10556_ _19209_/Q _19800_/Q _19962_/Q _19177_/Q _10319_/A _10497_/X vssd1 vssd1 vccd1
+ vccd1 _10557_/B sky130_fd_sc_hd__mux4_1
XFILLER_128_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12615__B _12641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16063_ _12188_/X _14554_/X _12071_/B vssd1 vssd1 vccd1 vccd1 _16063_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16802__S _16808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10487_ _10480_/Y _10482_/Y _10484_/Y _10486_/Y _09821_/A vssd1 vssd1 vccd1 vccd1
+ _10487_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13275_ _18733_/Q vssd1 vssd1 vccd1 vccd1 _14501_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_154_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15014_ _14956_/X _14943_/X _15014_/S vssd1 vssd1 vccd1 vccd1 _15014_/X sky130_fd_sc_hd__mux2_1
X_12226_ _12249_/B _12226_/B vssd1 vssd1 vccd1 vccd1 _12227_/D sky130_fd_sc_hd__nand2_1
XFILLER_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12157_ _13511_/B vssd1 vssd1 vccd1 vccd1 _18104_/A sky130_fd_sc_hd__clkbuf_4
X_19822_ _19951_/CLK _19822_/D vssd1 vssd1 vccd1 vccd1 _19822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11108_ _11108_/A vssd1 vssd1 vccd1 vccd1 _11108_/X sky130_fd_sc_hd__clkbuf_4
X_16965_ _16965_/A vssd1 vssd1 vccd1 vccd1 _19440_/D sky130_fd_sc_hd__clkbuf_1
X_19753_ _20012_/CLK _19753_/D vssd1 vssd1 vccd1 vccd1 _19753_/Q sky130_fd_sc_hd__dfxtp_1
X_12088_ _12088_/A _15183_/A vssd1 vssd1 vccd1 vccd1 _12091_/A sky130_fd_sc_hd__xnor2_1
XFILLER_77_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15942__A _15942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ _11032_/Y _11034_/Y _11036_/Y _11038_/Y _11166_/A vssd1 vssd1 vccd1 vccd1
+ _11039_/X sky130_fd_sc_hd__o221a_1
X_15916_ _15916_/A vssd1 vssd1 vccd1 vccd1 _15978_/B sky130_fd_sc_hd__clkbuf_4
X_18704_ _18744_/CLK _18704_/D vssd1 vssd1 vccd1 vccd1 _18704_/Q sky130_fd_sc_hd__dfxtp_1
X_19684_ _19810_/CLK _19684_/D vssd1 vssd1 vccd1 vccd1 _19684_/Q sky130_fd_sc_hd__dfxtp_1
X_16896_ _16896_/A vssd1 vssd1 vccd1 vccd1 _19409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09940__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18635_ _19683_/CLK _18635_/D vssd1 vssd1 vccd1 vccd1 _18635_/Q sky130_fd_sc_hd__dfxtp_1
X_15847_ _15847_/A vssd1 vssd1 vccd1 vccd1 _15847_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14558__A _15833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11129__S0 _11258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18566_ _20005_/CLK _18566_/D vssd1 vssd1 vccd1 vccd1 _18566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _09471_/C _11867_/X _15777_/X _15769_/X vssd1 vssd1 vccd1 vccd1 _18957_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17517_ _17517_/A vssd1 vssd1 vccd1 vccd1 _19664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11454__B1 _11292_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14729_ _14729_/A vssd1 vssd1 vccd1 vccd1 _14738_/S sky130_fd_sc_hd__buf_2
X_18497_ _19861_/CLK _18497_/D vssd1 vssd1 vccd1 vccd1 _18497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17448_ _17128_/X _19632_/Q _17448_/S vssd1 vssd1 vccd1 vccd1 _17449_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14943__A1 _15138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17379_ _19601_/Q _17026_/X _17387_/S vssd1 vssd1 vccd1 vccd1 _17380_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12806__A _15553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14293__A _14479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__A1 _18472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11301__S0 _11230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19118_ _19644_/CLK _19118_/D vssd1 vssd1 vccd1 vccd1 _19118_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12954__B1 _12890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19049_ _19936_/CLK _19049_/D vssd1 vssd1 vccd1 vccd1 _19049_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17808__S _17808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16712__S _16714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09704_ _11435_/A vssd1 vssd1 vccd1 vccd1 _11164_/A sky130_fd_sc_hd__buf_2
XANTENNA__11157__A _11157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11142__C1 _09873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10496__B2 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _09668_/S vssd1 vssd1 vccd1 vccd1 _09635_/X sky130_fd_sc_hd__buf_4
XANTENNA__09350__A2 _09347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11693__B1 _12890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09566_ _09566_/A vssd1 vssd1 vccd1 vccd1 _09567_/A sky130_fd_sc_hd__buf_2
XFILLER_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15998__S _15998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18374__S _18374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09497_ _12536_/A _11912_/A vssd1 vssd1 vccd1 vccd1 _14782_/C sky130_fd_sc_hd__nand2_1
XFILLER_24_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10343__S1 _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14934__A1 _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ _19933_/Q _19547_/Q _19997_/Q _19116_/Q _09995_/A _10400_/A vssd1 vssd1 vccd1
+ vccd1 _10411_/B sky130_fd_sc_hd__mux4_1
XANTENNA__16136__A0 _13385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _09828_/A _11389_/X _11404_/A vssd1 vssd1 vccd1 vccd1 _11390_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10341_ _19214_/Q _19805_/Q _19967_/Q _19182_/Q _10166_/S _10223_/X vssd1 vssd1 vccd1
+ vccd1 _10342_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17718__S _17730_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10420__A1 _09547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16622__S _16630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14931__A _14931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13060_ _18653_/Q _11889_/X _13055_/X _13059_/X vssd1 vssd1 vccd1 vccd1 _13560_/B
+ sky130_fd_sc_hd__a211o_2
X_10272_ _10064_/X _10271_/X _09980_/X vssd1 vssd1 vccd1 vccd1 _10272_/X sky130_fd_sc_hd__o21a_1
XFILLER_155_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12011_ _12448_/S _11994_/A _12008_/X _12010_/X vssd1 vssd1 vccd1 vccd1 _12011_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12451__A _12452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17453__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16750_ _19345_/Q _13838_/X _16758_/S vssd1 vssd1 vccd1 vccd1 _16751_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15762__A _15762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13962_ _18561_/Q _13964_/C _13961_/Y vssd1 vssd1 vccd1 vccd1 _18561_/D sky130_fd_sc_hd__o21a_1
XANTENNA__14870__A0 _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15701_ _18927_/Q _18548_/Q _15703_/S vssd1 vssd1 vccd1 vccd1 _15702_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10031__S0 _10275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ _12913_/A vssd1 vssd1 vccd1 vccd1 _16691_/B sky130_fd_sc_hd__buf_4
X_16681_ _16387_/X _19315_/Q _16685_/S vssd1 vssd1 vccd1 vccd1 _16682_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09972__S0 _09967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13893_ _13900_/A vssd1 vssd1 vccd1 vccd1 _13893_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13282__A _17055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18420_ _17732_/X _20039_/Q _18422_/S vssd1 vssd1 vccd1 vccd1 _18421_/A sky130_fd_sc_hd__mux2_1
X_15632_ _15632_/A vssd1 vssd1 vccd1 vccd1 _18896_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12844_ _12844_/A _12844_/B vssd1 vssd1 vccd1 vccd1 _12844_/Y sky130_fd_sc_hd__nor2_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14622__A0 _12508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _18351_/A vssd1 vssd1 vccd1 vccd1 _20008_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _18865_/Q _18897_/Q _15567_/S vssd1 vssd1 vccd1 vccd1 _15564_/A sky130_fd_sc_hd__mux2_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12480_/X _12773_/Y _12799_/B _12583_/X vssd1 vssd1 vccd1 vccd1 _12775_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10334__S1 _10153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__S0 _11532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17302_ _17125_/X _19567_/Q _17304_/S vssd1 vssd1 vccd1 vccd1 _17303_/A sky130_fd_sc_hd__mux2_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15701__S _15703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16375__A0 _16374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14514_/A _14518_/C vssd1 vssd1 vccd1 vccd1 _14514_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11726_ _14159_/A vssd1 vssd1 vccd1 vccd1 _15715_/B sky130_fd_sc_hd__buf_4
XFILLER_30_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18282_ _18350_/S vssd1 vssd1 vccd1 vccd1 _18291_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15498_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _15494_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17233_ _17233_/A vssd1 vssd1 vccd1 vccd1 _19536_/D sky130_fd_sc_hd__clkbuf_1
X_14445_ _14445_/A _14445_/B vssd1 vssd1 vccd1 vccd1 _18709_/D sky130_fd_sc_hd__nor2_1
XANTENNA__13728__A2 _13727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ _11657_/A _11657_/B vssd1 vssd1 vccd1 vccd1 _11657_/Y sky130_fd_sc_hd__nor2_4
XFILLER_30_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11739__A1 _18753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12626__A _18477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10608_ _10836_/A _10608_/B vssd1 vssd1 vccd1 vccd1 _10608_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10098__S0 _10094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17164_ _17180_/A vssd1 vssd1 vccd1 vccd1 _17177_/S sky130_fd_sc_hd__buf_4
XFILLER_156_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14376_ _14378_/B _14381_/D _18689_/Q vssd1 vssd1 vccd1 vccd1 _14377_/A sky130_fd_sc_hd__a21o_1
X_11588_ _11588_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16115_ _16115_/A vssd1 vssd1 vccd1 vccd1 _19079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17628__S _17628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13327_ _13664_/A _13306_/X _13288_/B _18887_/Q vssd1 vssd1 vccd1 vccd1 _13328_/C
+ sky130_fd_sc_hd__a31o_1
X_17095_ _17095_/A vssd1 vssd1 vccd1 vccd1 _19484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10539_ _10539_/A _12849_/B vssd1 vssd1 vccd1 vccd1 _10540_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16046_ _16046_/A vssd1 vssd1 vccd1 vccd1 _19051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13258_ _13473_/A _18851_/Q vssd1 vssd1 vccd1 vccd1 _13258_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14560__B _18995_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12209_ _12209_/A _12209_/B _12209_/C _15219_/A vssd1 vssd1 vccd1 vccd1 _12323_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA__10175__B1 _09843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13189_ _13189_/A vssd1 vssd1 vccd1 vccd1 _13189_/X sky130_fd_sc_hd__buf_2
XFILLER_69_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19805_ _19999_/CLK _19805_/D vssd1 vssd1 vccd1 vccd1 _19805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17997_ _17997_/A vssd1 vssd1 vccd1 vccd1 _19865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17363__S _17365_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19736_ _19994_/CLK _19736_/D vssd1 vssd1 vccd1 vccd1 _19736_/Q sky130_fd_sc_hd__dfxtp_1
X_16948_ _16948_/A vssd1 vssd1 vccd1 vccd1 _19432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10478__A1 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09670__A _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16879_ _16342_/X _19402_/Q _16881_/S vssd1 vssd1 vccd1 vccd1 _16880_/A sky130_fd_sc_hd__mux2_1
X_19667_ _19796_/CLK _19667_/D vssd1 vssd1 vccd1 vccd1 _19667_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_10_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09420_ _18960_/Q _18959_/Q _11772_/B vssd1 vssd1 vccd1 vccd1 _09420_/X sky130_fd_sc_hd__and3_1
X_18618_ _18653_/CLK _18618_/D vssd1 vssd1 vccd1 vccd1 _18618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19598_ _19951_/CLK _19598_/D vssd1 vssd1 vccd1 vccd1 _19598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ _18829_/Q vssd1 vssd1 vccd1 vccd1 _14789_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18194__S _18202_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18549_ _18773_/CLK _18549_/D vssd1 vssd1 vccd1 vccd1 _18549_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15611__S _15611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09282_ _11664_/A _09282_/B _09282_/C _09282_/D vssd1 vssd1 vccd1 vccd1 _09491_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_100_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15708__A3 _13700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12927__B1 _12881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10402__A1 _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15847__A _15847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16442__S _16446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09845__A _15980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18043__A0 _18837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09580__A _10200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11666__B1 _11657_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__S1 _10011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09618_ _11068_/A vssd1 vssd1 vccd1 vccd1 _11206_/A sky130_fd_sc_hd__buf_2
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ _18843_/Q vssd1 vssd1 vccd1 vccd1 _10890_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09549_ _09549_/A vssd1 vssd1 vccd1 vccd1 _09550_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16617__S _16617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12560_ _18777_/Q vssd1 vssd1 vccd1 vccd1 _12562_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10641__A1 _10690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _11510_/B _10818_/A _11508_/Y vssd1 vssd1 vccd1 vccd1 _11511_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12491_ _12517_/S vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12446__A _12446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14230_ _18646_/Q _14242_/C vssd1 vssd1 vccd1 vccd1 _14234_/B sky130_fd_sc_hd__nand2_1
XFILLER_109_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11442_ _19224_/Q _19719_/Q _11442_/S vssd1 vssd1 vccd1 vccd1 _11442_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09458__C _18970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11373_ _11206_/A _11372_/X _09681_/A vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__o21a_1
X_14161_ _18625_/Q _14164_/C _14160_/X vssd1 vssd1 vccd1 vccd1 _14161_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10324_ _10192_/X _10312_/Y _10316_/Y _10323_/Y _09876_/A vssd1 vssd1 vccd1 vccd1
+ _10324_/X sky130_fd_sc_hd__o311a_1
XANTENNA_input60_A io_ibus_inst[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ _13350_/S _13108_/X _13110_/Y _13111_/X _13297_/A vssd1 vssd1 vccd1 vccd1
+ _13113_/B sky130_fd_sc_hd__a221o_1
XANTENNA__09755__A _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14092_ _14095_/A _14095_/C _14059_/X vssd1 vssd1 vccd1 vccd1 _14092_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10255_ _09597_/A _10253_/Y _10254_/Y _10054_/X vssd1 vssd1 vccd1 vccd1 _10255_/X
+ sky130_fd_sc_hd__a211o_1
X_17920_ _19831_/Q _17046_/X _17926_/S vssd1 vssd1 vccd1 vccd1 _17921_/A sky130_fd_sc_hd__mux2_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _13042_/X _18430_/Q _13116_/S vssd1 vssd1 vccd1 vccd1 _13044_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13894__A1 _12501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17851_ _17851_/A vssd1 vssd1 vccd1 vccd1 _19800_/D sky130_fd_sc_hd__clkbuf_1
X_10186_ _19681_/Q _19447_/Q _18512_/Q _19777_/Q _09655_/A _10185_/X vssd1 vssd1 vccd1
+ vccd1 _10186_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11509__B _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output147_A _12403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16802_ _16352_/X _19368_/Q _16808_/S vssd1 vssd1 vccd1 vccd1 _16803_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17782_ _17697_/X _19770_/Q _17782_/S vssd1 vssd1 vccd1 vccd1 _17783_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15923__C _15923_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14994_ _15102_/A vssd1 vssd1 vccd1 vccd1 _14994_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18034__A0 _09425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16733_ _16733_/A vssd1 vssd1 vccd1 vccd1 _19337_/D sky130_fd_sc_hd__clkbuf_1
X_19521_ _19846_/CLK _19521_/D vssd1 vssd1 vccd1 vccd1 _19521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _18556_/Q _13945_/B _13945_/C vssd1 vssd1 vccd1 vccd1 _13946_/C sky130_fd_sc_hd__and3_1
XFILLER_47_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17911__S _17915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19452_ _20040_/CLK _19452_/D vssd1 vssd1 vccd1 vccd1 _19452_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11525__A _15976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16664_ _16664_/A vssd1 vssd1 vccd1 vccd1 _19307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13876_ _15715_/B vssd1 vssd1 vccd1 vccd1 _13946_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_34_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18403_ _17707_/X _20031_/Q _18407_/S vssd1 vssd1 vccd1 vccd1 _18404_/A sky130_fd_sc_hd__mux2_1
X_15615_ _15615_/A vssd1 vssd1 vccd1 vccd1 _18888_/D sky130_fd_sc_hd__clkbuf_1
X_19383_ _20040_/CLK _19383_/D vssd1 vssd1 vccd1 vccd1 _19383_/Q sky130_fd_sc_hd__dfxtp_1
X_12827_ _12827_/A _12827_/B vssd1 vssd1 vccd1 vccd1 _12827_/Y sky130_fd_sc_hd__nor2_4
X_16595_ _16595_/A vssd1 vssd1 vccd1 vccd1 _19276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18334_ _18334_/A vssd1 vssd1 vccd1 vccd1 _20000_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17212__A _17280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15546_ _15546_/A _15546_/B vssd1 vssd1 vccd1 vccd1 _15546_/X sky130_fd_sc_hd__or2_1
X_12758_ _15531_/A _12758_/B vssd1 vssd1 vccd1 vccd1 _12762_/A sky130_fd_sc_hd__xor2_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14555__B _14555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18265_ _18265_/A vssd1 vssd1 vccd1 vccd1 _18274_/S sky130_fd_sc_hd__buf_4
X_11709_ _18754_/Q _11670_/A _13164_/B _19897_/Q vssd1 vssd1 vccd1 vccd1 _11709_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15477_ _15151_/X _15204_/X _15476_/X _15413_/X vssd1 vssd1 vccd1 vccd1 _15477_/X
+ sky130_fd_sc_hd__a211o_1
X_12689_ _12689_/A _12715_/A vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__xor2_4
XFILLER_129_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17216_ _17216_/A vssd1 vssd1 vccd1 vccd1 _19528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14428_ _14433_/C _14431_/C _14427_/X vssd1 vssd1 vccd1 vccd1 _14428_/Y sky130_fd_sc_hd__a21oi_1
X_18196_ _17720_/X _19939_/Q _18202_/S vssd1 vssd1 vccd1 vccd1 _18197_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17147_ _17684_/A vssd1 vssd1 vccd1 vccd1 _17147_/X sky130_fd_sc_hd__buf_2
XFILLER_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14359_ _14407_/A vssd1 vssd1 vccd1 vccd1 _14399_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10396__B1 _09843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14571__A _15833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09665__A _10822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17078_ _17078_/A vssd1 vssd1 vccd1 vccd1 _17078_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12137__A1 _12165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16029_ _13263_/X _19044_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16030_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13187__A _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18189__S _18191_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19719_ _19720_/CLK _19719_/D vssd1 vssd1 vccd1 vccd1 _19719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17821__S _17821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09403_ _09403_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _09405_/A sky130_fd_sc_hd__nor2_2
XFILLER_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13650__A _13650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _18981_/Q _17098_/B vssd1 vssd1 vccd1 vccd1 _09698_/A sky130_fd_sc_hd__or2b_1
XFILLER_166_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09265_ _11932_/A _11932_/B _09265_/C _09265_/D vssd1 vssd1 vccd1 vccd1 _09292_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12266__A _15934_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09196_ _09521_/A _11950_/A vssd1 vssd1 vccd1 vccd1 _09197_/B sky130_fd_sc_hd__nor2_1
XFILLER_135_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12376__A1 _13650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17268__S _17276_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12713__B _12713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13097__A _17020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10139__B1 _09547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10514__A _15956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _19153_/Q _19414_/Q _19313_/Q _19648_/Q _10095_/S _10028_/X vssd1 vssd1 vccd1
+ vccd1 _10041_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10234__S0 _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_88_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11991_ _11964_/A _14901_/A vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__and2b_1
XFILLER_75_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _13737_/A _13737_/C vssd1 vssd1 vccd1 vccd1 _13730_/Y sky130_fd_sc_hd__xnor2_1
X_10942_ _19922_/Q _19536_/Q _19986_/Q _19105_/Q _10907_/S _10624_/A vssd1 vssd1 vccd1
+ vccd1 _10943_/B sky130_fd_sc_hd__mux4_1
XFILLER_44_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13661_ _13656_/X _13657_/X _13659_/Y _13660_/X _19013_/Q vssd1 vssd1 vccd1 vccd1
+ _13661_/X sky130_fd_sc_hd__a32o_2
X_10873_ _19362_/Q _19697_/Q _10921_/S vssd1 vssd1 vccd1 vccd1 _10873_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15400_ _15400_/A vssd1 vssd1 vccd1 vccd1 _15400_/X sky130_fd_sc_hd__clkbuf_2
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12612_/A vssd1 vssd1 vccd1 vccd1 _15463_/A sky130_fd_sc_hd__clkbuf_2
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _17716_/A vssd1 vssd1 vccd1 vccd1 _16380_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _18875_/Q _13593_/B vssd1 vssd1 vccd1 vccd1 _13603_/C sky130_fd_sc_hd__or2_2
XFILLER_40_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15331_ _14985_/X _15330_/X _15331_/S vssd1 vssd1 vccd1 vccd1 _15331_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10614__B2 _10668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17967__A _18024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12543_ _12544_/A _14860_/A vssd1 vssd1 vccd1 vccd1 _12545_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18050_ _18839_/Q _13553_/X _18050_/S vssd1 vssd1 vccd1 vccd1 _18050_/X sky130_fd_sc_hd__mux2_1
X_15262_ _15059_/X _15064_/X _15298_/S vssd1 vssd1 vccd1 vccd1 _15262_/X sky130_fd_sc_hd__mux2_1
X_12474_ _18526_/Q _18527_/Q _18530_/Q _18533_/Q vssd1 vssd1 vccd1 vccd1 _12476_/C
+ sky130_fd_sc_hd__and4_1
X_17001_ _17001_/A vssd1 vssd1 vccd1 vccd1 _17001_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14213_ _14239_/A _14215_/B vssd1 vssd1 vccd1 vccd1 _14213_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ _11425_/A _11425_/B vssd1 vssd1 vccd1 vccd1 _11425_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15487__A _15487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15193_ _15190_/X _15192_/X _15247_/A vssd1 vssd1 vccd1 vccd1 _15194_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10378__B1 _10162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14144_ _18621_/Q _18620_/Q _18619_/Q _14144_/D vssd1 vssd1 vccd1 vccd1 _14156_/D
+ sky130_fd_sc_hd__and4_1
X_11356_ _19384_/Q vssd1 vssd1 vccd1 vccd1 _11356_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13316__A0 _18854_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ _10312_/A _10307_/B vssd1 vssd1 vccd1 vccd1 _10307_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14075_ _18600_/Q _14072_/B _14074_/Y vssd1 vssd1 vccd1 vccd1 _18600_/D sky130_fd_sc_hd__o21a_1
X_18952_ _18956_/CLK _18952_/D vssd1 vssd1 vccd1 vccd1 _18952_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10424__A _10424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11287_ _11287_/A _11287_/B vssd1 vssd1 vccd1 vccd1 _11287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13026_ _13026_/A vssd1 vssd1 vccd1 vccd1 _18429_/D sky130_fd_sc_hd__clkbuf_1
X_17903_ _17903_/A vssd1 vssd1 vccd1 vccd1 _19823_/D sky130_fd_sc_hd__clkbuf_1
X_10238_ _10231_/Y _10233_/Y _10235_/Y _10237_/Y _09822_/A vssd1 vssd1 vccd1 vccd1
+ _10238_/X sky130_fd_sc_hd__o221a_1
XANTENNA__15934__B _15934_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18883_ _18918_/CLK _18883_/D vssd1 vssd1 vccd1 vccd1 _18883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10169_ _10082_/A _10166_/X _10168_/X vssd1 vssd1 vccd1 vccd1 _10169_/X sky130_fd_sc_hd__a21o_1
X_17834_ _17880_/S vssd1 vssd1 vccd1 vccd1 _17843_/S sky130_fd_sc_hd__buf_4
XFILLER_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17765_ _17672_/X _19762_/Q _17771_/S vssd1 vssd1 vccd1 vccd1 _17766_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14977_ _15151_/A vssd1 vssd1 vccd1 vccd1 _14977_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19504_ _19990_/CLK _19504_/D vssd1 vssd1 vccd1 vccd1 _19504_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17641__S _17650_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16716_ _16762_/S vssd1 vssd1 vccd1 vccd1 _16725_/S sky130_fd_sc_hd__clkbuf_4
X_13928_ _14507_/A vssd1 vssd1 vccd1 vccd1 _13967_/A sky130_fd_sc_hd__buf_2
XFILLER_81_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17696_ _17696_/A vssd1 vssd1 vccd1 vccd1 _19737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19435_ _20023_/CLK _19435_/D vssd1 vssd1 vccd1 vccd1 _19435_/Q sky130_fd_sc_hd__dfxtp_1
X_16647_ _16647_/A vssd1 vssd1 vccd1 vccd1 _19299_/D sky130_fd_sc_hd__clkbuf_1
X_13859_ _13859_/A vssd1 vssd1 vccd1 vccd1 _18517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19366_ _19959_/CLK _19366_/D vssd1 vssd1 vccd1 vccd1 _19366_/Q sky130_fd_sc_hd__dfxtp_1
X_16578_ _19269_/Q _13800_/X _16580_/S vssd1 vssd1 vccd1 vccd1 _16579_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18317_ _18317_/A vssd1 vssd1 vccd1 vccd1 _19992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15529_ _15211_/X _15531_/B _15081_/X _15528_/X vssd1 vssd1 vccd1 vccd1 _15529_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19297_ _19985_/CLK _19297_/D vssd1 vssd1 vccd1 vccd1 _19297_/Q sky130_fd_sc_hd__dfxtp_1
X_18248_ _19962_/Q _17691_/A _18252_/S vssd1 vssd1 vccd1 vccd1 _18249_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17088__S _17088_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15397__A _15397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18179_ _18179_/A vssd1 vssd1 vccd1 vccd1 _19931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09395__A _11777_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09952_ _09824_/A _09951_/X _09765_/A vssd1 vssd1 vccd1 vccd1 _09952_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13858__A1 _13857_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09883_ _09883_/A vssd1 vssd1 vccd1 vccd1 _09884_/A sky130_fd_sc_hd__clkbuf_4
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15480__A0 _18857_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16167__S _16173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09317_ _11950_/A _09500_/B vssd1 vssd1 vccd1 vccd1 _11980_/D sky130_fd_sc_hd__or2_1
XANTENNA__09289__B _09289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16691__A _16691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _09316_/B vssd1 vssd1 vccd1 vccd1 _09248_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_132_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ _09230_/A _09283_/A vssd1 vssd1 vccd1 vccd1 _09311_/A sky130_fd_sc_hd__or2_1
XFILLER_135_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11210_ _11287_/A _11209_/X _11058_/X vssd1 vssd1 vccd1 vccd1 _11210_/X sky130_fd_sc_hd__o21a_1
XFILLER_134_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12190_ _12191_/A _12477_/C _18525_/Q vssd1 vssd1 vccd1 vccd1 _12192_/A sky130_fd_sc_hd__a21oi_1
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11141_ _11001_/A _11138_/X _11140_/X _09683_/A vssd1 vssd1 vccd1 vccd1 _11141_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16630__S _16630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11072_ _11070_/X _11071_/X _11003_/A vssd1 vssd1 vccd1 vccd1 _11072_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput77 _12413_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[15] sky130_fd_sc_hd__buf_2
Xoutput88 _12671_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[25] sky130_fd_sc_hd__buf_2
XFILLER_103_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput99 _12150_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[6] sky130_fd_sc_hd__buf_2
XFILLER_163_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10023_ _10470_/S vssd1 vssd1 vccd1 vccd1 _10328_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14900_ _14897_/X _14899_/X _14916_/S vssd1 vssd1 vccd1 vccd1 _14900_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17027__A _17094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_1_clock clkbuf_1_0_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_103_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15880_ _09261_/A _15875_/X _15879_/X input52/X vssd1 vssd1 vccd1 vccd1 _15881_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input23_A io_dbus_rdata[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ _12870_/B _12807_/B _14869_/A vssd1 vssd1 vccd1 vccd1 _14832_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09471__C _09471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13077__A2 _13071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17550_ _19681_/Q vssd1 vssd1 vccd1 vccd1 _17551_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14762_ _12866_/A _11660_/A _09272_/C _14761_/Y _14812_/A vssd1 vssd1 vccd1 vccd1
+ _14763_/D sky130_fd_sc_hd__a311o_1
X_11974_ _11650_/X _14758_/B _11653_/X _11661_/X vssd1 vssd1 vccd1 vccd1 _11999_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA_clkbuf_leaf_57_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16501_ _16501_/A vssd1 vssd1 vccd1 vccd1 _19234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13713_ _13713_/A vssd1 vssd1 vccd1 vccd1 _18480_/D sky130_fd_sc_hd__clkbuf_1
X_17481_ _17176_/X _19647_/Q _17481_/S vssd1 vssd1 vccd1 vccd1 _17482_/A sky130_fd_sc_hd__mux2_1
X_10925_ _10920_/Y _10922_/Y _10719_/A _10924_/Y vssd1 vssd1 vccd1 vccd1 _10925_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14693_ _14693_/A vssd1 vssd1 vccd1 vccd1 _18798_/D sky130_fd_sc_hd__clkbuf_1
X_16432_ _16432_/A vssd1 vssd1 vccd1 vccd1 _19204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19220_ _20037_/CLK _19220_/D vssd1 vssd1 vccd1 vccd1 _19220_/Q sky130_fd_sc_hd__dfxtp_1
X_13644_ _18471_/Q _13643_/X _13670_/S vssd1 vssd1 vccd1 vccd1 _13645_/A sky130_fd_sc_hd__mux2_1
X_10856_ _10856_/A vssd1 vssd1 vccd1 vccd1 _10856_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15774__A1 _09261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19151_ _20003_/CLK _19151_/D vssd1 vssd1 vccd1 vccd1 _19151_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16363_/A vssd1 vssd1 vccd1 vccd1 _19179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13575_ _18462_/Q _13574_/X _13575_/S vssd1 vssd1 vccd1 vccd1 _13576_/A sky130_fd_sc_hd__mux2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10419__A _18853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ _10787_/A vssd1 vssd1 vccd1 vccd1 _10787_/X sky130_fd_sc_hd__buf_4
XFILLER_169_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18102_ _18101_/X _19902_/Q _18112_/S vssd1 vssd1 vccd1 vccd1 _18103_/A sky130_fd_sc_hd__mux2_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15314_ _15073_/X _15313_/X _15331_/S vssd1 vssd1 vccd1 vccd1 _15314_/X sky130_fd_sc_hd__mux2_1
X_19082_ _19864_/CLK _19082_/D vssd1 vssd1 vccd1 vccd1 _19082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12526_ _12521_/Y _12525_/Y _12814_/S vssd1 vssd1 vccd1 vccd1 _12526_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11260__A1 _11050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15526__A1 _18861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10694__S0 _10521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16294_ _16294_/A vssd1 vssd1 vccd1 vccd1 _19158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18033_ _18033_/A vssd1 vssd1 vccd1 vccd1 _19881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _15025_/X _15035_/X _15347_/S vssd1 vssd1 vccd1 vccd1 _15245_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12457_ _12514_/B vssd1 vssd1 vccd1 vccd1 _15385_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output91_A _12743_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11012__A1 _11291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__S0 _10319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _11960_/A _12823_/B vssd1 vssd1 vccd1 vccd1 _11408_/X sky130_fd_sc_hd__or2_1
X_15176_ _15176_/A vssd1 vssd1 vccd1 vccd1 _18838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12388_ _12334_/A _12334_/B _12364_/A _12387_/X vssd1 vssd1 vccd1 vccd1 _12389_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_125_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14127_ _14135_/D vssd1 vssd1 vccd1 vccd1 _14133_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11339_ _19194_/Q _19785_/Q _19947_/Q _19162_/Q _10618_/A _11021_/A vssd1 vssd1 vccd1
+ vccd1 _11340_/B sky130_fd_sc_hd__mux4_1
X_19984_ _20016_/CLK _19984_/D vssd1 vssd1 vccd1 vccd1 _19984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18935_ _18967_/CLK _18935_/D vssd1 vssd1 vccd1 vccd1 _18935_/Q sky130_fd_sc_hd__dfxtp_1
X_14058_ _18594_/Q _14053_/B _14057_/Y vssd1 vssd1 vccd1 vccd1 _18594_/D sky130_fd_sc_hd__o21a_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12512__A1 _11904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ _18795_/Q _11841_/A _11817_/X _12165_/A _13008_/X vssd1 vssd1 vccd1 vccd1
+ _13009_/X sky130_fd_sc_hd__a221o_1
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18866_ _18997_/CLK _18866_/D vssd1 vssd1 vccd1 vccd1 _18866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17817_ _19785_/Q _17001_/X _17821_/S vssd1 vssd1 vccd1 vccd1 _17818_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18797_ _19062_/CLK _18797_/D vssd1 vssd1 vccd1 vccd1 _18797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17748_ _17748_/A vssd1 vssd1 vccd1 vccd1 _19754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17679_ _17678_/X _19732_/Q _17682_/S vssd1 vssd1 vccd1 vccd1 _17680_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12809__A _14993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19418_ _20038_/CLK _19418_/D vssd1 vssd1 vccd1 vccd1 _19418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_194_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19656_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19349_ _20039_/CLK _19349_/D vssd1 vssd1 vccd1 vccd1 _19349_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10329__A _10329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17400__A _17411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10437__S0 _10328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13359__B _13359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_132_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18547_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09935_ _09929_/A _09934_/X _09690_/A vssd1 vssd1 vccd1 vccd1 _09935_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09866_ _09868_/A _09865_/X _09568_/X vssd1 vssd1 vccd1 vccd1 _09866_/X sky130_fd_sc_hd__o21a_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_147_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _18745_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_86_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _10382_/A vssd1 vssd1 vccd1 vccd1 _09798_/A sky130_fd_sc_hd__buf_2
XANTENNA__18377__S _18385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clock clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10710_/A vssd1 vssd1 vccd1 vccd1 _10710_/X sky130_fd_sc_hd__buf_2
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16953__A0 _16345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11690_/A vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10641_ _10690_/A _10637_/X _10640_/X vssd1 vssd1 vccd1 vccd1 _10641_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10239__A _18859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13360_ _13360_/A _18857_/Q vssd1 vssd1 vccd1 vccd1 _13360_/X sky130_fd_sc_hd__or2_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10572_ _10572_/A _10572_/B vssd1 vssd1 vccd1 vccd1 _10572_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12311_ _12188_/X _12306_/X _12307_/X _12310_/Y vssd1 vssd1 vccd1 vccd1 _12312_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13291_ _18474_/Q _11755_/X _12881_/X _18698_/Q _13290_/X vssd1 vssd1 vccd1 vccd1
+ _13291_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15030_ _14872_/X _14908_/X _15039_/S vssd1 vssd1 vccd1 vccd1 _15030_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10428__S0 _10152_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ _12242_/A _14868_/A vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__or2_1
XFILLER_123_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ _11997_/X _12171_/X _12172_/X vssd1 vssd1 vccd1 vccd1 _12173_/X sky130_fd_sc_hd__a21o_4
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09763__A _10438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ _11124_/A vssd1 vssd1 vccd1 vccd1 _11125_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15484__B _15487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16981_ _16981_/A vssd1 vssd1 vccd1 vccd1 _19447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18720_ _18744_/CLK _18720_/D vssd1 vssd1 vccd1 vccd1 _18720_/Q sky130_fd_sc_hd__dfxtp_1
X_15932_ _19003_/Q _15942_/A vssd1 vssd1 vccd1 vccd1 _15932_/X sky130_fd_sc_hd__and2_1
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11055_ _19135_/Q _19396_/Q _19295_/Q _19630_/Q _11367_/S _11320_/A vssd1 vssd1 vccd1
+ vccd1 _11056_/B sky130_fd_sc_hd__mux4_1
X_10006_ _19217_/Q _19808_/Q _19970_/Q _19185_/Q _10275_/A _09747_/A vssd1 vssd1 vccd1
+ vccd1 _10007_/B sky130_fd_sc_hd__mux4_1
XFILLER_37_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11517__B _12850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15863_ _15883_/A vssd1 vssd1 vccd1 vccd1 _15881_/A sky130_fd_sc_hd__clkbuf_1
X_18651_ _18653_/CLK _18651_/D vssd1 vssd1 vccd1 vccd1 _18651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18287__S _18291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17602_ _17154_/X _19704_/Q _17606_/S vssd1 vssd1 vccd1 vccd1 _17603_/A sky130_fd_sc_hd__mux2_1
X_14814_ _14814_/A _14814_/B _14814_/C _11980_/D vssd1 vssd1 vccd1 vccd1 _14815_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15794_ _15879_/A vssd1 vssd1 vccd1 vccd1 _15834_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18582_ _18745_/CLK _18582_/D vssd1 vssd1 vccd1 vccd1 _18582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14828__B _15004_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17533_ _17533_/A vssd1 vssd1 vccd1 vccd1 _19672_/D sky130_fd_sc_hd__clkbuf_1
X_14745_ _14745_/A _14745_/B vssd1 vssd1 vccd1 vccd1 _14800_/A sky130_fd_sc_hd__nor2_2
XFILLER_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11957_ _11949_/X _12432_/B _12432_/C vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__and3b_2
XANTENNA__11533__A _11533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17464_ _17151_/X _19639_/Q _17470_/S vssd1 vssd1 vccd1 vccd1 _17465_/A sky130_fd_sc_hd__mux2_1
X_10908_ _09830_/A _10907_/X _10947_/A vssd1 vssd1 vccd1 vccd1 _10908_/X sky130_fd_sc_hd__a21o_1
X_14676_ _14676_/A vssd1 vssd1 vccd1 vccd1 _18790_/D sky130_fd_sc_hd__clkbuf_1
X_11888_ _13081_/A vssd1 vssd1 vccd1 vccd1 _12889_/A sky130_fd_sc_hd__buf_2
X_19203_ _20020_/CLK _19203_/D vssd1 vssd1 vccd1 vccd1 _19203_/Q sky130_fd_sc_hd__dfxtp_1
X_16415_ _16472_/S vssd1 vssd1 vccd1 vccd1 _16424_/S sky130_fd_sc_hd__clkbuf_4
X_13627_ _19009_/Q _13627_/B vssd1 vssd1 vccd1 vccd1 _13627_/X sky130_fd_sc_hd__or2_1
X_10839_ _10832_/Y _10834_/Y _10836_/Y _10838_/Y _09551_/A vssd1 vssd1 vccd1 vccd1
+ _10839_/X sky130_fd_sc_hd__o221a_2
X_17395_ _17395_/A vssd1 vssd1 vccd1 vccd1 _19608_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16535__S _16541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14750__C_N _09471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16346_ _16345_/X _19174_/Q _16346_/S vssd1 vssd1 vccd1 vccd1 _16347_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09938__A _10277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11233__A1 _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19134_ _19757_/CLK _19134_/D vssd1 vssd1 vccd1 vccd1 _19134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13558_ _18460_/Q _13557_/X _13575_/S vssd1 vssd1 vccd1 vccd1 _13559_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10441__C1 _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19065_ _19978_/CLK _19065_/D vssd1 vssd1 vccd1 vccd1 _19065_/Q sky130_fd_sc_hd__dfxtp_1
X_12509_ _12347_/X _12507_/X _12508_/Y _12350_/X vssd1 vssd1 vccd1 vccd1 _12509_/X
+ sky130_fd_sc_hd__a31o_1
X_16277_ _16277_/A vssd1 vssd1 vccd1 vccd1 _19150_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13489_ _18821_/Q _12880_/X _11817_/X _18788_/Q vssd1 vssd1 vccd1 vccd1 _13489_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18016_ _19874_/Q _17081_/X _18020_/S vssd1 vssd1 vccd1 vccd1 _18017_/A sky130_fd_sc_hd__mux2_1
X_15228_ _15206_/X _15226_/X _15331_/S vssd1 vssd1 vccd1 vccd1 _15228_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15159_ _15384_/A vssd1 vssd1 vccd1 vccd1 _15159_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15394__B _15397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19967_ _19999_/CLK _19967_/D vssd1 vssd1 vccd1 vccd1 _19967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _20026_/CLK sky130_fd_sc_hd__clkbuf_16
X_09720_ _11348_/S vssd1 vssd1 vccd1 vccd1 _09721_/A sky130_fd_sc_hd__clkbuf_4
X_18918_ _18918_/CLK _18918_/D vssd1 vssd1 vccd1 vccd1 _18918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19898_ _19899_/CLK _19898_/D vssd1 vssd1 vccd1 vccd1 _19898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09651_ _10655_/S vssd1 vssd1 vccd1 vccd1 _09652_/A sky130_fd_sc_hd__buf_2
XFILLER_83_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18849_ _18851_/CLK _18849_/D vssd1 vssd1 vccd1 vccd1 _18849_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09582_ _10069_/A vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_79_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 _19942_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13213__A2 _12876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09848__A _09848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10432__C1 _09806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10493__S _10493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19949_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15910__A1 _11292_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17276__S _17276_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16180__S _16184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09583__A _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09918_ _19252_/Q _19747_/Q _09918_/S vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__mux2_1
XFILLER_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10522__A _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20038_ _20038_/CLK _20038_/D vssd1 vssd1 vccd1 vccd1 _20038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09849_ _09849_/A vssd1 vssd1 vccd1 vccd1 _09849_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10241__B _12858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _12866_/A _12866_/B _12860_/C vssd1 vssd1 vccd1 vccd1 _12861_/A sky130_fd_sc_hd__and3_2
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _13511_/B vssd1 vssd1 vccd1 vccd1 _12188_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12791_/A _12791_/B vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__and2_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13452__A2 _11755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _18744_/Q _14528_/B _14529_/Y vssd1 vssd1 vccd1 vccd1 _18744_/D sky130_fd_sc_hd__o21a_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _18748_/Q _11677_/B _11701_/A _18774_/Q vssd1 vssd1 vccd1 vccd1 _11743_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14461_ _14495_/A _14461_/B _14461_/C vssd1 vssd1 vccd1 vccd1 _18719_/D sky130_fd_sc_hd__nor3_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _14547_/A _14546_/A vssd1 vssd1 vccd1 vccd1 _13510_/B sky130_fd_sc_hd__or2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16200_ _13323_/X _19117_/Q _16206_/S vssd1 vssd1 vccd1 vccd1 _16201_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13412_ _13188_/A _18860_/Q _12957_/X vssd1 vssd1 vccd1 vccd1 _13412_/Y sky130_fd_sc_hd__a21oi_1
X_10624_ _10624_/A vssd1 vssd1 vccd1 vccd1 _10625_/A sky130_fd_sc_hd__buf_2
X_17180_ _17180_/A vssd1 vssd1 vccd1 vccd1 _17193_/S sky130_fd_sc_hd__buf_4
X_14392_ _14400_/D vssd1 vssd1 vccd1 vccd1 _14398_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16131_ _13354_/X _19087_/Q _16133_/S vssd1 vssd1 vccd1 vccd1 _16132_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11766__A2 _11764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13343_ _17065_/A vssd1 vssd1 vccd1 vccd1 _17707_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10555_ _10557_/A _10554_/X _10107_/A vssd1 vssd1 vccd1 vccd1 _10555_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16062_ _16062_/A vssd1 vssd1 vccd1 vccd1 _19058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13274_ _14078_/A _11683_/X _11733_/X _18633_/Q vssd1 vssd1 vccd1 vccd1 _13274_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15901__A1 _15900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10486_ _10480_/A _10485_/X _10382_/X vssd1 vssd1 vccd1 vccd1 _10486_/Y sky130_fd_sc_hd__o21ai_1
X_15013_ _14953_/X _14955_/X _15014_/S vssd1 vssd1 vccd1 vccd1 _15013_/X sky130_fd_sc_hd__mux2_1
X_12225_ _12234_/A _12277_/D vssd1 vssd1 vccd1 vccd1 _12226_/B sky130_fd_sc_hd__or2_1
XANTENNA__11074__S0 _11063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12912__A _18940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19821_ _19821_/CLK _19821_/D vssd1 vssd1 vccd1 vccd1 _19821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12156_ _15633_/B vssd1 vssd1 vccd1 vccd1 _12556_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_111_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11528__A _15980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ _11107_/A vssd1 vssd1 vccd1 vccd1 _11108_/A sky130_fd_sc_hd__buf_2
XANTENNA__12479__A0 _12470_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19752_ _20010_/CLK _19752_/D vssd1 vssd1 vccd1 vccd1 _19752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16964_ _16361_/X _19440_/Q _16964_/S vssd1 vssd1 vccd1 vccd1 _16965_/A sky130_fd_sc_hd__mux2_1
X_12087_ _12143_/A vssd1 vssd1 vccd1 vccd1 _15183_/A sky130_fd_sc_hd__buf_2
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18703_ _18819_/CLK _18703_/D vssd1 vssd1 vccd1 vccd1 _18703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11038_ _11032_/A _11037_/X _09774_/A vssd1 vssd1 vccd1 vccd1 _11038_/Y sky130_fd_sc_hd__o21ai_1
X_15915_ _15915_/A vssd1 vssd1 vccd1 vccd1 _18998_/D sky130_fd_sc_hd__clkbuf_1
X_19683_ _19683_/CLK _19683_/D vssd1 vssd1 vccd1 vccd1 _19683_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15417__A0 _18852_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16895_ _16364_/X _19409_/Q _16903_/S vssd1 vssd1 vccd1 vccd1 _16896_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11151__B1 _11095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18634_ _19683_/CLK _18634_/D vssd1 vssd1 vccd1 vccd1 _18634_/Q sky130_fd_sc_hd__dfxtp_1
X_15846_ _15846_/A vssd1 vssd1 vccd1 vccd1 _18976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11129__S1 _11050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18565_ _20005_/CLK _18565_/D vssd1 vssd1 vccd1 vccd1 _18565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15777_ _15777_/A _15783_/B vssd1 vssd1 vccd1 vccd1 _15777_/X sky130_fd_sc_hd__or2_1
X_12989_ _18618_/Q _11686_/A _13082_/A _14459_/B vssd1 vssd1 vccd1 vccd1 _12989_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17516_ _19664_/Q vssd1 vssd1 vccd1 vccd1 _17517_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__11454__A1 _11223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14728_ _14728_/A vssd1 vssd1 vccd1 vccd1 _18814_/D sky130_fd_sc_hd__clkbuf_1
X_18496_ _19731_/CLK _18496_/D vssd1 vssd1 vccd1 vccd1 _18496_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17447_ _17447_/A vssd1 vssd1 vccd1 vccd1 _19631_/D sky130_fd_sc_hd__clkbuf_1
X_14659_ _18786_/Q _13733_/X _14667_/S vssd1 vssd1 vccd1 vccd1 _14660_/B sky130_fd_sc_hd__mux2_1
XANTENNA__16265__S _16269_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14574__A _14577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17378_ _17424_/S vssd1 vssd1 vccd1 vccd1 _17387_/S sky130_fd_sc_hd__buf_2
XFILLER_146_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11757__A2 _11755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12806__B _12807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19117_ _19966_/CLK _19117_/D vssd1 vssd1 vccd1 vccd1 _19117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16329_ _17665_/A vssd1 vssd1 vccd1 vccd1 _16329_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048_ _19999_/CLK _19048_/D vssd1 vssd1 vccd1 vccd1 _19048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15609__S _15611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10193__A1 _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17824__S _17832_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__A _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09703_ _19386_/Q vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14749__A _14749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09634_ _09868_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09634_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17125__A _17662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13653__A _18884_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10040__S1 _10028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09565_ _09565_/A vssd1 vssd1 vccd1 vccd1 _09566_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09496_ _09496_/A _11941_/B vssd1 vssd1 vccd1 vccd1 _11912_/A sky130_fd_sc_hd__nor2_2
XFILLER_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09578__A _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14395__B1 _14366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17795__A _17795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18390__S _18396_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16903__S _16903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10340_ _10344_/A _10340_/B vssd1 vssd1 vccd1 vccd1 _10340_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15344__C1 _15275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10271_ _19215_/Q _19806_/Q _19968_/Q _19183_/Q _10059_/S _10261_/X vssd1 vssd1 vccd1
+ vccd1 _10271_/X sky130_fd_sc_hd__mux4_2
X_12010_ _12722_/B vssd1 vssd1 vccd1 vccd1 _12010_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10803__S0 _10787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10184__A1 _10182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13039__S _13350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11779__A_N _12060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13961_ _18561_/Q _13964_/C _11884_/X vssd1 vssd1 vccd1 vccd1 _13961_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14870__A1 _15449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13563__A _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ _18940_/Q vssd1 vssd1 vccd1 vccd1 _15735_/A sky130_fd_sc_hd__buf_4
XFILLER_74_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15700_ _15700_/A vssd1 vssd1 vccd1 vccd1 _18926_/D sky130_fd_sc_hd__clkbuf_1
X_16680_ _16680_/A vssd1 vssd1 vccd1 vccd1 _19314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09972__S1 _09612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ _12501_/A _13883_/X _12481_/X _12484_/Y _13890_/X vssd1 vssd1 vccd1 vccd1
+ _18535_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12843_ _12843_/A _12844_/B vssd1 vssd1 vccd1 vccd1 _12843_/Y sky130_fd_sc_hd__nor2_8
X_15631_ _18896_/Q _18928_/Q _15901_/S vssd1 vssd1 vccd1 vccd1 _15632_/A sky130_fd_sc_hd__mux2_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14622__A1 _11764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_opt_4_0_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18350_ _17735_/X _20008_/Q _18350_/S vssd1 vssd1 vccd1 vccd1 _18351_/A sky130_fd_sc_hd__mux2_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15562_ _15562_/A vssd1 vssd1 vccd1 vccd1 _18864_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _18786_/Q _12774_/B vssd1 vssd1 vccd1 vccd1 _12799_/B sky130_fd_sc_hd__and2_1
XFILLER_61_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17301_/A vssd1 vssd1 vccd1 vccd1 _19566_/D sky130_fd_sc_hd__clkbuf_1
X_14513_ _14513_/A vssd1 vssd1 vccd1 vccd1 _14518_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11531__S1 _09614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11725_ _13926_/A vssd1 vssd1 vccd1 vccd1 _14159_/A sky130_fd_sc_hd__buf_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18281_ _18337_/A vssd1 vssd1 vccd1 vccd1 _18350_/S sky130_fd_sc_hd__buf_6
XANTENNA__16085__S _16089_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15493_ _18858_/Q _15053_/X _15482_/Y _15492_/X vssd1 vssd1 vccd1 vccd1 _18858_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13502__S _13502_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17232_ _17128_/X _19536_/Q _17232_/S vssd1 vssd1 vccd1 vccd1 _17233_/A sky130_fd_sc_hd__mux2_1
X_14444_ _18709_/Q _18708_/Q _14440_/C _15807_/A vssd1 vssd1 vccd1 vccd1 _14445_/B
+ sky130_fd_sc_hd__a31o_1
X_11656_ _11667_/A _14761_/B _11975_/A vssd1 vssd1 vccd1 vccd1 _11656_/Y sky130_fd_sc_hd__nor3_1
XFILLER_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12626__B _12722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17163_ _17700_/A vssd1 vssd1 vccd1 vccd1 _17163_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17909__S _17915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ _19208_/Q _19799_/Q _19961_/Q _19176_/Q _10655_/S _09607_/A vssd1 vssd1 vccd1
+ vccd1 _10608_/B sky130_fd_sc_hd__mux4_1
X_14375_ _14378_/B _14381_/D _14374_/Y vssd1 vssd1 vccd1 vccd1 _18688_/D sky130_fd_sc_hd__o21a_1
XANTENNA__16813__S _16819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11587_ _11629_/A _11586_/C _11586_/A vssd1 vssd1 vccd1 vccd1 _11588_/B sky130_fd_sc_hd__a21oi_1
XFILLER_7_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16114_ _13219_/X _19079_/Q _16122_/S vssd1 vssd1 vccd1 vccd1 _16115_/A sky130_fd_sc_hd__mux2_1
X_13326_ _18886_/Q _18887_/Q _13326_/C vssd1 vssd1 vccd1 vccd1 _13357_/C sky130_fd_sc_hd__and3_1
X_17094_ _19484_/Q _17093_/X _17094_/S vssd1 vssd1 vccd1 vccd1 _17095_/A sky130_fd_sc_hd__mux2_1
X_10538_ _10539_/A _12849_/B vssd1 vssd1 vccd1 vccd1 _10540_/A sky130_fd_sc_hd__and2_1
XFILLER_156_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_180_clock_A _18998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16045_ _13385_/X _19051_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16046_/A sky130_fd_sc_hd__mux2_1
X_13257_ _13257_/A vssd1 vssd1 vccd1 vccd1 _13257_/Y sky130_fd_sc_hd__inv_2
X_10469_ _19371_/Q _19706_/Q _10469_/S vssd1 vssd1 vccd1 vccd1 _10469_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ _12208_/A vssd1 vssd1 vccd1 vccd1 _12322_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10175__A1 _09702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13188_ _13188_/A vssd1 vssd1 vccd1 vccd1 _13188_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10175__B2 _18860_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19804_ _19966_/CLK _19804_/D vssd1 vssd1 vccd1 vccd1 _19804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17644__S _17650_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12139_ _12139_/A _12139_/B vssd1 vssd1 vccd1 vccd1 _12140_/A sky130_fd_sc_hd__and2_1
XANTENNA__10162__A _10162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17996_ _19865_/Q _17052_/X _17998_/S vssd1 vssd1 vccd1 vccd1 _17997_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19735_ _19993_/CLK _19735_/D vssd1 vssd1 vccd1 vccd1 _19735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16947_ _16336_/X _19432_/Q _16953_/S vssd1 vssd1 vccd1 vccd1 _16948_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19666_ _20023_/CLK _19666_/D vssd1 vssd1 vccd1 vccd1 _19666_/Q sky130_fd_sc_hd__dfxtp_1
X_16878_ _16878_/A vssd1 vssd1 vccd1 vccd1 _19401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18617_ _18653_/CLK _18617_/D vssd1 vssd1 vccd1 vccd1 _18617_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11705__B _14227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15829_ _15829_/A vssd1 vssd1 vccd1 vccd1 _18971_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13416__A2 _11815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19597_ _19951_/CLK _19597_/D vssd1 vssd1 vccd1 vccd1 _19597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09350_ _09425_/B _09347_/X _09215_/X _09349_/Y vssd1 vssd1 vccd1 vccd1 _12061_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18548_ _18548_/CLK _18548_/D vssd1 vssd1 vccd1 vccd1 _18548_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11978__A2 _11971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09281_ _09274_/A _09272_/A _09279_/X _09280_/Y vssd1 vssd1 vccd1 vccd1 _09289_/B
+ sky130_fd_sc_hd__o211a_2
X_18479_ _18544_/CLK _18479_/D vssd1 vssd1 vccd1 vccd1 _18479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17315__A0 _17144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10089__S1 _10028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17819__S _17821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10337__A _10434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16723__S _16725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11286__S0 _11273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__B1 _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11060__C1 _11133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13648__A _13648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09845__B _12864_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13888__C1 _13946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13352__A1 _12967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12155__A2 _12150_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15863__A _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14301__B1 _14792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14852__A1 _09289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14479__A _14479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18043__A1 hold7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09617_ _19524_/Q vssd1 vssd1 vccd1 vccd1 _11068_/A sky130_fd_sc_hd__inv_2
XFILLER_83_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18385__S _18385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16694__A _16762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11418__A1 _11131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ _19526_/Q vssd1 vssd1 vccd1 vccd1 _09549_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09479_ _13307_/A vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__buf_2
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11510_ _11508_/Y _11510_/B vssd1 vssd1 vccd1 vccd1 _11510_/X sky130_fd_sc_hd__and2b_1
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12490_ _15397_/A _12490_/B vssd1 vssd1 vccd1 vccd1 _12493_/A sky130_fd_sc_hd__xor2_4
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11441_ _19352_/Q _19687_/Q _11441_/S vssd1 vssd1 vccd1 vccd1 _11441_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11277__S0 _11121_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14942__A _15094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12394__A2 _12390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14160_ _14427_/A vssd1 vssd1 vccd1 vccd1 _14160_/X sky130_fd_sc_hd__buf_2
XFILLER_164_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11372_ _19321_/Q _19592_/Q _19816_/Q _19560_/Q _10980_/A _10972_/A vssd1 vssd1 vccd1
+ vccd1 _11372_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09890__S0 _11553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ _13110_/A _13131_/C _12957_/A vssd1 vssd1 vccd1 vccd1 _13111_/X sky130_fd_sc_hd__o21a_1
XFILLER_166_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10323_ _10312_/A _10317_/X _10322_/X vssd1 vssd1 vccd1 vccd1 _10323_/Y sky130_fd_sc_hd__o21ai_1
X_14091_ _18606_/Q _14088_/B _14090_/Y vssd1 vssd1 vccd1 vccd1 _18606_/D sky130_fd_sc_hd__o21a_1
XANTENNA_input53_A io_ibus_inst[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13042_ _17656_/A vssd1 vssd1 vccd1 vccd1 _13042_/X sky130_fd_sc_hd__clkbuf_2
X_10254_ _10254_/A _19247_/Q vssd1 vssd1 vccd1 vccd1 _10254_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17464__S _17470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17850_ _19800_/Q _17049_/X _17854_/S vssd1 vssd1 vccd1 vccd1 _17851_/A sky130_fd_sc_hd__mux2_1
X_10185_ _10185_/A vssd1 vssd1 vccd1 vccd1 _10185_/X sky130_fd_sc_hd__buf_2
XFILLER_132_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16801_ _16801_/A vssd1 vssd1 vccd1 vccd1 _19367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17781_ _17781_/A vssd1 vssd1 vccd1 vccd1 _19769_/D sky130_fd_sc_hd__clkbuf_1
X_14993_ _14993_/A _14993_/B _14993_/C vssd1 vssd1 vccd1 vccd1 _15102_/A sky130_fd_sc_hd__or3_1
XFILLER_115_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19520_ _20007_/CLK _19520_/D vssd1 vssd1 vccd1 vccd1 _19520_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18034__A1 _14562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16732_ _19337_/Q _13813_/X _16736_/S vssd1 vssd1 vccd1 vccd1 _16733_/A sky130_fd_sc_hd__mux2_1
X_13944_ _13945_/B _13945_/C _18556_/Q vssd1 vssd1 vccd1 vccd1 _13946_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__16045__A0 _13385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_127_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19451_ _19877_/CLK _19451_/D vssd1 vssd1 vccd1 vccd1 _19451_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11525__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16663_ _16361_/X _19307_/Q _16663_/S vssd1 vssd1 vccd1 vccd1 _16664_/A sky130_fd_sc_hd__mux2_1
X_13875_ _12204_/A _12204_/B _13870_/X vssd1 vssd1 vccd1 vccd1 _18525_/D sky130_fd_sc_hd__a21o_1
XANTENNA__16808__S _16808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18402_ _18402_/A vssd1 vssd1 vccd1 vccd1 _20030_/D sky130_fd_sc_hd__clkbuf_1
X_15614_ _13688_/A _18920_/Q _15622_/S vssd1 vssd1 vccd1 vccd1 _15615_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12826_ _12827_/A _12826_/B vssd1 vssd1 vccd1 vccd1 _12826_/Y sky130_fd_sc_hd__nor2_8
X_19382_ _20007_/CLK _19382_/D vssd1 vssd1 vccd1 vccd1 _19382_/Q sky130_fd_sc_hd__dfxtp_1
X_16594_ _19276_/Q _13822_/X _16602_/S vssd1 vssd1 vccd1 vccd1 _16595_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18333_ _17710_/X _20000_/Q _18335_/S vssd1 vssd1 vccd1 vccd1 _18334_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13740__B _19024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _15151_/X _15047_/B _15544_/X _15413_/X vssd1 vssd1 vccd1 vccd1 _15545_/X
+ sky130_fd_sc_hd__a211o_1
X_12757_ _14993_/A _15520_/A _12736_/B vssd1 vssd1 vccd1 vccd1 _12758_/B sky130_fd_sc_hd__a21bo_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11708_ _12946_/A vssd1 vssd1 vccd1 vccd1 _13164_/B sky130_fd_sc_hd__buf_2
X_18264_ _18264_/A vssd1 vssd1 vccd1 vccd1 _19969_/D sky130_fd_sc_hd__clkbuf_1
X_15476_ _15544_/A _15476_/B _15476_/C vssd1 vssd1 vccd1 vccd1 _15476_/X sky130_fd_sc_hd__and3_1
X_12688_ _15972_/C _18923_/Q _12782_/S vssd1 vssd1 vccd1 vccd1 _12715_/A sky130_fd_sc_hd__mux2_8
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17215_ _17103_/X _19528_/Q _17221_/S vssd1 vssd1 vccd1 vccd1 _17216_/A sky130_fd_sc_hd__mux2_1
X_14427_ _14427_/A vssd1 vssd1 vccd1 vccd1 _14427_/X sky130_fd_sc_hd__clkbuf_2
X_11639_ _11639_/A _11639_/B vssd1 vssd1 vccd1 vccd1 _11639_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_156_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10157__A _10434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18195_ _18195_/A vssd1 vssd1 vccd1 vccd1 _19938_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16543__S _16545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17146_ _17146_/A vssd1 vssd1 vccd1 vccd1 _19504_/D sky130_fd_sc_hd__clkbuf_1
X_14358_ _18684_/Q _14356_/C _14357_/Y vssd1 vssd1 vccd1 vccd1 _18684_/D sky130_fd_sc_hd__o21a_1
XFILLER_143_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10396__A1 _09702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10396__B2 _18854_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13309_ _13306_/X _13326_/C _13308_/Y vssd1 vssd1 vccd1 vccd1 _13309_/X sky130_fd_sc_hd__a21o_1
X_17077_ _17077_/A vssd1 vssd1 vccd1 vccd1 _19478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14289_ _18662_/Q _14285_/B _14288_/Y vssd1 vssd1 vccd1 vccd1 _18662_/D sky130_fd_sc_hd__o21a_1
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16028_ _16028_/A vssd1 vssd1 vccd1 vccd1 _19043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14531__B1 _14507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09633__S0 _09598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17374__S _17376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17979_ _19857_/Q _17026_/X _17987_/S vssd1 vssd1 vccd1 vccd1 _17980_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13407__S _13464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19718_ _19846_/CLK _19718_/D vssd1 vssd1 vccd1 vccd1 _19718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19649_ _19942_/CLK _19649_/D vssd1 vssd1 vccd1 vccd1 _19649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09402_ _11703_/A _11671_/A _09402_/C _09402_/D vssd1 vssd1 vccd1 vccd1 _09410_/B
+ sky130_fd_sc_hd__nor4_1
XANTENNA__13931__A _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ _18936_/Q vssd1 vssd1 vccd1 vccd1 _17098_/B sky130_fd_sc_hd__buf_4
XFILLER_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09264_ _11961_/B _09264_/B _09264_/C _09316_/B vssd1 vssd1 vccd1 vccd1 _09265_/D
+ sky130_fd_sc_hd__or4_2
XANTENNA__11281__C1 _11133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16453__S _16457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09195_ _09274_/A vssd1 vssd1 vccd1 vccd1 _11950_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17839__A1 _17033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10234__S1 _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__09591__A _10724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11990_ _12044_/A _14898_/A vssd1 vssd1 vccd1 vccd1 _11993_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__14002__A _14010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10941_ _18842_/Q _09538_/A _09546_/A _10940_/X vssd1 vssd1 vccd1 vccd1 _12239_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16628__S _16630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18409__A _18409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13660_ _13660_/A vssd1 vssd1 vccd1 vccd1 _13660_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10872_ _19234_/Q _19729_/Q _10872_/S vssd1 vssd1 vccd1 vccd1 _10872_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12611_ _14749_/A _12657_/A _12682_/A _12610_/Y vssd1 vssd1 vccd1 vccd1 _12612_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_169_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13560__B _13560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13587_/X _13588_/X _13589_/Y _13590_/X _19004_/Q vssd1 vssd1 vccd1 vccd1
+ _13591_/X sky130_fd_sc_hd__a32o_4
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15330_ _15189_/X _15191_/X _15347_/S vssd1 vssd1 vccd1 vccd1 _15330_/X sky130_fd_sc_hd__mux2_1
X_12542_ _10444_/A _18917_/Q _12687_/A vssd1 vssd1 vccd1 vccd1 _14860_/A sky130_fd_sc_hd__mux2_2
XANTENNA__10170__S0 _10152_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17459__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15261_ _18842_/Q _09433_/X _15260_/X vssd1 vssd1 vccd1 vccd1 _18842_/D sky130_fd_sc_hd__o21a_1
XFILLER_61_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ _12501_/A _12501_/C vssd1 vssd1 vccd1 vccd1 _12478_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14672__A _14672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17000_ _17000_/A vssd1 vssd1 vccd1 vccd1 _19454_/D sky130_fd_sc_hd__clkbuf_1
X_14212_ _18643_/Q _18642_/Q _14212_/C vssd1 vssd1 vccd1 vccd1 _14215_/B sky130_fd_sc_hd__and3_1
XANTENNA__09766__A _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _19192_/Q _19783_/Q _19945_/Q _19160_/Q _11409_/S _11320_/A vssd1 vssd1 vccd1
+ vccd1 _11425_/B sky130_fd_sc_hd__mux4_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15192_ _15191_/X _14982_/X _15298_/S vssd1 vssd1 vccd1 vccd1 _15192_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15487__B _15487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10378__A1 _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09863__S0 _09598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__B1 _09843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14143_ _14143_/A _14143_/B _14143_/C vssd1 vssd1 vccd1 vccd1 _18620_/D sky130_fd_sc_hd__nor3_1
XANTENNA_clkbuf_leaf_53_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11355_ _11404_/A vssd1 vssd1 vccd1 vccd1 _11401_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10306_ _19935_/Q _19549_/Q _19999_/Q _19118_/Q _10354_/S _10182_/X vssd1 vssd1 vccd1
+ vccd1 _10307_/B sky130_fd_sc_hd__mux4_1
XFILLER_153_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14074_ _14090_/A _14078_/C vssd1 vssd1 vccd1 vccd1 _14074_/Y sky130_fd_sc_hd__nor2_1
X_18951_ _18956_/CLK _18951_/D vssd1 vssd1 vccd1 vccd1 _18951_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_106_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ _19195_/Q _19786_/Q _19948_/Q _19163_/Q _11273_/A _11073_/X vssd1 vssd1 vccd1
+ vccd1 _11287_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09615__S0 _09598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17902_ _19823_/Q _17020_/X _17904_/S vssd1 vssd1 vccd1 vccd1 _17903_/A sky130_fd_sc_hd__mux2_1
X_13025_ _13023_/X _18429_/Q _13116_/S vssd1 vssd1 vccd1 vccd1 _13026_/A sky130_fd_sc_hd__mux2_1
X_10237_ _10344_/A _10236_/X _09798_/A vssd1 vssd1 vccd1 vccd1 _10237_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11422__S0 _11212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18882_ _18918_/CLK _18882_/D vssd1 vssd1 vccd1 vccd1 _18882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17833_ _17833_/A vssd1 vssd1 vccd1 vccd1 _19792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10168_ _10210_/A _10167_/X _10001_/A vssd1 vssd1 vccd1 vccd1 _10168_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17922__S _17926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17764_ _17764_/A vssd1 vssd1 vccd1 vccd1 _19761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10099_ _19344_/Q _19615_/Q _19839_/Q _19583_/Q _10277_/S _10082_/A vssd1 vssd1 vccd1
+ vccd1 _10099_/X sky130_fd_sc_hd__mux4_1
X_14976_ _09347_/X _14803_/X _14972_/X _14975_/X vssd1 vssd1 vccd1 vccd1 _18833_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19503_ _19636_/CLK _19503_/D vssd1 vssd1 vccd1 vccd1 _19503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16715_ _16715_/A vssd1 vssd1 vccd1 vccd1 _19329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16569__A1 _13787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13927_ _14745_/A vssd1 vssd1 vccd1 vccd1 _14507_/A sky130_fd_sc_hd__clkbuf_1
X_17695_ _17694_/X _19737_/Q _17698_/S vssd1 vssd1 vccd1 vccd1 _17696_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15442__S _15480_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19434_ _19764_/CLK _19434_/D vssd1 vssd1 vccd1 vccd1 _19434_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17223__A _17280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16646_ _16336_/X _19299_/Q _16652_/S vssd1 vssd1 vccd1 vccd1 _16647_/A sky130_fd_sc_hd__mux2_1
X_13858_ _18517_/Q _13857_/X _13858_/S vssd1 vssd1 vccd1 vccd1 _13859_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15241__A1 _12221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19365_ _19764_/CLK _19365_/D vssd1 vssd1 vccd1 vccd1 _19365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12809_ _14993_/A vssd1 vssd1 vccd1 vccd1 _14990_/A sky130_fd_sc_hd__clkbuf_2
X_16577_ _16577_/A vssd1 vssd1 vccd1 vccd1 _19268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12367__A _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13789_ _13789_/A vssd1 vssd1 vccd1 vccd1 _18495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18316_ _17684_/X _19992_/Q _18324_/S vssd1 vssd1 vccd1 vccd1 _18317_/A sky130_fd_sc_hd__mux2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ _15553_/A _15531_/A vssd1 vssd1 vccd1 vccd1 _15528_/X sky130_fd_sc_hd__or2_1
Xclkbuf_2_3_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_19296_ _19985_/CLK _19296_/D vssd1 vssd1 vccd1 vccd1 _19296_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09379__C _11777_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18247_ _18247_/A vssd1 vssd1 vccd1 vccd1 _19961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14582__A _14595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15459_ _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15459_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09676__A _10073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18178_ _17694_/X _19931_/Q _18180_/S vssd1 vssd1 vccd1 vccd1 _18179_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17129_ _17128_/X _19499_/Q _17129_/S vssd1 vssd1 vccd1 vccd1 _17130_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09951_ _19380_/Q _19715_/Q _10094_/S vssd1 vssd1 vccd1 vccd1 _09951_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09882_ _09882_/A vssd1 vssd1 vccd1 vccd1 _09883_/A sky130_fd_sc_hd__clkbuf_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11413__S0 _11328_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12830__A _12831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09931__B1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17832__S _17832_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12818__B1 _18788_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15848__A1_N input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15480__A1 _15479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15232__A1 _15139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09316_ _09316_/A _09316_/B vssd1 vssd1 vccd1 vccd1 _09500_/B sky130_fd_sc_hd__or2_1
XFILLER_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16691__B _16691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09247_ _18973_/Q _09247_/B _09247_/C vssd1 vssd1 vccd1 vccd1 _09316_/B sky130_fd_sc_hd__or3_4
XFILLER_31_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09586__A _09586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13546__B2 _18999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ _18974_/Q vssd1 vssd1 vccd1 vccd1 _09283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15100__B _15100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11140_ _11140_/A _11140_/B vssd1 vssd1 vccd1 vccd1 _11140_/X sky130_fd_sc_hd__or2_1
Xclkbuf_4_5_0_clock clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_122_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18237__A1 _17675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput78 _12443_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[16] sky130_fd_sc_hd__buf_2
X_11071_ _18431_/Q _19460_/Q _19497_/Q _19071_/Q _11049_/S _10973_/A vssd1 vssd1 vccd1
+ vccd1 _11071_/X sky130_fd_sc_hd__mux4_1
Xoutput89 _12693_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[26] sky130_fd_sc_hd__buf_2
XFILLER_103_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10022_ _10529_/S vssd1 vssd1 vccd1 vccd1 _10470_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_76_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14830_ _15419_/A vssd1 vssd1 vccd1 vccd1 _14830_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10260__A _10260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09471__D _14750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input16_A io_dbus_rdata[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11973_ _12285_/A vssd1 vssd1 vccd1 vccd1 _12366_/B sky130_fd_sc_hd__clkbuf_2
X_14761_ _15738_/A _14761_/B _14761_/C vssd1 vssd1 vccd1 vccd1 _14761_/Y sky130_fd_sc_hd__nor3_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16500_ _19234_/Q _13790_/X _16508_/S vssd1 vssd1 vccd1 vccd1 _16501_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17043__A _17075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10924_ _10936_/A _10924_/B vssd1 vssd1 vccd1 vccd1 _10924_/Y sky130_fd_sc_hd__nor2_1
X_13712_ _18480_/Q _13711_/X _13752_/S vssd1 vssd1 vccd1 vccd1 _13713_/A sky130_fd_sc_hd__mux2_1
X_17480_ _17480_/A vssd1 vssd1 vccd1 vccd1 _19646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14692_ _18798_/Q _13572_/X _14694_/S vssd1 vssd1 vccd1 vccd1 _14693_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10391__S0 _10469_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ _19204_/Q _13797_/X _16435_/S vssd1 vssd1 vccd1 vccd1 _16432_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13290__B _13290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17978__A _18024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ _10893_/A vssd1 vssd1 vccd1 vccd1 _10856_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13643_ _11748_/X _13642_/Y _13689_/S vssd1 vssd1 vccd1 vccd1 _13643_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19150_ _19999_/CLK _19150_/D vssd1 vssd1 vccd1 vccd1 _19150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11245__C1 _09817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13785__A1 _13784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16362_ _16361_/X _19179_/Q _16362_/S vssd1 vssd1 vccd1 vccd1 _16363_/A sky130_fd_sc_hd__mux2_1
X_13574_ _13572_/X _13573_/Y _13583_/S vssd1 vssd1 vccd1 vccd1 _13574_/X sky130_fd_sc_hd__mux2_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _10954_/S vssd1 vssd1 vccd1 vccd1 _10787_/A sky130_fd_sc_hd__buf_2
XFILLER_9_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10143__S0 _10141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18101_ _18854_/Q _13677_/X _18101_/S vssd1 vssd1 vccd1 vccd1 _18101_/X sky130_fd_sc_hd__mux2_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15313_ _15166_/X _15168_/X _15347_/S vssd1 vssd1 vccd1 vccd1 _15313_/X sky130_fd_sc_hd__mux2_1
X_12525_ _12525_/A _12576_/C vssd1 vssd1 vccd1 vccd1 _12525_/Y sky130_fd_sc_hd__nor2_1
X_19081_ _19864_/CLK _19081_/D vssd1 vssd1 vccd1 vccd1 _19081_/Q sky130_fd_sc_hd__dfxtp_1
X_16293_ _13481_/X _19158_/Q _16295_/S vssd1 vssd1 vccd1 vccd1 _16294_/A sky130_fd_sc_hd__mux2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12915__A _15735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18032_ _18027_/X _19881_/Q _18044_/S vssd1 vssd1 vccd1 vccd1 _18033_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12456_ _11904_/X _12848_/B _12455_/Y vssd1 vssd1 vccd1 vccd1 _12514_/B sky130_fd_sc_hd__a21oi_1
X_15244_ _15244_/A vssd1 vssd1 vccd1 vccd1 _15244_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09836__S0 _09733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12634__B _12856_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ _09701_/A _11397_/X _11406_/X _09841_/A _18834_/Q vssd1 vssd1 vccd1 vccd1
+ _12823_/B sky130_fd_sc_hd__a32o_2
X_15175_ _18838_/Q _15173_/X _15480_/S vssd1 vssd1 vccd1 vccd1 _15176_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10446__S1 _10320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12387_ _12329_/A _12361_/A _12361_/B vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__o21ba_1
XFILLER_153_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output84_A _12574_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ _18615_/Q _18614_/Q _18745_/Q _14126_/D vssd1 vssd1 vccd1 vccd1 _14135_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_4_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ _09847_/A _11327_/X _11337_/X _09536_/A _18835_/Q vssd1 vssd1 vccd1 vccd1
+ _11452_/A sky130_fd_sc_hd__a32o_2
XFILLER_154_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19983_ _20015_/CLK _19983_/D vssd1 vssd1 vccd1 vccd1 _19983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18228__A1 _17662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14057_ _14090_/A _14062_/C vssd1 vssd1 vccd1 vccd1 _14057_/Y sky130_fd_sc_hd__nor2_1
X_18934_ _18967_/CLK _18934_/D vssd1 vssd1 vccd1 vccd1 _18934_/Q sky130_fd_sc_hd__dfxtp_1
X_11269_ _12827_/B _11223_/X _12828_/B _12118_/A vssd1 vssd1 vccd1 vccd1 _11269_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13008_ _18459_/Q _11740_/X _12944_/A _18683_/Q _13007_/X vssd1 vssd1 vccd1 vccd1
+ _13008_/X sky130_fd_sc_hd__a221o_1
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12512__A2 _12850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18865_ _18997_/CLK _18865_/D vssd1 vssd1 vccd1 vccd1 _18865_/Q sky130_fd_sc_hd__dfxtp_1
X_17816_ _17816_/A vssd1 vssd1 vccd1 vccd1 _19784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18796_ _19887_/CLK _18796_/D vssd1 vssd1 vccd1 vccd1 _18796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12276__A1 _12234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17747_ _17646_/X _19754_/Q _17749_/S vssd1 vssd1 vccd1 vccd1 _17748_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14959_ _15103_/B vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14577__A _14577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11484__C1 _09874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17678_ _17678_/A vssd1 vssd1 vccd1 vccd1 _17678_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19417_ _19747_/CLK _19417_/D vssd1 vssd1 vccd1 vccd1 _19417_/Q sky130_fd_sc_hd__dfxtp_1
X_16629_ _16629_/A vssd1 vssd1 vccd1 vccd1 _19291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13776__A1 _13774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19348_ _20037_/CLK _19348_/D vssd1 vssd1 vccd1 vccd1 _19348_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10134__S0 _09653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11787__B1 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19279_ _19936_/CLK _19279_/D vssd1 vssd1 vccd1 vccd1 _19279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16714__A1 _13787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10685__S1 _10010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12544__B _14860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13656__A _13656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09934_ _20037_/Q _19875_/Q _19284_/Q _19054_/Q _09668_/S _09614_/A vssd1 vssd1 vccd1
+ vccd1 _09934_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09865_ _18453_/Q _19482_/Q _19519_/Q _19093_/Q _09635_/X _09851_/A vssd1 vssd1 vccd1
+ vccd1 _09865_/X sky130_fd_sc_hd__mux4_1
XANTENNA_input8_A io_dbus_rdata[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11711__B1 _14555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _09796_/A vssd1 vssd1 vccd1 vccd1 _10382_/A sky130_fd_sc_hd__buf_2
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16178__S _16184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14487__A _14495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16906__S _16914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10640_ _10638_/X _10639_/X _10630_/A vssd1 vssd1 vccd1 vccd1 _10640_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ _19672_/Q _19438_/Q _18503_/Q _19768_/Q _10521_/X _10522_/X vssd1 vssd1 vccd1
+ vccd1 _10572_/B sky130_fd_sc_hd__mux4_1
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12310_ _12344_/A _12308_/Y _12374_/C _12366_/B vssd1 vssd1 vccd1 vccd1 _12310_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_10_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13290_ _19901_/Q _13290_/B vssd1 vssd1 vccd1 vccd1 _13290_/X sky130_fd_sc_hd__and2_1
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12241_ _12242_/A _14868_/A vssd1 vssd1 vccd1 vccd1 _12241_/X sky130_fd_sc_hd__and2_1
XANTENNA__10428__S1 _10153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10202__B1 _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ _12191_/A _12234_/B vssd1 vssd1 vccd1 vccd1 _12172_/X sky130_fd_sc_hd__and2_1
XFILLER_162_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11123_ _11328_/A vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16980_ _16384_/X _19447_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16981_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11054_ _11410_/S vssd1 vssd1 vccd1 vccd1 _11367_/S sky130_fd_sc_hd__buf_4
X_15931_ _19002_/Q _15927_/X _15928_/X _15930_/Y vssd1 vssd1 vccd1 vccd1 _19002_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10005_ _10005_/A vssd1 vssd1 vccd1 vccd1 _10275_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11086__A _11086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18650_ _18653_/CLK _18650_/D vssd1 vssd1 vccd1 vccd1 _18650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15862_ _15862_/A vssd1 vssd1 vccd1 vccd1 _18981_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17601_ _17601_/A vssd1 vssd1 vccd1 vccd1 _19703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14813_ _14813_/A _14813_/B _14813_/C vssd1 vssd1 vccd1 vccd1 _14814_/C sky130_fd_sc_hd__or3_1
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18581_ _18744_/CLK _18581_/D vssd1 vssd1 vccd1 vccd1 _18581_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output122_A _12853_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15793_ input45/X vssd1 vssd1 vccd1 vccd1 _15793_/Y sky130_fd_sc_hd__inv_6
XANTENNA__13455__B1 _11687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17532_ _19672_/Q vssd1 vssd1 vccd1 vccd1 _17533_/A sky130_fd_sc_hd__clkbuf_1
X_14744_ _15856_/A _14744_/B vssd1 vssd1 vccd1 vccd1 _14745_/B sky130_fd_sc_hd__nor2_2
XFILLER_18_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11956_ _11956_/A _11956_/B _11956_/C vssd1 vssd1 vccd1 vccd1 _12432_/C sky130_fd_sc_hd__and3_1
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10364__S0 _10356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17463_ _17463_/A vssd1 vssd1 vccd1 vccd1 _19638_/D sky130_fd_sc_hd__clkbuf_1
X_10907_ _19234_/Q _19729_/Q _10907_/S vssd1 vssd1 vccd1 vccd1 _10907_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11887_ _09411_/Y _16836_/A _11773_/A vssd1 vssd1 vccd1 vccd1 _11887_/Y sky130_fd_sc_hd__a21oi_1
X_14675_ _18790_/Q _14554_/X _14683_/S vssd1 vssd1 vccd1 vccd1 _14676_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19202_ _19957_/CLK _19202_/D vssd1 vssd1 vccd1 vccd1 _19202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16414_ _16414_/A vssd1 vssd1 vccd1 vccd1 _19196_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14955__A0 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10838_ _10723_/A _10837_/X _10719_/X vssd1 vssd1 vccd1 vccd1 _10838_/Y sky130_fd_sc_hd__o21ai_1
X_13626_ _13626_/A vssd1 vssd1 vccd1 vccd1 _18468_/D sky130_fd_sc_hd__clkbuf_1
X_17394_ _19608_/Q _17049_/X _17398_/S vssd1 vssd1 vccd1 vccd1 _17395_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10116__S0 _09595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19133_ _19758_/CLK _19133_/D vssd1 vssd1 vccd1 vccd1 _19133_/Q sky130_fd_sc_hd__dfxtp_1
X_16345_ _17681_/A vssd1 vssd1 vccd1 vccd1 _16345_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12430__A1 _15847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769_ _19140_/Q _19401_/Q _19300_/Q _19635_/Q _10921_/S _10663_/A vssd1 vssd1 vccd1
+ vccd1 _10770_/B sky130_fd_sc_hd__mux4_1
X_13557_ _13553_/X _13556_/Y _13583_/S vssd1 vssd1 vccd1 vccd1 _13557_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19064_ _20010_/CLK _19064_/D vssd1 vssd1 vccd1 vccd1 _19064_/Q sky130_fd_sc_hd__dfxtp_1
X_12508_ _12508_/A _12532_/C vssd1 vssd1 vccd1 vccd1 _12508_/Y sky130_fd_sc_hd__nand2_1
X_16276_ _13344_/X _19150_/Q _16280_/S vssd1 vssd1 vccd1 vccd1 _16277_/A sky130_fd_sc_hd__mux2_1
X_13488_ _18709_/Q _12881_/X _13487_/X vssd1 vssd1 vccd1 vccd1 _13488_/X sky130_fd_sc_hd__a21o_1
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18015_ _18015_/A vssd1 vssd1 vccd1 vccd1 _19873_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15956__A _15964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17647__S _17650_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15227_ _15348_/S vssd1 vssd1 vccd1 vccd1 _15331_/S sky130_fd_sc_hd__clkbuf_2
X_12439_ _12411_/A _14877_/A _12386_/A vssd1 vssd1 vccd1 vccd1 _12439_/X sky130_fd_sc_hd__a21bo_1
XFILLER_126_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14860__A _14860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12194__B1 _12186_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15158_ _15099_/X _15154_/Y _15157_/X _15105_/X vssd1 vssd1 vccd1 vccd1 _15162_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14109_ _18612_/Q _14107_/B _14108_/Y vssd1 vssd1 vccd1 vccd1 _18612_/D sky130_fd_sc_hd__o21a_1
X_19966_ _19966_/CLK _19966_/D vssd1 vssd1 vccd1 vccd1 _19966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15089_ _15428_/A vssd1 vssd1 vccd1 vccd1 _15089_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18917_ _18918_/CLK _18917_/D vssd1 vssd1 vccd1 vccd1 _18917_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09392__C _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19897_ _19899_/CLK _19897_/D vssd1 vssd1 vccd1 vccd1 _19897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09650_ _09650_/A vssd1 vssd1 vccd1 vccd1 _10655_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18848_ _19792_/CLK _18848_/D vssd1 vssd1 vccd1 vccd1 _18848_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_clock clock vssd1 vssd1 vccd1 vccd1 clkbuf_0_clock/X sky130_fd_sc_hd__clkbuf_16
XFILLER_27_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09581_ _10266_/A vssd1 vssd1 vccd1 vccd1 _10069_/A sky130_fd_sc_hd__clkbuf_4
X_18779_ _18819_/CLK _18779_/D vssd1 vssd1 vccd1 vccd1 _18779_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13446__B1 _13368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_175_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17411__A _17411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_164_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09864__A _11538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13386__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09917_ _19683_/Q _19449_/Q _18514_/Q _19779_/Q _09920_/S _09647_/A vssd1 vssd1 vccd1
+ vccd1 _09917_/X sky130_fd_sc_hd__mux4_1
XANTENNA__18388__S _18396_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20037_ _20037_/CLK _20037_/D vssd1 vssd1 vccd1 vccd1 _20037_/Q sky130_fd_sc_hd__dfxtp_1
X_09848_ _09848_/A vssd1 vssd1 vccd1 vccd1 _09849_/A sky130_fd_sc_hd__buf_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09779_/A vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15977__A2 _14803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _12918_/B vssd1 vssd1 vccd1 vccd1 _13511_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12790_ _12790_/A vssd1 vssd1 vccd1 vccd1 _12790_/X sky130_fd_sc_hd__buf_2
XFILLER_73_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14010__A _14010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _18471_/Q _11740_/X _14672_/A _18807_/Q vssd1 vssd1 vccd1 vccd1 _11743_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12660__A1 _09261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11772_/A _11772_/B vssd1 vssd1 vccd1 vccd1 _14546_/A sky130_fd_sc_hd__or2b_1
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14460_ _14459_/B _14459_/C _18719_/Q vssd1 vssd1 vccd1 vccd1 _14461_/C sky130_fd_sc_hd__a21oi_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10623_ _10750_/S vssd1 vssd1 vccd1 vccd1 _10691_/S sky130_fd_sc_hd__clkbuf_4
X_13411_ _13714_/B _13427_/C vssd1 vssd1 vccd1 vccd1 _13411_/Y sky130_fd_sc_hd__xnor2_1
X_14391_ _18693_/Q _18692_/Q _18691_/Q _14391_/D vssd1 vssd1 vccd1 vccd1 _14400_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_128_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16130_ _16130_/A vssd1 vssd1 vccd1 vccd1 _19086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13342_ _13005_/X _13328_/X _13339_/X _13341_/X vssd1 vssd1 vccd1 vccd1 _17065_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_154_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10554_ _18441_/Q _19470_/Q _19507_/Q _19081_/Q _10125_/S _10497_/X vssd1 vssd1 vccd1
+ vccd1 _10554_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13273_ _18601_/Q vssd1 vssd1 vccd1 vccd1 _14078_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16061_ _19058_/Q _12161_/B _16073_/S vssd1 vssd1 vccd1 vccd1 _16062_/A sky130_fd_sc_hd__mux2_1
X_10485_ _20028_/Q _19866_/Q _19275_/Q _19045_/Q _09729_/A _10473_/X vssd1 vssd1 vccd1
+ vccd1 _10485_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09774__A _09774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15012_ _15009_/X _15011_/X _15113_/S vssd1 vssd1 vccd1 vccd1 _15012_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12224_ _12234_/A _12277_/D vssd1 vssd1 vccd1 vccd1 _12249_/B sky130_fd_sc_hd__nand2_1
XFILLER_170_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19820_ _19950_/CLK _19820_/D vssd1 vssd1 vccd1 vccd1 _19820_/Q sky130_fd_sc_hd__dfxtp_1
X_12155_ _12791_/A _12150_/Y _12153_/X _12154_/X vssd1 vssd1 vccd1 vccd1 _12155_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09493__B _15899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_64_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_193_clock clkbuf_opt_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19816_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11106_ _19385_/Q vssd1 vssd1 vccd1 vccd1 _11107_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19751_ _20010_/CLK _19751_/D vssd1 vssd1 vccd1 vccd1 _19751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16963_ _16963_/A vssd1 vssd1 vccd1 vccd1 _19439_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11528__B _12864_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12086_ _12537_/A _09495_/A _12084_/X _12085_/Y vssd1 vssd1 vccd1 vccd1 _12143_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_150_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18298__S _18302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18702_ _19912_/CLK _18702_/D vssd1 vssd1 vccd1 vccd1 _18702_/Q sky130_fd_sc_hd__dfxtp_1
X_11037_ _18432_/Q _19461_/Q _19498_/Q _19072_/Q _10892_/A _11022_/X vssd1 vssd1 vccd1
+ vccd1 _11037_/X sky130_fd_sc_hd__mux4_1
X_15914_ hold6/A _15913_/X _15914_/S vssd1 vssd1 vccd1 vccd1 _15915_/A sky130_fd_sc_hd__mux2_1
X_19682_ _20036_/CLK _19682_/D vssd1 vssd1 vccd1 vccd1 _19682_/Q sky130_fd_sc_hd__dfxtp_1
X_16894_ _16905_/A vssd1 vssd1 vccd1 vccd1 _16903_/S sky130_fd_sc_hd__buf_6
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15417__A1 _15416_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18633_ _19683_/CLK _18633_/D vssd1 vssd1 vccd1 vccd1 _18633_/Q sky130_fd_sc_hd__dfxtp_1
X_15845_ _15861_/A _17201_/B vssd1 vssd1 vccd1 vccd1 _15846_/A sky130_fd_sc_hd__and2_1
XANTENNA__10859__S _10859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15016__A _15016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18564_ _20005_/CLK _18564_/D vssd1 vssd1 vccd1 vccd1 _18564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15776_ _09263_/A _15765_/X _15775_/X _15769_/X vssd1 vssd1 vccd1 vccd1 _18956_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _18718_/Q vssd1 vssd1 vccd1 vccd1 _14459_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17515_ _17515_/A vssd1 vssd1 vccd1 vccd1 _19663_/D sky130_fd_sc_hd__clkbuf_1
X_14727_ _18814_/Q _11898_/X _14727_/S vssd1 vssd1 vccd1 vccd1 _14728_/A sky130_fd_sc_hd__mux2_1
X_18495_ _20018_/CLK _18495_/D vssd1 vssd1 vccd1 vccd1 _18495_/Q sky130_fd_sc_hd__dfxtp_1
X_11939_ _11939_/A _12290_/B _11939_/C vssd1 vssd1 vccd1 vccd1 _11940_/D sky130_fd_sc_hd__and3_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_131_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18544_/CLK sky130_fd_sc_hd__clkbuf_16
X_17446_ _17125_/X _19631_/Q _17448_/S vssd1 vssd1 vccd1 vccd1 _17447_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14658_ _14658_/A vssd1 vssd1 vccd1 vccd1 _18785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13600__A0 _11833_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ _19007_/Q _13609_/B vssd1 vssd1 vccd1 vccd1 _13609_/X sky130_fd_sc_hd__or2_1
X_17377_ _17377_/A vssd1 vssd1 vccd1 vccd1 _19600_/D sky130_fd_sc_hd__clkbuf_1
X_14589_ _14595_/A _14589_/B vssd1 vssd1 vccd1 vccd1 _14590_/A sky130_fd_sc_hd__and2_1
X_19116_ _19581_/CLK _19116_/D vssd1 vssd1 vccd1 vccd1 _19116_/Q sky130_fd_sc_hd__dfxtp_1
X_16328_ _16328_/A vssd1 vssd1 vccd1 vccd1 _19168_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_146_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _18693_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19047_ _19966_/CLK _19047_/D vssd1 vssd1 vccd1 vccd1 _19047_/Q sky130_fd_sc_hd__dfxtp_1
X_16259_ _16259_/A vssd1 vssd1 vccd1 vccd1 _19142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09684__A _10719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10623__A _10750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19949_ _19949_/CLK _19949_/D vssd1 vssd1 vccd1 vccd1 _19949_/Q sky130_fd_sc_hd__dfxtp_1
X_09702_ _09702_/A vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__buf_4
XANTENNA__15625__S _15901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18001__S _18009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11142__A1 _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09633_ _19222_/Q _19813_/Q _19975_/Q _19190_/Q _09598_/X _09614_/X vssd1 vssd1 vccd1
+ vccd1 _09634_/B sky130_fd_sc_hd__mux4_1
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11693__A2 _13081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15959__A2 _15951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09564_ _10107_/A vssd1 vssd1 vccd1 vccd1 _09565_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12269__B _12298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10102__C1 _09807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ _09495_/A vssd1 vssd1 vccd1 vccd1 _12536_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13198__A2 _13619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10956__A1 _10856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17287__S _17293_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10270_ _10270_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10270_/X sky130_fd_sc_hd__or2_1
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10803__S1 _10788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13960_ _18560_/Q _13957_/C _13959_/Y vssd1 vssd1 vccd1 vccd1 _18560_/D sky130_fd_sc_hd__o21a_1
XFILLER_101_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09533__S _15127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ _14225_/D vssd1 vssd1 vccd1 vccd1 _18352_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13891_ _12446_/A _13883_/X _12450_/Y _12453_/X _13890_/X vssd1 vssd1 vccd1 vccd1
+ _18534_/D sky130_fd_sc_hd__o221a_1
XFILLER_74_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15630_ _15630_/A vssd1 vssd1 vccd1 vccd1 _18895_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _12842_/A _12844_/B vssd1 vssd1 vccd1 vccd1 _12842_/Y sky130_fd_sc_hd__nor2_2
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _18864_/Q _15560_/X _15567_/S vssd1 vssd1 vccd1 vccd1 _15562_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16366__S _16378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _18786_/Q _12774_/B vssd1 vssd1 vccd1 vccd1 _12773_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17300_ _17122_/X _19566_/Q _17304_/S vssd1 vssd1 vccd1 vccd1 _17301_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14528_/A _14512_/B _14512_/C vssd1 vssd1 vccd1 vccd1 _18737_/D sky130_fd_sc_hd__nor3_1
X_18280_ _18280_/A _18280_/B vssd1 vssd1 vccd1 vccd1 _18337_/A sky130_fd_sc_hd__or2_4
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11715_/X _11717_/X _11721_/Y _11723_/X _19010_/Q vssd1 vssd1 vccd1 vccd1
+ _11724_/X sky130_fd_sc_hd__a32o_4
XFILLER_42_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _15089_/X _15490_/X _15491_/Y _15954_/A vssd1 vssd1 vccd1 vccd1 _15492_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_opt_8_0_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17231_/A vssd1 vssd1 vccd1 vccd1 _19535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14443_ _18708_/Q _14440_/C _18709_/Q vssd1 vssd1 vccd1 vccd1 _14445_/A sky130_fd_sc_hd__a21oi_1
X_11655_ _11655_/A _11657_/B vssd1 vssd1 vccd1 vccd1 _11667_/C sky130_fd_sc_hd__nor2_4
Xclkbuf_leaf_63_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19864_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10708__A _10919_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12397__B1 _13648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17162_ _17162_/A vssd1 vssd1 vccd1 vccd1 _19509_/D sky130_fd_sc_hd__clkbuf_1
X_10606_ _10832_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _10606_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11586_ _11586_/A _11629_/A _11586_/C vssd1 vssd1 vccd1 vccd1 _11588_/A sky130_fd_sc_hd__and3_1
X_14374_ _14378_/B _14381_/D _14366_/X vssd1 vssd1 vccd1 vccd1 _14374_/Y sky130_fd_sc_hd__a21oi_1
X_16113_ _16135_/A vssd1 vssd1 vccd1 vccd1 _16122_/S sky130_fd_sc_hd__buf_2
XFILLER_171_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13325_ _13325_/A vssd1 vssd1 vccd1 vccd1 _18445_/D sky130_fd_sc_hd__clkbuf_1
X_10537_ _09883_/A _10525_/X _10536_/X _09913_/A _10512_/Y vssd1 vssd1 vccd1 vccd1
+ _12849_/B sky130_fd_sc_hd__o32a_4
XANTENNA_clkbuf_leaf_123_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17093_ _17093_/A vssd1 vssd1 vccd1 vccd1 _17093_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12923__A _13502_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16044_ _16044_/A vssd1 vssd1 vccd1 vccd1 _16053_/S sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_78_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _20006_/CLK sky130_fd_sc_hd__clkbuf_16
X_10468_ _10480_/A _10468_/B vssd1 vssd1 vccd1 vccd1 _10468_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13256_ _13642_/A _13256_/B _13256_/C vssd1 vssd1 vccd1 vccd1 _13256_/X sky130_fd_sc_hd__and3_1
XFILLER_124_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _12263_/A vssd1 vssd1 vccd1 vccd1 _15234_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13361__A2 _11896_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13187_ _13245_/A vssd1 vssd1 vccd1 vccd1 _13188_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10399_ _19372_/Q _19707_/Q _10447_/S vssd1 vssd1 vccd1 vccd1 _10400_/B sky130_fd_sc_hd__mux2_1
XFILLER_151_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19803_ _19997_/CLK _19803_/D vssd1 vssd1 vccd1 vccd1 _19803_/Q sky130_fd_sc_hd__dfxtp_1
X_12138_ _13508_/A _12131_/X _12132_/X _12137_/Y _12402_/B vssd1 vssd1 vccd1 vccd1
+ _12139_/B sky130_fd_sc_hd__a311o_1
X_17995_ _17995_/A vssd1 vssd1 vccd1 vccd1 _19864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13754__A _16992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19734_ _19993_/CLK _19734_/D vssd1 vssd1 vccd1 vccd1 _19734_/Q sky130_fd_sc_hd__dfxtp_1
X_16946_ _16946_/A vssd1 vssd1 vccd1 vccd1 _19431_/D sky130_fd_sc_hd__clkbuf_1
X_12069_ _18760_/Q _12069_/B vssd1 vssd1 vccd1 vccd1 _12071_/C sky130_fd_sc_hd__xor2_1
XFILLER_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10558__S0 _10125_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19665_ _19731_/CLK _19665_/D vssd1 vssd1 vccd1 vccd1 _19665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13473__B _18863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16877_ _16339_/X _19401_/Q _16881_/S vssd1 vssd1 vccd1 vccd1 _16878_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16063__A1 _12188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18616_ _18653_/CLK _18616_/D vssd1 vssd1 vccd1 vccd1 _18616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17660__S _17666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15828_ _15831_/A _15828_/B vssd1 vssd1 vccd1 vccd1 _15829_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_16_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19950_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19596_ _19821_/CLK _19596_/D vssd1 vssd1 vccd1 vccd1 _19596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_48_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18547_ _18547_/CLK _18547_/D vssd1 vssd1 vccd1 vccd1 _18547_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__16276__S _16280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15759_ _09467_/X _15752_/X _15758_/Y _15756_/X vssd1 vssd1 vccd1 vccd1 _18949_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10635__B1 _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__A _10069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09280_ _09521_/A vssd1 vssd1 vccd1 vccd1 _09280_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_61_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18478_ _19900_/CLK _18478_/D vssd1 vssd1 vccd1 vccd1 _18478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10730__S0 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17429_ _17097_/X _19623_/Q _17437_/S vssd1 vssd1 vccd1 vccd1 _17430_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11721__B _19010_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10618__A _10618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12833__A _12833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17835__S _17843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11363__B2 _12956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12979__S _13003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14852__A2 _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09616_ _11538_/A _09616_/B vssd1 vssd1 vccd1 vccd1 _09616_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09547_ _09547_/A vssd1 vssd1 vccd1 vccd1 _09547_/X sky130_fd_sc_hd__buf_2
XANTENNA__14495__A _14495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09589__A _10921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09478_ _19486_/Q vssd1 vssd1 vccd1 vccd1 _13307_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_169_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15103__B _15103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16914__S _16914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _11440_/A _11440_/B vssd1 vssd1 vccd1 vccd1 _11440_/X sky130_fd_sc_hd__or2_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11277__S1 _11077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13040__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13040__B2 _12874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11371_ _19129_/Q _19390_/Q _19289_/Q _19624_/Q _11328_/X _11322_/X vssd1 vssd1 vccd1
+ vccd1 _11371_/X sky130_fd_sc_hd__mux4_2
XFILLER_125_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10322_ _10462_/A _10321_/X _10192_/A vssd1 vssd1 vccd1 vccd1 _10322_/X sky130_fd_sc_hd__o21a_1
X_13110_ _13110_/A _13131_/C vssd1 vssd1 vccd1 vccd1 _13110_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14090_ _14090_/A _14095_/C vssd1 vssd1 vccd1 vccd1 _14090_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17745__S _17749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13041_ _17014_/A vssd1 vssd1 vccd1 vccd1 _17656_/A sky130_fd_sc_hd__clkbuf_2
X_10253_ _19742_/Q vssd1 vssd1 vccd1 vccd1 _10253_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16817__A0 _16374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10184_ _10182_/X _10183_/X _10112_/A vssd1 vssd1 vccd1 vccd1 _10184_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input46_A io_ibus_inst[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16800_ _16348_/X _19367_/Q _16808_/S vssd1 vssd1 vccd1 vccd1 _16801_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17490__A0 _17189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17046__A _17046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17780_ _17694_/X _19769_/Q _17782_/S vssd1 vssd1 vccd1 vccd1 _17781_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14992_ _15055_/S _14996_/B vssd1 vssd1 vccd1 vccd1 _15002_/B sky130_fd_sc_hd__nand2_1
XFILLER_120_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16731_ _16731_/A vssd1 vssd1 vccd1 vccd1 _19336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13943_ _13945_/B _13945_/C _13942_/Y vssd1 vssd1 vccd1 vccd1 _18555_/D sky130_fd_sc_hd__o21a_1
XFILLER_101_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19450_ _20006_/CLK _19450_/D vssd1 vssd1 vccd1 vccd1 _19450_/Q sky130_fd_sc_hd__dfxtp_1
X_16662_ _16662_/A vssd1 vssd1 vccd1 vccd1 _19306_/D sky130_fd_sc_hd__clkbuf_1
X_13874_ _12790_/X _12171_/X _12172_/X _17203_/A vssd1 vssd1 vccd1 vccd1 _18524_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18401_ _17704_/X _20030_/Q _18407_/S vssd1 vssd1 vccd1 vccd1 _18402_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15613_ _15624_/A vssd1 vssd1 vccd1 vccd1 _15622_/S sky130_fd_sc_hd__clkbuf_2
X_19381_ _20006_/CLK _19381_/D vssd1 vssd1 vccd1 vccd1 _19381_/Q sky130_fd_sc_hd__dfxtp_1
X_12825_ _12827_/A _12825_/B vssd1 vssd1 vccd1 vccd1 _12825_/Y sky130_fd_sc_hd__nor2_8
X_16593_ _16604_/A vssd1 vssd1 vccd1 vccd1 _16602_/S sky130_fd_sc_hd__buf_4
XFILLER_62_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16096__S _16100_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12918__A _18827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18332_ _18332_/A vssd1 vssd1 vccd1 vccd1 _19999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ _15544_/A _15544_/B _15544_/C vssd1 vssd1 vccd1 vccd1 _15544_/X sky130_fd_sc_hd__and3_1
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12756_/A vssd1 vssd1 vccd1 vccd1 _14993_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _19969_/Q _17713_/A _18263_/S vssd1 vssd1 vccd1 vccd1 _18264_/A sky130_fd_sc_hd__mux2_1
X_11707_ _11707_/A vssd1 vssd1 vccd1 vccd1 _12946_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ _15305_/A _15470_/Y _15474_/Y vssd1 vssd1 vccd1 vccd1 _15476_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__10438__A _10438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16824__S _16830_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12687_ _12687_/A vssd1 vssd1 vccd1 vccd1 _12782_/S sky130_fd_sc_hd__clkbuf_4
X_17214_ _17214_/A vssd1 vssd1 vccd1 vccd1 _19527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14426_ _18703_/Q vssd1 vssd1 vccd1 vccd1 _14433_/C sky130_fd_sc_hd__clkbuf_1
X_18194_ _17716_/X _19938_/Q _18202_/S vssd1 vssd1 vccd1 vccd1 _18195_/A sky130_fd_sc_hd__mux2_1
X_11638_ _10242_/X _11647_/B _10246_/B vssd1 vssd1 vccd1 vccd1 _11639_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13031__B2 _18763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17145_ _17144_/X _19504_/Q _17145_/S vssd1 vssd1 vccd1 vccd1 _17146_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10872__S _10872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14357_ _18684_/Q _14356_/C _14332_/X vssd1 vssd1 vccd1 vccd1 _14357_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _11565_/X _11567_/X _11568_/X _11572_/A _09837_/X vssd1 vssd1 vccd1 vccd1
+ _11574_/B sky130_fd_sc_hd__o221a_1
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10396__A2 _10384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13308_ _13306_/X _13326_/C _13307_/X vssd1 vssd1 vccd1 vccd1 _13308_/Y sky130_fd_sc_hd__o21ai_1
X_17076_ _19478_/Q _17074_/X _17088_/S vssd1 vssd1 vccd1 vccd1 _17077_/A sky130_fd_sc_hd__mux2_1
X_14288_ _14288_/A _14297_/D vssd1 vssd1 vccd1 vccd1 _14288_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16027_ _13250_/X _19043_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15964__A _15964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ _13238_/X _18440_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _13240_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10779__S0 _10704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__S1 _09614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15175__S _15480_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17978_ _18024_/S vssd1 vssd1 vccd1 vccd1 _17987_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_111_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19717_ _20007_/CLK _19717_/D vssd1 vssd1 vccd1 vccd1 _19717_/Q sky130_fd_sc_hd__dfxtp_1
X_16929_ _16310_/X _19424_/Q _16931_/S vssd1 vssd1 vccd1 vccd1 _16930_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17390__S _17398_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19648_ _19971_/CLK _19648_/D vssd1 vssd1 vccd1 vccd1 _19648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10951__S0 _10907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09401_ _09401_/A _09408_/B vssd1 vssd1 vccd1 vccd1 _09402_/D sky130_fd_sc_hd__nor2_4
XFILLER_111_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14598__A1 _11833_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19579_ _19965_/CLK _19579_/D vssd1 vssd1 vccd1 vccd1 _19579_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15795__B1 _15789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12828__A _15899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09332_ _18983_/Q _18938_/Q vssd1 vssd1 vccd1 vccd1 _09697_/C sky130_fd_sc_hd__xnor2_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09263_ _09263_/A _09273_/A _18991_/Q vssd1 vssd1 vccd1 vccd1 _09264_/C sky130_fd_sc_hd__or3b_1
XANTENNA__16734__S _16736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09194_ _18974_/Q vssd1 vssd1 vccd1 vccd1 _09274_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17565__S _17573_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11336__A1 _11131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11887__A2 _16836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18396__S _18396_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17224__A0 _17115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ _10925_/X _10930_/X _10939_/X _09550_/A vssd1 vssd1 vccd1 vccd1 _10940_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10942__S0 _10907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ _10936_/A _10871_/B vssd1 vssd1 vccd1 vccd1 _10871_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12738__A _12738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_clock clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_71_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _12634_/A _12855_/B vssd1 vssd1 vccd1 vccd1 _12610_/Y sky130_fd_sc_hd__nor2_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13660_/A vssd1 vssd1 vccd1 vccd1 _13590_/X sky130_fd_sc_hd__clkbuf_2
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12541_ _12541_/A _15424_/A vssd1 vssd1 vccd1 vccd1 _12544_/A sky130_fd_sc_hd__xor2_1
XANTENNA__16644__S _16652_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10170__S1 _10153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15260_ _12246_/X _15146_/X _15259_/X _15951_/A vssd1 vssd1 vccd1 vccd1 _15260_/X
+ sky130_fd_sc_hd__a211o_1
X_12472_ _12472_/A vssd1 vssd1 vccd1 vccd1 _12522_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__14672__B _14672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14211_ _18642_/Q _14212_/C _14210_/Y vssd1 vssd1 vccd1 vccd1 _18642_/D sky130_fd_sc_hd__o21a_1
XANTENNA__11024__B1 _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11423_ _11332_/A _11422_/X _11003_/A vssd1 vssd1 vccd1 vccd1 _11423_/Y sky130_fd_sc_hd__o21ai_1
X_15191_ _15065_/X _15063_/X _15198_/S vssd1 vssd1 vccd1 vccd1 _15191_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12473__A _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11575__B2 _18864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__S1 _09851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11354_ _19130_/Q _19391_/Q _19290_/Q _19625_/Q _11155_/A _11172_/A vssd1 vssd1 vccd1
+ vccd1 _11354_/X sky130_fd_sc_hd__mux4_1
X_14142_ _18620_/Q _14142_/B _14142_/C vssd1 vssd1 vccd1 vccd1 _14143_/C sky130_fd_sc_hd__and3_1
XFILLER_4_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10783__C1 _09550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17475__S _17481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ _10305_/A _10305_/B vssd1 vssd1 vccd1 vccd1 _10305_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14073_ _14073_/A vssd1 vssd1 vccd1 vccd1 _14078_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18950_ _18958_/CLK _18950_/D vssd1 vssd1 vccd1 vccd1 _18950_/Q sky130_fd_sc_hd__dfxtp_2
X_11285_ _11070_/X _11284_/X _11003_/A vssd1 vssd1 vccd1 vccd1 _11285_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18160__A _18206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11327__A1 _09559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__S1 _09614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10236_ _20035_/Q _19873_/Q _19282_/Q _19052_/Q _10330_/S _10013_/A vssd1 vssd1 vccd1
+ vccd1 _10236_/X sky130_fd_sc_hd__mux4_1
X_13024_ _13502_/S vssd1 vssd1 vccd1 vccd1 _13116_/S sky130_fd_sc_hd__clkbuf_4
X_17901_ _17901_/A vssd1 vssd1 vccd1 vccd1 _19822_/D sky130_fd_sc_hd__clkbuf_1
X_18881_ _18918_/CLK _18881_/D vssd1 vssd1 vccd1 vccd1 _18881_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output152_A _12534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11422__S1 _11077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17832_ _19792_/Q _17023_/X _17832_/S vssd1 vssd1 vccd1 vccd1 _17833_/A sky130_fd_sc_hd__mux2_1
X_10167_ _19251_/Q _19746_/Q _10279_/A vssd1 vssd1 vccd1 vccd1 _10167_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17763_ _17668_/X _19761_/Q _17771_/S vssd1 vssd1 vccd1 vccd1 _17764_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10098_ _19152_/Q _19413_/Q _19312_/Q _19647_/Q _10094_/S _10278_/A vssd1 vssd1 vccd1
+ vccd1 _10098_/X sky130_fd_sc_hd__mux4_1
X_14975_ _12871_/Y _15482_/B _15940_/A vssd1 vssd1 vccd1 vccd1 _14975_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16819__S _16819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17215__A0 _17103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19502_ _19633_/CLK _19502_/D vssd1 vssd1 vccd1 vccd1 _19502_/Q sky130_fd_sc_hd__dfxtp_1
X_16714_ _19329_/Q _13787_/X _16714_/S vssd1 vssd1 vccd1 vccd1 _16715_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13926_ _13926_/A vssd1 vssd1 vccd1 vccd1 _14745_/A sky130_fd_sc_hd__buf_4
X_17694_ _17694_/A vssd1 vssd1 vccd1 vccd1 _17694_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19433_ _19796_/CLK _19433_/D vssd1 vssd1 vccd1 vccd1 _19433_/Q sky130_fd_sc_hd__dfxtp_1
X_16645_ _16645_/A vssd1 vssd1 vccd1 vccd1 _19298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13857_ _17093_/A vssd1 vssd1 vccd1 vccd1 _13857_/X sky130_fd_sc_hd__buf_2
XFILLER_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19364_ _19796_/CLK _19364_/D vssd1 vssd1 vccd1 vccd1 _19364_/Q sky130_fd_sc_hd__dfxtp_1
X_12808_ _15552_/A _14970_/B vssd1 vssd1 vccd1 vccd1 _12811_/A sky130_fd_sc_hd__nor2_2
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16576_ _19268_/Q _13797_/X _16580_/S vssd1 vssd1 vccd1 vccd1 _16577_/A sky130_fd_sc_hd__mux2_1
X_13788_ _18495_/Q _13787_/X _13788_/S vssd1 vssd1 vccd1 vccd1 _13789_/A sky130_fd_sc_hd__mux2_1
X_18315_ _18337_/A vssd1 vssd1 vccd1 vccd1 _18324_/S sky130_fd_sc_hd__buf_2
XFILLER_43_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ _15531_/A _15531_/B vssd1 vssd1 vccd1 vccd1 _15527_/Y sky130_fd_sc_hd__nand2_1
X_12739_ _12740_/A _15520_/B vssd1 vssd1 vccd1 vccd1 _12741_/A sky130_fd_sc_hd__and2_1
X_19295_ _19758_/CLK _19295_/D vssd1 vssd1 vccd1 vccd1 _19295_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16554__S _16558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18246_ _19961_/Q _17688_/A _18252_/S vssd1 vssd1 vccd1 vccd1 _18247_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09957__A _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15458_ _15458_/A vssd1 vssd1 vccd1 vccd1 _15458_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14409_ _18698_/Q _14411_/C _14409_/C vssd1 vssd1 vccd1 vccd1 _14410_/C sky130_fd_sc_hd__and3_1
X_18177_ _18177_/A vssd1 vssd1 vccd1 vccd1 _19930_/D sky130_fd_sc_hd__clkbuf_1
X_15389_ _15329_/X _15332_/X _15388_/X _15342_/X vssd1 vssd1 vccd1 vccd1 _15389_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17128_ _17665_/A vssd1 vssd1 vccd1 vccd1 _17128_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17385__S _17387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17059_ _17075_/A vssd1 vssd1 vccd1 vccd1 _17072_/S sky130_fd_sc_hd__clkbuf_8
X_09950_ _19252_/Q _19747_/Q _09950_/S vssd1 vssd1 vccd1 vccd1 _09950_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18070__A _18104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09692__A _09862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _09881_/A vssd1 vssd1 vccd1 vccd1 _09882_/A sky130_fd_sc_hd__buf_4
XFILLER_140_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11413__S1 _11073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12830__B _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09931__A1 _09933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10350__B _12854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09315_ _14822_/B _09315_/B vssd1 vssd1 vccd1 vccd1 _14782_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11254__B1 _09559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16464__S _16468_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ _09309_/A _09514_/A _09276_/C vssd1 vssd1 vccd1 vccd1 _09246_/X sky130_fd_sc_hd__or3_1
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09177_ _18975_/Q vssd1 vssd1 vccd1 vccd1 _09230_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14712__S _14716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11070_ _11332_/A vssd1 vssd1 vccd1 vccd1 _11070_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput79 _12470_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[17] sky130_fd_sc_hd__buf_2
XFILLER_163_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10021_ _10521_/A vssd1 vssd1 vccd1 vccd1 _10529_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_131_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09922__A1 _10069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14760_ _15539_/A vssd1 vssd1 vccd1 vccd1 _15553_/A sky130_fd_sc_hd__buf_2
X_11972_ input66/X _15633_/A vssd1 vssd1 vccd1 vccd1 _12285_/A sky130_fd_sc_hd__and2_2
XFILLER_72_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13711_ _13707_/Y _13710_/X _16066_/S vssd1 vssd1 vccd1 vccd1 _13711_/X sky130_fd_sc_hd__mux2_1
X_10923_ _19664_/Q _19430_/Q _18495_/Q _19760_/Q _10703_/A _10663_/A vssd1 vssd1 vccd1
+ vccd1 _10924_/B sky130_fd_sc_hd__mux4_1
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13571__B _19002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14691_ _14691_/A vssd1 vssd1 vccd1 vccd1 _18797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16420__A1 _13781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16430_ _16430_/A vssd1 vssd1 vccd1 vccd1 _19203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ _13642_/A _13646_/C vssd1 vssd1 vccd1 vccd1 _13642_/Y sky130_fd_sc_hd__xnor2_2
X_10854_ _10854_/A vssd1 vssd1 vccd1 vccd1 _10893_/A sky130_fd_sc_hd__buf_2
XFILLER_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _17697_/A vssd1 vssd1 vccd1 vccd1 _16361_/X sky130_fd_sc_hd__clkbuf_2
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _13580_/A _13580_/C vssd1 vssd1 vccd1 vccd1 _13573_/Y sky130_fd_sc_hd__xnor2_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _09848_/A _10772_/X _10784_/Y _09538_/A _18845_/Q vssd1 vssd1 vccd1 vccd1
+ _15938_/C sky130_fd_sc_hd__a32o_4
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10143__S1 _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18100_ _18100_/A vssd1 vssd1 vccd1 vccd1 _19901_/D sky130_fd_sc_hd__clkbuf_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _18845_/Q _15278_/X _15311_/X vssd1 vssd1 vccd1 vccd1 _18845_/D sky130_fd_sc_hd__o21a_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09777__A _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19080_ _20026_/CLK _19080_/D vssd1 vssd1 vccd1 vccd1 _19080_/Q sky130_fd_sc_hd__dfxtp_1
X_12524_ _18536_/Q _18537_/Q _12524_/C vssd1 vssd1 vccd1 vccd1 _12576_/C sky130_fd_sc_hd__and3_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _16292_/A vssd1 vssd1 vccd1 vccd1 _19157_/D sky130_fd_sc_hd__clkbuf_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12915__B _16691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18031_ _18134_/S vssd1 vssd1 vccd1 vccd1 _18044_/S sky130_fd_sc_hd__clkbuf_4
X_15243_ _15243_/A vssd1 vssd1 vccd1 vccd1 _15243_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12455_ _11982_/X _14763_/C _12318_/Y vssd1 vssd1 vccd1 vccd1 _12455_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__09836__S1 _09768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11406_ _09772_/A _11399_/X _11401_/X _11405_/X _09802_/A vssd1 vssd1 vccd1 vccd1
+ _11406_/X sky130_fd_sc_hd__a311o_2
X_15174_ _15945_/A vssd1 vssd1 vccd1 vccd1 _15480_/S sky130_fd_sc_hd__clkbuf_4
X_12386_ _12386_/A _12386_/B vssd1 vssd1 vccd1 vccd1 _12389_/A sky130_fd_sc_hd__and2_2
XFILLER_126_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14125_ _14143_/A _14125_/B _14125_/C vssd1 vssd1 vccd1 vccd1 _18614_/D sky130_fd_sc_hd__nor3_1
X_11337_ _09559_/A _11330_/X _11332_/X _11336_/X _09872_/A vssd1 vssd1 vccd1 vccd1
+ _11337_/X sky130_fd_sc_hd__a311o_1
XFILLER_114_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19982_ _19982_/CLK _19982_/D vssd1 vssd1 vccd1 vccd1 _19982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14056_ _14056_/A vssd1 vssd1 vccd1 vccd1 _14062_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18933_ _18974_/CLK _18933_/D vssd1 vssd1 vccd1 vccd1 _18933_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output77_A _12413_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11268_ _18838_/Q _09537_/A _09546_/A _11267_/X vssd1 vssd1 vccd1 vccd1 _12118_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__17933__S _17937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ _19886_/Q _13209_/B vssd1 vssd1 vccd1 vccd1 _13007_/X sky130_fd_sc_hd__and2_1
X_10219_ _19681_/Q _19447_/Q _18512_/Q _19777_/Q _10388_/S _10223_/A vssd1 vssd1 vccd1
+ vccd1 _10220_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11199_ _11199_/A _11199_/B vssd1 vssd1 vccd1 vccd1 _11199_/X sky130_fd_sc_hd__and2_1
X_18864_ _18911_/CLK _18864_/D vssd1 vssd1 vccd1 vccd1 _18864_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17987__A1 _17039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17815_ _19784_/Q _16998_/X _17821_/S vssd1 vssd1 vccd1 vccd1 _17816_/A sky130_fd_sc_hd__mux2_1
X_18795_ _19887_/CLK _18795_/D vssd1 vssd1 vccd1 vccd1 _18795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13762__A _16998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17234__A _17280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17746_ _17746_/A vssd1 vssd1 vccd1 vccd1 _19753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14958_ _14954_/X _14957_/X _15121_/S vssd1 vssd1 vccd1 vccd1 _14958_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14670__A0 _11801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _18548_/Q _12820_/A _12796_/X _12800_/X _13904_/X vssd1 vssd1 vccd1 vccd1
+ _18548_/D sky130_fd_sc_hd__o221a_1
XFILLER_63_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17677_ _17677_/A vssd1 vssd1 vccd1 vccd1 _19731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14889_ _14931_/A vssd1 vssd1 vccd1 vccd1 _15020_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12378__A _12378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19416_ _19972_/CLK _19416_/D vssd1 vssd1 vccd1 vccd1 _19416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16628_ _16310_/X _19291_/Q _16630_/S vssd1 vssd1 vccd1 vccd1 _16629_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19347_ _19972_/CLK _19347_/D vssd1 vssd1 vccd1 vccd1 _19347_/Q sky130_fd_sc_hd__dfxtp_1
X_16559_ _16559_/A vssd1 vssd1 vccd1 vccd1 _19260_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10134__S1 _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11331__S0 _11328_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19278_ _20031_/CLK _19278_/D vssd1 vssd1 vccd1 vccd1 _19278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17911__A1 _17033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18229_ _18229_/A vssd1 vssd1 vccd1 vccd1 _19953_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14725__A1 _11879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10626__A _10626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_171_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13937__A _13946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12841__A _12841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09933_/X sky130_fd_sc_hd__or2_1
XANTENNA__15150__A1 _18837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11398__S0 _11356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17843__S _17843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11457__A _15923_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09864_ _11538_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09864_/X sky130_fd_sc_hd__or2_1
XFILLER_112_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11711__B2 _12452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10070__S0 _09597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09380__A2 _14227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _10579_/A vssd1 vssd1 vccd1 vccd1 _09796_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17144__A _17681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11570__S0 _11553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_96_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13216__B2 _13350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10570_ _10563_/Y _10565_/Y _10567_/Y _10569_/Y _09821_/A vssd1 vssd1 vccd1 vccd1
+ _10570_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09597__A _09597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09229_ _09481_/A _09481_/B _09481_/C _09481_/D vssd1 vssd1 vccd1 vccd1 _11951_/A
+ sky130_fd_sc_hd__nand4b_4
XANTENNA__15913__A0 _12082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14716__A1 _13661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14008__A _14044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12727__B1 _12234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ _12239_/Y _18906_/Q _12358_/S vssd1 vssd1 vccd1 vccd1 _14868_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10202__A1 _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12171_ _12155_/X _12159_/X _12168_/X _12170_/X vssd1 vssd1 vccd1 vccd1 _12171_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11122_ _11122_/A _11122_/B vssd1 vssd1 vccd1 vccd1 _11122_/X sky130_fd_sc_hd__and2_1
XFILLER_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11053_ _19522_/Q vssd1 vssd1 vccd1 vccd1 _11410_/S sky130_fd_sc_hd__clkbuf_2
X_15930_ _15936_/A _15930_/B vssd1 vssd1 vccd1 vccd1 _15930_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10004_ _10279_/A vssd1 vssd1 vccd1 vccd1 _10005_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18091__A0 _18851_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ _15861_/A _16837_/B vssd1 vssd1 vccd1 vccd1 _15862_/A sky130_fd_sc_hd__and2_1
XANTENNA__16369__S _16378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17600_ _17151_/X _19703_/Q _17606_/S vssd1 vssd1 vccd1 vccd1 _17601_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14812_ _14812_/A _14812_/B _14812_/C _11937_/B vssd1 vssd1 vccd1 vccd1 _14813_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18580_ _18744_/CLK _18580_/D vssd1 vssd1 vccd1 vccd1 _18580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15792_ _15792_/A vssd1 vssd1 vccd1 vccd1 _18961_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13455__A1 _14336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17531_ _17531_/A vssd1 vssd1 vccd1 vccd1 _19671_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17989__A _18011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14743_ _14743_/A vssd1 vssd1 vccd1 vccd1 _18821_/D sky130_fd_sc_hd__clkbuf_1
X_11955_ _09310_/C _09276_/X _11912_/A _14818_/A _09492_/A vssd1 vssd1 vccd1 vccd1
+ _11956_/C sky130_fd_sc_hd__o2111a_1
XANTENNA_output115_A _12844_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17462_ _17147_/X _19638_/Q _17470_/S vssd1 vssd1 vccd1 vccd1 _17463_/A sky130_fd_sc_hd__mux2_1
X_10906_ _19362_/Q _19697_/Q _10906_/S vssd1 vssd1 vccd1 vccd1 _10906_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14674_ _14742_/S vssd1 vssd1 vccd1 vccd1 _14683_/S sky130_fd_sc_hd__clkbuf_2
X_11886_ _14665_/A vssd1 vssd1 vccd1 vccd1 _16836_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19201_ _19824_/CLK _19201_/D vssd1 vssd1 vccd1 vccd1 _19201_/Q sky130_fd_sc_hd__dfxtp_1
X_16413_ _19196_/Q _13771_/X _16413_/S vssd1 vssd1 vccd1 vccd1 _16414_/A sky130_fd_sc_hd__mux2_1
X_13625_ _18468_/Q _13623_/X _13670_/S vssd1 vssd1 vccd1 vccd1 _13626_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14955__A1 _15078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10837_ _20020_/Q _19858_/Q _19267_/Q _19037_/Q _09650_/A _10049_/A vssd1 vssd1 vccd1
+ vccd1 _10837_/X sky130_fd_sc_hd__mux4_1
X_17393_ _17393_/A vssd1 vssd1 vccd1 vccd1 _19607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10116__S1 _10260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19132_ _19981_/CLK _19132_/D vssd1 vssd1 vccd1 vccd1 _19132_/Q sky130_fd_sc_hd__dfxtp_1
X_16344_ _16344_/A vssd1 vssd1 vccd1 vccd1 _19173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13556_ _13565_/B _13556_/B vssd1 vssd1 vccd1 vccd1 _13556_/Y sky130_fd_sc_hd__nand2_1
X_10768_ _19332_/Q _19603_/Q _19827_/Q _19571_/Q _11468_/S _10597_/A vssd1 vssd1 vccd1
+ vccd1 _10768_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19063_ _19063_/CLK _19063_/D vssd1 vssd1 vccd1 vccd1 _19063_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15904__A0 _15847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ _12508_/A _12532_/C vssd1 vssd1 vccd1 vccd1 _12507_/X sky130_fd_sc_hd__or2_1
X_16275_ _16275_/A vssd1 vssd1 vccd1 vccd1 _19149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16832__S _16834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ _19912_/Q _13290_/B _12982_/A _18485_/Q vssd1 vssd1 vccd1 vccd1 _13487_/X
+ sky130_fd_sc_hd__a22o_1
X_10699_ _18848_/Q vssd1 vssd1 vccd1 vccd1 _10699_/Y sky130_fd_sc_hd__inv_2
X_18014_ _19873_/Q _17078_/X _18020_/S vssd1 vssd1 vccd1 vccd1 _18015_/A sky130_fd_sc_hd__mux2_1
X_15226_ _14941_/A _14894_/X _15280_/S vssd1 vssd1 vccd1 vccd1 _15226_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12438_ _12438_/A vssd1 vssd1 vccd1 vccd1 _12438_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15956__B _15956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15157_ _15155_/X _15160_/B _15102_/X _15156_/X vssd1 vssd1 vccd1 vccd1 _15157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12369_ _12369_/A _12392_/B vssd1 vssd1 vccd1 vccd1 _12369_/X sky130_fd_sc_hd__and2_1
XFILLER_141_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14108_ _14146_/A _14108_/B vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__nor2_1
X_19965_ _19965_/CLK _19965_/D vssd1 vssd1 vccd1 vccd1 _19965_/Q sky130_fd_sc_hd__dfxtp_1
X_15088_ _15071_/X _15075_/X _15086_/X _15491_/A vssd1 vssd1 vccd1 vccd1 _15088_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_141_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17663__S _17666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15972__A _15978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18916_ _19350_/CLK _18916_/D vssd1 vssd1 vccd1 vccd1 _18916_/Q sky130_fd_sc_hd__dfxtp_1
X_14039_ _18588_/Q _14036_/B _14038_/Y vssd1 vssd1 vccd1 vccd1 _18588_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10181__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19896_ _19896_/CLK _19896_/D vssd1 vssd1 vccd1 vccd1 _19896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09993__S0 _09967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18847_ _19792_/CLK _18847_/D vssd1 vssd1 vccd1 vccd1 _18847_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09580_ _10200_/A vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13446__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18778_ _19900_/CLK _18778_/D vssd1 vssd1 vccd1 vccd1 _18778_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_118_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17729_ _17729_/A vssd1 vssd1 vccd1 vccd1 _17729_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13749__A2 _19025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12836__A _12836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11304__S0 _11158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17573__S _17573_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09916_ _15978_/C _12863_/B vssd1 vssd1 vccd1 vccd1 _11581_/A sky130_fd_sc_hd__nand2_2
XFILLER_59_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20036_ _20036_/CLK _20036_/D vssd1 vssd1 vccd1 vccd1 _20036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _09847_/A vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__buf_4
XFILLER_100_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11915__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09778_ _10162_/A vssd1 vssd1 vccd1 vccd1 _09779_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13437__A1 _18674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11870_/A vssd1 vssd1 vccd1 vccd1 _11740_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11671_/A vssd1 vssd1 vccd1 vccd1 _11772_/A sky130_fd_sc_hd__buf_2
XFILLER_42_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13410_ _18892_/Q vssd1 vssd1 vccd1 vccd1 _13714_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10622_ _11486_/S vssd1 vssd1 vccd1 vccd1 _10750_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_139_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14390_ _14390_/A _14390_/B vssd1 vssd1 vccd1 vccd1 _14390_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12412__A2 _12389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ input15/X _13340_/X _13319_/X vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _10553_/A _10553_/B vssd1 vssd1 vccd1 vccd1 _10553_/X sky130_fd_sc_hd__or2_1
XFILLER_167_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16652__S _16652_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16060_ _16076_/S vssd1 vssd1 vccd1 vccd1 _16073_/S sky130_fd_sc_hd__buf_2
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15362__A1 _18848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ _18809_/Q _13269_/X _12984_/X _18776_/Q _13271_/X vssd1 vssd1 vccd1 vccd1
+ _13272_/X sky130_fd_sc_hd__a221o_2
X_10484_ _10484_/A _10484_/B vssd1 vssd1 vccd1 vccd1 _10484_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15011_ _14948_/X _14933_/X _15023_/S vssd1 vssd1 vccd1 vccd1 _15011_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12176__B2 _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ _18526_/Q vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13577__A _19003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17049__A _17049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11384__C1 _19526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ _12154_/A vssd1 vssd1 vccd1 vccd1 _12154_/X sky130_fd_sc_hd__buf_2
XFILLER_123_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11105_ _11158_/S _19231_/Q vssd1 vssd1 vccd1 vccd1 _11105_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19750_ _19842_/CLK _19750_/D vssd1 vssd1 vccd1 vccd1 _19750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16962_ _16358_/X _19439_/Q _16964_/S vssd1 vssd1 vccd1 vccd1 _16963_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12085_ _12085_/A _12827_/B vssd1 vssd1 vccd1 vccd1 _12085_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10034__S0 _10277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18701_ _19912_/CLK _18701_/D vssd1 vssd1 vccd1 vccd1 _18701_/Q sky130_fd_sc_hd__dfxtp_1
X_11036_ _11149_/A _11036_/B vssd1 vssd1 vccd1 vccd1 _11036_/Y sky130_fd_sc_hd__nor2_1
X_15913_ _12082_/X _11223_/X _15916_/A vssd1 vssd1 vccd1 vccd1 _15913_/X sky130_fd_sc_hd__mux2_1
X_16893_ _16893_/A vssd1 vssd1 vccd1 vccd1 _19408_/D sky130_fd_sc_hd__clkbuf_1
X_19681_ _19940_/CLK _19681_/D vssd1 vssd1 vccd1 vccd1 _19681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18632_ _19683_/CLK _18632_/D vssd1 vssd1 vccd1 vccd1 _18632_/Q sky130_fd_sc_hd__dfxtp_1
X_15844_ _09458_/A _15842_/X _15843_/X input40/X vssd1 vssd1 vccd1 vccd1 _17201_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14201__A _14239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15775_ _15775_/A _15775_/B vssd1 vssd1 vccd1 vccd1 _15775_/X sky130_fd_sc_hd__or2_1
X_18563_ _19909_/CLK _18563_/D vssd1 vssd1 vccd1 vccd1 _18563_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _18650_/Q vssd1 vssd1 vccd1 vccd1 _14278_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14726_/A vssd1 vssd1 vccd1 vccd1 _18813_/D sky130_fd_sc_hd__clkbuf_1
X_17514_ _19663_/Q vssd1 vssd1 vccd1 vccd1 _17515_/A sky130_fd_sc_hd__clkbuf_1
X_11938_ _09197_/B _09188_/A _09190_/X _09206_/Y vssd1 vssd1 vccd1 vccd1 _11940_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18494_ _19985_/CLK _18494_/D vssd1 vssd1 vccd1 vccd1 _18494_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _17445_/A vssd1 vssd1 vccd1 vccd1 _19630_/D sky130_fd_sc_hd__clkbuf_1
X_14657_ _14663_/A _14657_/B vssd1 vssd1 vccd1 vccd1 _14658_/A sky130_fd_sc_hd__and2_1
X_11869_ _11869_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _11869_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__15050__A0 _09425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ _13608_/A vssd1 vssd1 vccd1 vccd1 _18466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17376_ _19600_/Q _17023_/X _17376_/S vssd1 vssd1 vccd1 vccd1 _17377_/A sky130_fd_sc_hd__mux2_1
X_14588_ _12231_/A _13572_/X _14598_/S vssd1 vssd1 vccd1 vccd1 _14589_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13600__A1 _13599_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19115_ _19706_/CLK _19115_/D vssd1 vssd1 vccd1 vccd1 _19115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16327_ _16326_/X _19168_/Q _16330_/S vssd1 vssd1 vccd1 vccd1 _16328_/A sky130_fd_sc_hd__mux2_1
X_13539_ _13690_/A vssd1 vssd1 vccd1 vccd1 _13575_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_146_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10176__A _15974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19046_ _19581_/CLK _19046_/D vssd1 vssd1 vccd1 vccd1 _19046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16258_ _13202_/X _19142_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _16259_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15209_ _15366_/A vssd1 vssd1 vccd1 vccd1 _15209_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14561__C1 _11717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16189_ _13238_/X _19112_/Q _16195_/S vssd1 vssd1 vccd1 vccd1 _16190_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_44_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19948_ _19948_/CLK _19948_/D vssd1 vssd1 vccd1 vccd1 _19948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14864__A0 _15270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _09701_/A vssd1 vssd1 vccd1 vccd1 _09702_/A sky130_fd_sc_hd__buf_4
XFILLER_67_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19879_ _19880_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 _19879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15408__A2 _15410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ _09933_/A vssd1 vssd1 vccd1 vccd1 _09868_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11735__A _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09563_ _09563_/A vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__buf_2
XFILLER_71_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09494_ _11951_/A _11925_/B _09436_/C vssd1 vssd1 vccd1 vccd1 _09495_/A sky130_fd_sc_hd__or3b_4
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11850__B1 _11843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16472__S _16472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__A _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15344__A1 _12390_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10814__A _18845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18399__S _18407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13107__B1 _13104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11118__C1 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18046__A0 _18838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20019_ _20021_/CLK _20019_/D vssd1 vssd1 vccd1 vccd1 _20019_/Q sky130_fd_sc_hd__dfxtp_1
X_12910_ _18937_/Q _17098_/B vssd1 vssd1 vccd1 vccd1 _14225_/D sky130_fd_sc_hd__or2_4
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13890_ _14385_/A vssd1 vssd1 vccd1 vccd1 _13890_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12841_ _12841_/A _12844_/B vssd1 vssd1 vccd1 vccd1 _12841_/Y sky130_fd_sc_hd__nor2_2
XFILLER_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13860__A _16836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15405_/X _15558_/X _15559_/X _14826_/A _12812_/Y vssd1 vssd1 vccd1 vccd1
+ _15560_/X sky130_fd_sc_hd__a32o_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12338_/A _12770_/X _12771_/Y vssd1 vssd1 vccd1 vccd1 _12772_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14510_/B _14510_/C _18737_/Q vssd1 vssd1 vccd1 vccd1 _14512_/C sky130_fd_sc_hd__a21oi_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11831_/A vssd1 vssd1 vccd1 vccd1 _11723_/X sky130_fd_sc_hd__buf_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _15491_/A _15491_/B vssd1 vssd1 vccd1 vccd1 _15491_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17125_/X _19535_/Q _17232_/S vssd1 vssd1 vccd1 vccd1 _17231_/A sky130_fd_sc_hd__mux2_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _18708_/Q _14440_/C _14441_/Y vssd1 vssd1 vccd1 vccd1 _18708_/D sky130_fd_sc_hd__o21a_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11529_/A _11530_/X _11657_/A _11655_/A vssd1 vssd1 vccd1 vccd1 _11657_/B
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__15583__A1 _18906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17161_ _17160_/X _19509_/Q _17161_/S vssd1 vssd1 vccd1 vccd1 _17162_/A sky130_fd_sc_hd__mux2_1
X_10605_ _20025_/Q _19863_/Q _19272_/Q _19042_/Q _10724_/S _10654_/A vssd1 vssd1 vccd1
+ vccd1 _10606_/B sky130_fd_sc_hd__mux4_1
XFILLER_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14373_ _18687_/Q _18686_/Q _14373_/C _14373_/D vssd1 vssd1 vccd1 vccd1 _14381_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__16382__S _16394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11585_ _11635_/A _11634_/A _11634_/B _12856_/B _10104_/A vssd1 vssd1 vccd1 vccd1
+ _11585_/X sky130_fd_sc_hd__a32o_1
XFILLER_10_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16112_ _16112_/A vssd1 vssd1 vccd1 vccd1 _19078_/D sky130_fd_sc_hd__clkbuf_1
X_13324_ _13323_/X _18445_/Q _13366_/S vssd1 vssd1 vccd1 vccd1 _13325_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09785__A _09903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _10382_/A _10527_/Y _10531_/Y _10535_/Y _09806_/A vssd1 vssd1 vccd1 vccd1
+ _10536_/X sky130_fd_sc_hd__o311a_1
X_17092_ _17092_/A vssd1 vssd1 vccd1 vccd1 _19483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16043_ _16043_/A vssd1 vssd1 vccd1 vccd1 _19050_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14543__C1 _14540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13255_ _13256_/B _13267_/C vssd1 vssd1 vccd1 vccd1 _13255_/Y sky130_fd_sc_hd__nor2_1
X_10467_ _19674_/Q _19440_/Q _18505_/Q _19770_/Q _09729_/A _10223_/A vssd1 vssd1 vccd1
+ vccd1 _10468_/B sky130_fd_sc_hd__mux4_1
XFILLER_136_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12206_ _12658_/A _12834_/A _12260_/C _18989_/Q vssd1 vssd1 vccd1 vccd1 _12263_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13186_ _13224_/C _13186_/B vssd1 vssd1 vccd1 vccd1 _13186_/Y sky130_fd_sc_hd__nor2_1
X_10398_ _10398_/A vssd1 vssd1 vccd1 vccd1 _10400_/A sky130_fd_sc_hd__buf_2
XANTENNA__10443__B _12851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19802_ _20028_/CLK _19802_/D vssd1 vssd1 vccd1 vccd1 _19802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12137_ _12165_/A _12168_/S _12135_/X _12136_/Y _12188_/A vssd1 vssd1 vccd1 vccd1
+ _12137_/Y sky130_fd_sc_hd__a311oi_4
XFILLER_151_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17994_ _19864_/Q _17049_/X _17998_/S vssd1 vssd1 vccd1 vccd1 _17995_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11109__C1 _11108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18037__B1 _16069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19733_ _20023_/CLK _19733_/D vssd1 vssd1 vccd1 vccd1 _19733_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14310__A2 _14317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16945_ _16332_/X _19431_/Q _16953_/S vssd1 vssd1 vccd1 vccd1 _16946_/A sky130_fd_sc_hd__mux2_1
X_12068_ _09361_/X _12161_/B _12067_/X _12062_/A vssd1 vssd1 vccd1 vccd1 _12069_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10558__S1 _10492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _11019_/A vssd1 vssd1 vccd1 vccd1 _11388_/A sky130_fd_sc_hd__clkbuf_2
X_19664_ _19664_/CLK _19664_/D vssd1 vssd1 vccd1 vccd1 _19664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16876_ _16876_/A vssd1 vssd1 vccd1 vccd1 _19400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16063__A2 _14554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18615_ _18745_/CLK _18615_/D vssd1 vssd1 vccd1 vccd1 _18615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15827_ _18971_/Q _15816_/X _15820_/X input35/X vssd1 vssd1 vccd1 vccd1 _15828_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19595_ _19948_/CLK _19595_/D vssd1 vssd1 vccd1 vccd1 _19595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15758_ _15758_/A _15773_/B vssd1 vssd1 vccd1 vccd1 _15758_/Y sky130_fd_sc_hd__nand2_1
X_18546_ _18547_/CLK _18546_/D vssd1 vssd1 vccd1 vccd1 _18546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14709_ _14709_/A vssd1 vssd1 vccd1 vccd1 _18805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18477_ _18547_/CLK _18477_/D vssd1 vssd1 vccd1 vccd1 _18477_/Q sky130_fd_sc_hd__dfxtp_2
X_15689_ _15689_/A vssd1 vssd1 vccd1 vccd1 _18921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10730__S1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17428_ _17496_/S vssd1 vssd1 vccd1 vccd1 _17437_/S sky130_fd_sc_hd__buf_2
XFILLER_165_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17359_ _19592_/Q _16998_/X _17365_/S vssd1 vssd1 vccd1 vccd1 _17360_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11060__A1 _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19029_ _20012_/CLK _19029_/D vssd1 vssd1 vccd1 vccd1 _19029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18012__S _18020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09615_ _20039_/Q _19877_/Q _19286_/Q _19056_/Q _09598_/X _09614_/X vssd1 vssd1 vccd1
+ vccd1 _09616_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10874__A1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09546_ _09546_/A vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__buf_4
XFILLER_43_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_0_0_clock_A clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ _13439_/A _09433_/X _09476_/X vssd1 vssd1 vccd1 vccd1 _19488_/D sky130_fd_sc_hd__o21a_1
XFILLER_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_192_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19946_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13040__A2 _12906_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11051__A1 _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11370_ _11045_/X _11367_/X _11369_/X vssd1 vssd1 vccd1 vccd1 _11370_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10321_ _19342_/Q _19613_/Q _19837_/Q _19581_/Q _10319_/X _10320_/X vssd1 vssd1 vccd1
+ vccd1 _10321_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ input29/X _12906_/X _13039_/X _12874_/X vssd1 vssd1 vccd1 vccd1 _17014_/A
+ sky130_fd_sc_hd__a22o_4
X_10252_ _10054_/X _10251_/X _10064_/A vssd1 vssd1 vccd1 vccd1 _10252_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09694__A2_N _09540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10183_ _19378_/Q _19713_/Q _10314_/S vssd1 vssd1 vccd1 vccd1 _10183_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_130_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18926_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input39_A io_ibus_inst[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ _15099_/A vssd1 vssd1 vccd1 vccd1 _14991_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13066__S _13116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16730_ _19336_/Q _13810_/X _16736_/S vssd1 vssd1 vccd1 vccd1 _16731_/A sky130_fd_sc_hd__mux2_1
X_13942_ _13945_/B _13945_/C _11884_/X vssd1 vssd1 vccd1 vccd1 _13942_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16661_ _16358_/X _19306_/Q _16663_/S vssd1 vssd1 vccd1 vccd1 _16662_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_145_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19883_/CLK sky130_fd_sc_hd__clkbuf_16
X_13873_ _12139_/A _12139_/B _13870_/X vssd1 vssd1 vccd1 vccd1 _18523_/D sky130_fd_sc_hd__a21o_1
XFILLER_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18400_ _18400_/A vssd1 vssd1 vccd1 vccd1 _20029_/D sky130_fd_sc_hd__clkbuf_1
X_15612_ _15612_/A vssd1 vssd1 vccd1 vccd1 _18887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13590__A _13660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17062__A _17062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ _12824_/A vssd1 vssd1 vccd1 vccd1 _12824_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16592_ _16592_/A vssd1 vssd1 vccd1 vccd1 _19275_/D sky130_fd_sc_hd__clkbuf_1
X_19380_ _19747_/CLK _19380_/D vssd1 vssd1 vccd1 vccd1 _19380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12918__B _12918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18331_ _17707_/X _19999_/Q _18335_/S vssd1 vssd1 vccd1 vccd1 _18332_/A sky130_fd_sc_hd__mux2_1
X_15543_ _15305_/A _15538_/Y _15542_/Y vssd1 vssd1 vccd1 vccd1 _15544_/C sky130_fd_sc_hd__a21oi_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _12755_/A vssd1 vssd1 vccd1 vccd1 _15531_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10719__A _10719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18262_ _18262_/A vssd1 vssd1 vccd1 vccd1 _19968_/D sky130_fd_sc_hd__clkbuf_1
X_11706_ _11706_/A vssd1 vssd1 vccd1 vccd1 _14672_/A sky130_fd_sc_hd__buf_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15474_ _15474_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15474_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _15498_/A _12686_/B vssd1 vssd1 vccd1 vccd1 _12689_/A sky130_fd_sc_hd__xor2_4
XANTENNA__13567__B1 _13566_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17213_ _17097_/X _19527_/Q _17221_/S vssd1 vssd1 vccd1 vccd1 _17214_/A sky130_fd_sc_hd__mux2_1
X_14425_ _18702_/Q _14420_/C _14424_/Y vssd1 vssd1 vccd1 vccd1 _18702_/D sky130_fd_sc_hd__o21a_1
X_18193_ _18193_/A vssd1 vssd1 vccd1 vccd1 _18202_/S sky130_fd_sc_hd__buf_4
X_11637_ _11524_/A _11634_/A _11634_/B _10106_/Y vssd1 vssd1 vccd1 vccd1 _11647_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12934__A _12934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17144_ _17681_/A vssd1 vssd1 vccd1 vccd1 _17144_/X sky130_fd_sc_hd__buf_2
X_14356_ _14356_/A _14356_/B _14356_/C vssd1 vssd1 vccd1 vccd1 _18683_/D sky130_fd_sc_hd__nor3_1
X_11568_ _19686_/Q _19452_/Q _18517_/Q _19782_/Q _11553_/X _11554_/A vssd1 vssd1 vccd1
+ vccd1 _11568_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10396__A3 _10395_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13307_ _13307_/A vssd1 vssd1 vccd1 vccd1 _13307_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10519_ _20027_/Q _19865_/Q _19274_/Q _19044_/Q _10216_/A _10218_/A vssd1 vssd1 vccd1
+ vccd1 _10520_/B sky130_fd_sc_hd__mux4_1
X_17075_ _17075_/A vssd1 vssd1 vccd1 vccd1 _17088_/S sky130_fd_sc_hd__buf_4
XFILLER_7_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14287_ _18662_/Q _18661_/Q _18660_/Q _14287_/D vssd1 vssd1 vccd1 vccd1 _14297_/D
+ sky130_fd_sc_hd__and4_1
X_11499_ _19926_/Q _19540_/Q _19990_/Q _19109_/Q _11488_/S _10856_/X vssd1 vssd1 vccd1
+ vccd1 _11500_/B sky130_fd_sc_hd__mux4_1
X_16026_ _16026_/A vssd1 vssd1 vccd1 vccd1 _19042_/D sky130_fd_sc_hd__clkbuf_1
X_13238_ _17688_/A vssd1 vssd1 vccd1 vccd1 _13238_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10779__S1 _10048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13765__A _17001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13169_ _18727_/Q vssd1 vssd1 vccd1 vccd1 _14485_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17977_ _17977_/A vssd1 vssd1 vccd1 vccd1 _19856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15492__B1 _15954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19716_ _20006_/CLK _19716_/D vssd1 vssd1 vccd1 vccd1 _19716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15980__A _15982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16928_ _16928_/A vssd1 vssd1 vccd1 vccd1 _19423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19647_ _20035_/CLK _19647_/D vssd1 vssd1 vccd1 vccd1 _19647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16287__S _16291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16859_ _16313_/X _19393_/Q _16859_/S vssd1 vssd1 vccd1 vccd1 _16860_/A sky130_fd_sc_hd__mux2_1
X_09400_ _14227_/A _11697_/C vssd1 vssd1 vccd1 vccd1 _09408_/B sky130_fd_sc_hd__or2_4
XFILLER_53_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10951__S1 _10624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19578_ _20028_/CLK _19578_/D vssd1 vssd1 vccd1 vccd1 _19578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09331_ _09328_/Y _18939_/Q _18827_/Q _09696_/A _09698_/C vssd1 vssd1 vccd1 vccd1
+ _09337_/B sky130_fd_sc_hd__o2111a_1
X_18529_ _18868_/CLK _18529_/D vssd1 vssd1 vccd1 vccd1 _18529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09262_ _18988_/Q vssd1 vssd1 vccd1 vccd1 _09263_/A sky130_fd_sc_hd__buf_4
XANTENNA__11281__A1 _11003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15547__B2 _12791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13558__A0 _18460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09193_ _09230_/A vssd1 vssd1 vccd1 vccd1 _09521_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18007__S _18009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12844__A _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17846__S _17854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16750__S _16758_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10219__S0 _10388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_62_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19865_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_130_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11195__A _18837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10942__S1 _10624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_166_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10870_ _19665_/Q _19431_/Q _18496_/Q _19761_/Q _10919_/S _10596_/A vssd1 vssd1 vccd1
+ vccd1 _10871_/B sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_77_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19810_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09909_/A _09528_/X _15127_/S vssd1 vssd1 vccd1 vccd1 _09530_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16925__S _16931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12839__A_N _12833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12540_ _12540_/A vssd1 vssd1 vccd1 vccd1 _15424_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13549__A0 _18459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _18535_/Q vssd1 vssd1 vccd1 vccd1 _12501_/A sky130_fd_sc_hd__buf_2
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13013__A2 _13189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16226__A _16282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14210_ _14239_/A _14210_/B vssd1 vssd1 vccd1 vccd1 _14210_/Y sky130_fd_sc_hd__nor2_1
X_11422_ _18424_/Q _19453_/Q _19490_/Q _19064_/Q _11212_/A _11077_/A vssd1 vssd1 vccd1
+ vccd1 _11422_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15190_ _15188_/X _15189_/X _15190_/S vssd1 vssd1 vccd1 vccd1 _15190_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12772__A1 _12338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14141_ _14142_/B _14142_/C _18620_/Q vssd1 vssd1 vccd1 vccd1 _14143_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__17756__S _17760_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11353_ _11344_/A _11352_/X _09772_/A vssd1 vssd1 vccd1 vccd1 _11353_/X sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_15_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19951_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10304_ _19214_/Q _19805_/Q _19967_/Q _19182_/Q _09655_/A _10185_/X vssd1 vssd1 vccd1
+ vccd1 _10305_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14072_ _14088_/A _14072_/B _14072_/C vssd1 vssd1 vccd1 vccd1 _18599_/D sky130_fd_sc_hd__nor3_1
XFILLER_141_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11284_ _18427_/Q _19456_/Q _19493_/Q _19067_/Q _11121_/S _11077_/X vssd1 vssd1 vccd1
+ vccd1 _11284_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13023_ _17652_/A vssd1 vssd1 vccd1 vccd1 _13023_/X sky130_fd_sc_hd__clkbuf_2
X_17900_ _19822_/Q _17017_/X _17904_/S vssd1 vssd1 vccd1 vccd1 _17901_/A sky130_fd_sc_hd__mux2_1
X_10235_ _10342_/A _10235_/B vssd1 vssd1 vccd1 vccd1 _10235_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18880_ _18918_/CLK _18880_/D vssd1 vssd1 vccd1 vccd1 _18880_/Q sky130_fd_sc_hd__dfxtp_1
X_17831_ _17831_/A vssd1 vssd1 vccd1 vccd1 _19791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10166_ _19379_/Q _19714_/Q _10166_/S vssd1 vssd1 vccd1 vccd1 _10166_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output145_A _12352_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17762_ _17808_/S vssd1 vssd1 vccd1 vccd1 _17771_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_94_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10097_ _09940_/A _10094_/X _10096_/X vssd1 vssd1 vccd1 vccd1 _10097_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14974_ _15945_/A vssd1 vssd1 vccd1 vccd1 _15940_/A sky130_fd_sc_hd__clkbuf_2
X_19501_ _19637_/CLK _19501_/D vssd1 vssd1 vccd1 vccd1 _19501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16713_ _16713_/A vssd1 vssd1 vccd1 vccd1 _19328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13925_ _13946_/A _13925_/B _13925_/C vssd1 vssd1 vccd1 vccd1 _18550_/D sky130_fd_sc_hd__nor3_1
XFILLER_48_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17693_ _17693_/A vssd1 vssd1 vccd1 vccd1 _19736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19432_ _19861_/CLK _19432_/D vssd1 vssd1 vccd1 vccd1 _19432_/Q sky130_fd_sc_hd__dfxtp_1
X_16644_ _16332_/X _19298_/Q _16652_/S vssd1 vssd1 vccd1 vccd1 _16645_/A sky130_fd_sc_hd__mux2_1
X_13856_ _13856_/A vssd1 vssd1 vccd1 vccd1 _18516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ _15553_/B _12807_/B vssd1 vssd1 vccd1 vccd1 _14970_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19363_ _20023_/CLK _19363_/D vssd1 vssd1 vccd1 vccd1 _19363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16575_ _16575_/A vssd1 vssd1 vccd1 vccd1 _19267_/D sky130_fd_sc_hd__clkbuf_1
X_13787_ _17023_/A vssd1 vssd1 vccd1 vccd1 _13787_/X sky130_fd_sc_hd__clkbuf_2
X_10999_ _09683_/A _10989_/X _10993_/Y _10998_/Y _09873_/A vssd1 vssd1 vccd1 vccd1
+ _10999_/X sky130_fd_sc_hd__o221a_1
X_18314_ _18314_/A vssd1 vssd1 vccd1 vccd1 _19991_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12738_/A vssd1 vssd1 vccd1 vccd1 _15520_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15526_ _18861_/Q _15457_/X _15525_/X vssd1 vssd1 vccd1 vccd1 _18861_/D sky130_fd_sc_hd__o21a_1
XFILLER_124_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ _19757_/CLK _19294_/D vssd1 vssd1 vccd1 vccd1 _19294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18245_ _18245_/A vssd1 vssd1 vccd1 vccd1 _19960_/D sky130_fd_sc_hd__clkbuf_1
X_15457_ _15457_/A vssd1 vssd1 vccd1 vccd1 _15457_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12669_ _12729_/A _12645_/B _12640_/A vssd1 vssd1 vccd1 vccd1 _12670_/B sky130_fd_sc_hd__a21bo_1
XFILLER_129_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12664__A _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14408_ _14411_/C _14409_/C _18698_/Q vssd1 vssd1 vccd1 vccd1 _14410_/B sky130_fd_sc_hd__a21oi_1
X_18176_ _17691_/X _19930_/Q _18180_/S vssd1 vssd1 vccd1 vccd1 _18177_/A sky130_fd_sc_hd__mux2_1
X_15388_ _15365_/X _15331_/X _15387_/X _15324_/X vssd1 vssd1 vccd1 vccd1 _15388_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_116_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17666__S _17666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17127_ _17127_/A vssd1 vssd1 vccd1 vccd1 _19498_/D sky130_fd_sc_hd__clkbuf_1
X_14339_ _14373_/C vssd1 vssd1 vccd1 vccd1 _14364_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ _17058_/A vssd1 vssd1 vccd1 vccd1 _17058_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16009_ _13115_/X _19035_/Q _16009_/S vssd1 vssd1 vccd1 vccd1 _16010_/A sky130_fd_sc_hd__mux2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09880_/A vssd1 vssd1 vccd1 vccd1 _09881_/A sky130_fd_sc_hd__clkbuf_4
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11462__B _11462_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16745__S _16747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09314_ _09501_/B _09310_/C _09276_/X _09516_/B vssd1 vssd1 vccd1 vccd1 _14822_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10688__S0 _10691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09245_ _09245_/A vssd1 vssd1 vccd1 vccd1 _09309_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_166_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09176_ _09282_/B vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12754__A1 _14750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13951__B1 _11884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17576__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17142__A0 _17141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16480__S _16486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09883__A _09883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_92_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12506__A1 _12338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__A _11918_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10822__A _10822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10020_ _10749_/S vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__buf_2
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18200__S _18202_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11971_ _11971_/A _11971_/B vssd1 vssd1 vccd1 vccd1 _11971_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_57_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13710_ _13656_/X _13708_/X _13709_/Y _13660_/X _19020_/Q vssd1 vssd1 vccd1 vccd1
+ _13710_/X sky130_fd_sc_hd__a32o_2
X_10922_ _10664_/A _10921_/X _10929_/A vssd1 vssd1 vccd1 vccd1 _10922_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14690_ _18797_/Q _14548_/A _14694_/S vssd1 vssd1 vccd1 vccd1 _14691_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15759__A1 _09467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ _13641_/A vssd1 vssd1 vccd1 vccd1 _18470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10853_ _11015_/A vssd1 vssd1 vccd1 vccd1 _10854_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16655__S _16663_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16360_/A vssd1 vssd1 vccd1 vccd1 _19178_/D sky130_fd_sc_hd__clkbuf_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11245__A1 _09774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ _13528_/X _13570_/X _13571_/Y _13532_/X _19002_/Q vssd1 vssd1 vccd1 vccd1
+ _13572_/X sky130_fd_sc_hd__a32o_4
X_10784_ _10784_/A vssd1 vssd1 vccd1 vccd1 _10784_/Y sky130_fd_sc_hd__inv_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _12335_/Y _15279_/X _15310_/X _15275_/X vssd1 vssd1 vccd1 vccd1 _15311_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12993__A1 _14355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12523_ _18537_/Q _12523_/B vssd1 vssd1 vccd1 vccd1 _12525_/A sky130_fd_sc_hd__nor2_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _13463_/X _19157_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _16292_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12915__C _16150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18030_ _18115_/A vssd1 vssd1 vccd1 vccd1 _18134_/S sky130_fd_sc_hd__clkbuf_2
X_15242_ _18841_/Q _09433_/X _15241_/X vssd1 vssd1 vccd1 vccd1 _18841_/D sky130_fd_sc_hd__o21a_1
X_12454_ _12446_/A _12415_/X _12450_/Y _12453_/X vssd1 vssd1 vccd1 vccd1 _12454_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15931__A1 _19002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17486__S _17492_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ _11440_/A _11402_/X _11404_/X _09788_/A vssd1 vssd1 vccd1 vccd1 _11405_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13942__B1 _11884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15173_ _15093_/X _15163_/X _15172_/X _15048_/X _12124_/X vssd1 vssd1 vccd1 vccd1
+ _15173_/X sky130_fd_sc_hd__a32o_1
XFILLER_165_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12385_ _12385_/A _14879_/A vssd1 vssd1 vccd1 vccd1 _12386_/B sky130_fd_sc_hd__or2_1
XANTENNA__18171__A _18193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14124_ _18614_/Q _14124_/B _14529_/B vssd1 vssd1 vccd1 vccd1 _14125_/C sky130_fd_sc_hd__and3_1
X_11336_ _11131_/A _11333_/X _11335_/X _11058_/A vssd1 vssd1 vccd1 vccd1 _11336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19981_ _19981_/CLK _19981_/D vssd1 vssd1 vccd1 vccd1 _19981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14055_ _14245_/A vssd1 vssd1 vccd1 vccd1 _14090_/A sky130_fd_sc_hd__clkbuf_2
X_18932_ _18967_/CLK _18932_/D vssd1 vssd1 vccd1 vccd1 _18932_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11828__A _19005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ _09550_/A _11255_/X _11266_/X vssd1 vssd1 vccd1 vccd1 _11267_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13006_ _18555_/Q vssd1 vssd1 vccd1 vccd1 _13945_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10218_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10223_/A sky130_fd_sc_hd__buf_4
XFILLER_140_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18863_ _18911_/CLK _18863_/D vssd1 vssd1 vccd1 vccd1 _18863_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11198_ _19228_/Q _19723_/Q _11367_/S vssd1 vssd1 vccd1 vccd1 _11199_/B sky130_fd_sc_hd__mux2_1
XFILLER_67_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17814_ _17814_/A vssd1 vssd1 vccd1 vccd1 _19783_/D sky130_fd_sc_hd__clkbuf_1
X_10149_ _10149_/A vssd1 vssd1 vccd1 vccd1 _10376_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18794_ _19062_/CLK _18794_/D vssd1 vssd1 vccd1 vccd1 _18794_/Q sky130_fd_sc_hd__dfxtp_1
X_17745_ _17643_/X _19753_/Q _17749_/S vssd1 vssd1 vccd1 vccd1 _17746_/A sky130_fd_sc_hd__mux2_1
X_14957_ _14955_/X _14956_/X _14957_/S vssd1 vssd1 vccd1 vccd1 _14957_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12659__A _12753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _18547_/Q _12820_/A _12772_/Y _12775_/Y _13904_/X vssd1 vssd1 vccd1 vccd1
+ _18547_/D sky130_fd_sc_hd__o221a_1
X_17676_ _17675_/X _19731_/Q _17682_/S vssd1 vssd1 vccd1 vccd1 _17677_/A sky130_fd_sc_hd__mux2_1
X_14888_ _14884_/X _14887_/X _14916_/S vssd1 vssd1 vccd1 vccd1 _14888_/X sky130_fd_sc_hd__mux2_1
X_19415_ _19942_/CLK _19415_/D vssd1 vssd1 vccd1 vccd1 _19415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16627_ _16627_/A vssd1 vssd1 vccd1 vccd1 _19290_/D sky130_fd_sc_hd__clkbuf_1
X_13839_ _13839_/A vssd1 vssd1 vccd1 vccd1 _13852_/S sky130_fd_sc_hd__buf_4
XANTENNA__16565__S _16569_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19346_ _19942_/CLK _19346_/D vssd1 vssd1 vccd1 vccd1 _19346_/Q sky130_fd_sc_hd__dfxtp_1
X_16558_ _19260_/Q _13771_/X _16558_/S vssd1 vssd1 vccd1 vccd1 _16559_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11331__S1 _11322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15509_ _15509_/A _15509_/B vssd1 vssd1 vccd1 vccd1 _15509_/Y sky130_fd_sc_hd__nor2_1
X_19277_ _19836_/CLK _19277_/D vssd1 vssd1 vccd1 vccd1 _19277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16489_ _19229_/Q _13774_/X _16497_/S vssd1 vssd1 vccd1 vccd1 _16490_/A sky130_fd_sc_hd__mux2_1
X_18228_ _19953_/Q _17662_/A _18230_/S vssd1 vssd1 vccd1 vccd1 _18229_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17396__S _17398_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13933__B1 _11884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18159_ _18159_/A vssd1 vssd1 vccd1 vccd1 _19922_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_114_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18081__A _18115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10842__S0 _10797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12841__B _12844_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09932_ _19220_/Q _19811_/Q _19973_/Q _19188_/Q _09659_/S _09647_/A vssd1 vssd1 vccd1
+ vccd1 _09933_/B sky130_fd_sc_hd__mux4_1
XFILLER_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15150__A2 _15053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11398__S1 _11357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09863_ _19942_/Q _19556_/Q _20006_/Q _19125_/Q _09598_/X _09851_/A vssd1 vssd1 vccd1
+ vccd1 _09864_/B sky130_fd_sc_hd__mux4_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11457__B _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13953__A _14745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09794_/A vssd1 vssd1 vccd1 vccd1 _10579_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18020__S _18020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11473__A _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_39_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10817__A _15938_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09228_ _18961_/Q vssd1 vssd1 vccd1 vccd1 _09481_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__14177__B1 _14160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15913__A1 _11223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12727__A1 _12170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10833__S0 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ _12347_/A vssd1 vssd1 vccd1 vccd1 _12170_/X sky130_fd_sc_hd__buf_2
XFILLER_108_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11121_ _19230_/Q _19725_/Q _11121_/S vssd1 vssd1 vccd1 vccd1 _11122_/B sky130_fd_sc_hd__mux2_1
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09356__B1 _13340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11052_ _19327_/Q _19598_/Q _19822_/Q _19566_/Q _10977_/S _11045_/X vssd1 vssd1 vccd1
+ vccd1 _11052_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14959__A _15103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ _10573_/S vssd1 vssd1 vccd1 vccd1 _10279_/A sky130_fd_sc_hd__buf_4
XFILLER_103_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13863__A _13910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18091__A1 _11764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15860_ _09467_/X _15856_/X _15788_/X input46/X vssd1 vssd1 vccd1 vccd1 _16837_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input21_A io_dbus_rdata[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14101__B1 _14100_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ _14811_/A _14811_/B _14811_/C vssd1 vssd1 vccd1 vccd1 _14814_/B sky130_fd_sc_hd__or3_1
XFILLER_18_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15791_ _15833_/A _15791_/B vssd1 vssd1 vccd1 vccd1 _15792_/A sky130_fd_sc_hd__or2_1
XFILLER_123_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13455__A2 _13081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17530_ _19671_/Q vssd1 vssd1 vccd1 vccd1 _17531_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12663__A0 _15970_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14742_ _18821_/Q _13750_/B _14742_/S vssd1 vssd1 vccd1 vccd1 _14743_/A sky130_fd_sc_hd__mux2_1
X_11954_ _09198_/A _09309_/A _14761_/C vssd1 vssd1 vccd1 vccd1 _14818_/A sky130_fd_sc_hd__a21o_1
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10905_ _10905_/A _10905_/B vssd1 vssd1 vccd1 vccd1 _10905_/X sky130_fd_sc_hd__or2_1
XFILLER_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17461_ _17483_/A vssd1 vssd1 vccd1 vccd1 _17470_/S sky130_fd_sc_hd__buf_4
XFILLER_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14673_ _14729_/A vssd1 vssd1 vccd1 vccd1 _14742_/S sky130_fd_sc_hd__buf_2
XANTENNA__16385__S _16394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11885_ _15765_/A vssd1 vssd1 vccd1 vccd1 _15732_/B sky130_fd_sc_hd__buf_2
XFILLER_45_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output108_A _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19200_ _19824_/CLK _19200_/D vssd1 vssd1 vccd1 vccd1 _19200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16412_ _16412_/A vssd1 vssd1 vccd1 vccd1 _19195_/D sky130_fd_sc_hd__clkbuf_1
X_13624_ _13690_/A vssd1 vssd1 vccd1 vccd1 _13670_/S sky130_fd_sc_hd__buf_2
X_10836_ _10836_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _10836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17392_ _19607_/Q _17046_/X _17398_/S vssd1 vssd1 vccd1 vccd1 _17393_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12926__B _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19131_ _19981_/CLK _19131_/D vssd1 vssd1 vccd1 vccd1 _19131_/Q sky130_fd_sc_hd__dfxtp_1
X_16343_ _16342_/X _19173_/Q _16346_/S vssd1 vssd1 vccd1 vccd1 _16344_/A sky130_fd_sc_hd__mux2_1
X_13555_ _13554_/A _13554_/C _13046_/A vssd1 vssd1 vccd1 vccd1 _13556_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11830__B _19005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10767_ _10654_/A _10764_/X _10766_/X vssd1 vssd1 vccd1 vccd1 _10767_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ _12338_/X _12504_/X _12505_/Y vssd1 vssd1 vccd1 vccd1 _12506_/Y sky130_fd_sc_hd__a21oi_1
X_16274_ _13323_/X _19149_/Q _16280_/S vssd1 vssd1 vccd1 vccd1 _16275_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19062_ _19062_/CLK _19062_/D vssd1 vssd1 vccd1 vccd1 _19062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13486_ _18896_/Q _13486_/B vssd1 vssd1 vccd1 vccd1 _13486_/X sky130_fd_sc_hd__or2_1
XFILLER_157_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10698_ _10579_/X _10693_/X _10695_/Y _10697_/Y _09805_/A vssd1 vssd1 vccd1 vccd1
+ _10698_/X sky130_fd_sc_hd__o221a_1
X_18013_ _18013_/A vssd1 vssd1 vccd1 vccd1 _19872_/D sky130_fd_sc_hd__clkbuf_1
X_15225_ _18840_/Q _09433_/X _15224_/X vssd1 vssd1 vccd1 vccd1 _18840_/D sky130_fd_sc_hd__o21a_1
XFILLER_157_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12437_ _12437_/A _12467_/A vssd1 vssd1 vccd1 vccd1 _12442_/A sky130_fd_sc_hd__xor2_4
XFILLER_138_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15156_ _15517_/A _15160_/A vssd1 vssd1 vccd1 vccd1 _15156_/X sky130_fd_sc_hd__or2_1
X_12368_ _12368_/A _12416_/D vssd1 vssd1 vccd1 vccd1 _12392_/B sky130_fd_sc_hd__nand2_1
XFILLER_154_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14107_ _14143_/A _14107_/B _14107_/C vssd1 vssd1 vccd1 vccd1 _18611_/D sky130_fd_sc_hd__nor3_1
XANTENNA__17944__S _17948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11319_ _19354_/Q _19689_/Q _11410_/S vssd1 vssd1 vccd1 vccd1 _11320_/B sky130_fd_sc_hd__mux2_1
X_19964_ _20028_/CLK _19964_/D vssd1 vssd1 vccd1 vccd1 _19964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15087_ _15413_/A vssd1 vssd1 vccd1 vccd1 _15491_/A sky130_fd_sc_hd__clkbuf_2
X_12299_ _12299_/A _15270_/B vssd1 vssd1 vccd1 vccd1 _12299_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14038_ _14046_/A _14042_/C vssd1 vssd1 vccd1 vccd1 _14038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18915_ _19350_/CLK _18915_/D vssd1 vssd1 vccd1 vccd1 _18915_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15972__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19895_ _19912_/CLK _19895_/D vssd1 vssd1 vccd1 vccd1 _19895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17245__A _17267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18846_ _19855_/CLK _18846_/D vssd1 vssd1 vccd1 vccd1 _18846_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__09993__S1 _09637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18777_ _19900_/CLK _18777_/D vssd1 vssd1 vccd1 vccd1 _18777_/Q sky130_fd_sc_hd__dfxtp_1
X_15989_ _16057_/S vssd1 vssd1 vccd1 vccd1 _15998_/S sky130_fd_sc_hd__buf_4
XFILLER_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13446__A2 _13340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11293__A _11293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17728_ _17728_/A vssd1 vssd1 vccd1 vccd1 _19747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17593__A0 _17141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16295__S _16295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17659_ _17659_/A vssd1 vssd1 vccd1 vccd1 _17659_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13749__A3 _09341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__S1 _11108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19329_ _19824_/CLK _19329_/D vssd1 vssd1 vccd1 vccd1 _19329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13948__A _13958_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12852__A _12863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17854__S _17854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10291__S1 _10283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13134__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09915_ _09884_/X _09894_/X _09908_/Y _09913_/X _09914_/Y vssd1 vssd1 vccd1 vccd1
+ _12863_/B sky130_fd_sc_hd__o32a_4
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20035_ _20035_/CLK _20035_/D vssd1 vssd1 vccd1 vccd1 _20035_/Q sky130_fd_sc_hd__dfxtp_1
X_09846_ _18976_/Q _09465_/C _10077_/A vssd1 vssd1 vccd1 vccd1 _09847_/A sky130_fd_sc_hd__o21a_1
XFILLER_112_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09777_ _09777_/A vssd1 vssd1 vccd1 vccd1 _10162_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16994__A _17075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11670_/A vssd1 vssd1 vccd1 vccd1 _14547_/A sky130_fd_sc_hd__buf_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10621_ _10907_/S vssd1 vssd1 vccd1 vccd1 _11486_/S sky130_fd_sc_hd__buf_4
XANTENNA__14019__A _14102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13340_ _13340_/A vssd1 vssd1 vccd1 vccd1 _13340_/X sky130_fd_sc_hd__clkbuf_2
X_10552_ _19930_/Q _19544_/Q _19994_/Q _19113_/Q _10319_/A _10497_/X vssd1 vssd1 vccd1
+ vccd1 _10553_/B sky130_fd_sc_hd__mux4_1
XFILLER_167_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13271_ _18473_/Q _11755_/X _12881_/X _18697_/Q _13270_/X vssd1 vssd1 vccd1 vccd1
+ _13271_/X sky130_fd_sc_hd__a221o_1
X_10483_ _19211_/Q _19802_/Q _19964_/Q _19179_/Q _10279_/A _10473_/X vssd1 vssd1 vccd1
+ vccd1 _10484_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15010_ _15029_/A vssd1 vssd1 vccd1 vccd1 _15023_/S sky130_fd_sc_hd__clkbuf_2
X_12222_ _12503_/A vssd1 vssd1 vccd1 vccd1 _12770_/S sky130_fd_sc_hd__buf_2
XFILLER_108_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input69_A io_irq_uart_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13577__B _13577_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12153_ _15633_/C _12153_/B _12153_/C _12153_/D vssd1 vssd1 vccd1 vccd1 _12153_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _19726_/Q vssd1 vssd1 vccd1 vccd1 _11104_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16961_ _16961_/A vssd1 vssd1 vccd1 vccd1 _19438_/D sky130_fd_sc_hd__clkbuf_1
X_12084_ hold4/A _12083_/X _12084_/S vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18700_ _19912_/CLK _18700_/D vssd1 vssd1 vccd1 vccd1 _18700_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17065__A _17065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ _19921_/Q _19535_/Q _19985_/Q _19104_/Q _10962_/X _10893_/A vssd1 vssd1 vccd1
+ vccd1 _11036_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15912_ _15912_/A vssd1 vssd1 vccd1 vccd1 _18997_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10034__S1 _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19680_ _20033_/CLK _19680_/D vssd1 vssd1 vccd1 vccd1 _19680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11231__S0 _11230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16892_ _16361_/X _19408_/Q _16892_/S vssd1 vssd1 vccd1 vccd1 _16893_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18631_ _19683_/CLK _18631_/D vssd1 vssd1 vccd1 vccd1 _18631_/Q sky130_fd_sc_hd__dfxtp_1
X_15843_ _15879_/A vssd1 vssd1 vccd1 vccd1 _15843_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14625__A1 _13661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18562_ _19909_/CLK _18562_/D vssd1 vssd1 vccd1 vccd1 _18562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _09261_/A _15765_/X _15773_/Y _15769_/X vssd1 vssd1 vccd1 vccd1 _18955_/D
+ sky130_fd_sc_hd__o211a_1
X_12986_ _12134_/B _12984_/X _12985_/X vssd1 vssd1 vccd1 vccd1 _12986_/X sky130_fd_sc_hd__a21o_1
XFILLER_91_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _17513_/A vssd1 vssd1 vccd1 vccd1 _19662_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14725_ _18813_/Q _11879_/X _14727_/S vssd1 vssd1 vccd1 vccd1 _14726_/A sky130_fd_sc_hd__mux2_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _14819_/B _11937_/B vssd1 vssd1 vccd1 vccd1 _11937_/X sky130_fd_sc_hd__and2_1
X_18493_ _19758_/CLK _18493_/D vssd1 vssd1 vccd1 vccd1 _18493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _17122_/X _19630_/Q _17448_/S vssd1 vssd1 vccd1 vccd1 _17445_/A sky130_fd_sc_hd__mux2_1
X_11868_ _12060_/B _14159_/A _11860_/B vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14656_ _18785_/Q _13727_/X _14667_/S vssd1 vssd1 vccd1 vccd1 _14657_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10819_ _19363_/Q _19698_/Q _10821_/S vssd1 vssd1 vccd1 vccd1 _10820_/B sky130_fd_sc_hd__mux2_1
X_13607_ _18466_/Q _13606_/X _13617_/S vssd1 vssd1 vccd1 vccd1 _13608_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13061__A0 _18840_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17375_ _17375_/A vssd1 vssd1 vccd1 vccd1 _19599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14587_ _14587_/A vssd1 vssd1 vccd1 vccd1 _18764_/D sky130_fd_sc_hd__clkbuf_1
X_11799_ _13747_/A _18997_/Q _11730_/A vssd1 vssd1 vccd1 vccd1 _11799_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19114_ _20027_/CLK _19114_/D vssd1 vssd1 vccd1 vccd1 _19114_/Q sky130_fd_sc_hd__dfxtp_1
X_16326_ _17662_/A vssd1 vssd1 vccd1 vccd1 _16326_/X sky130_fd_sc_hd__clkbuf_1
X_13538_ hold7/A _13536_/Y _13583_/S vssd1 vssd1 vccd1 vccd1 _13538_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10176__B _12860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19045_ _20028_/CLK _19045_/D vssd1 vssd1 vccd1 vccd1 _19045_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13768__A _17004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16257_ _16257_/A vssd1 vssd1 vccd1 vccd1 _19141_/D sky130_fd_sc_hd__clkbuf_1
X_13469_ _18820_/Q _11841_/X _11843_/X _18787_/Q _13468_/X vssd1 vssd1 vccd1 vccd1
+ _13469_/X sky130_fd_sc_hd__a221o_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15208_ _15444_/A vssd1 vssd1 vccd1 vccd1 _15236_/A sky130_fd_sc_hd__clkbuf_2
X_16188_ _16188_/A vssd1 vssd1 vccd1 vccd1 _19111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10192__A _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15139_ _15139_/A _15183_/A vssd1 vssd1 vccd1 vccd1 _15139_/X sky130_fd_sc_hd__or2_1
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14313__B1 _18670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19947_ _19947_/CLK _19947_/D vssd1 vssd1 vccd1 vccd1 _19947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _09909_/A _09697_/X _09698_/X _09699_/Y vssd1 vssd1 vccd1 vccd1 _09701_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_96_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19878_ _20040_/CLK _19878_/D vssd1 vssd1 vccd1 vccd1 _19878_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10920__A _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09631_ _10073_/A vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__buf_2
XFILLER_110_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18829_ _19880_/CLK _18829_/D vssd1 vssd1 vccd1 vccd1 _18829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09562_ _09562_/A vssd1 vssd1 vccd1 vccd1 _09563_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09920__S _09920_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10102__A1 _09809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09493_ _11941_/A _15899_/A vssd1 vssd1 vccd1 vccd1 _12084_/S sky130_fd_sc_hd__nor2_2
XFILLER_24_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12847__A _12851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12566__B _12853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17318__A0 _17147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10169__A1 _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17584__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11905__A2 _11904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18046__A1 _13546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__A _12587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11213__S0 _11212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20018_ _20018_/CLK _20018_/D vssd1 vssd1 vccd1 vccd1 _20018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09829_ _11237_/A vssd1 vssd1 vccd1 vccd1 _09830_/A sky130_fd_sc_hd__buf_2
XFILLER_59_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _12840_/A vssd1 vssd1 vccd1 vccd1 _12840_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _18483_/Q _12012_/X _13648_/A vssd1 vssd1 vccd1 vccd1 _12771_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13291__B1 _12881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11722_/A vssd1 vssd1 vccd1 vccd1 _11831_/A sky130_fd_sc_hd__clkbuf_4
X_14510_ _18737_/Q _14510_/B _14510_/C vssd1 vssd1 vccd1 vccd1 _14512_/B sky130_fd_sc_hd__and3_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15071_/X _15194_/B _15489_/X _15491_/A vssd1 vssd1 vccd1 vccd1 _15490_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17309__A0 _17135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11653_ _12003_/C _11975_/A _11650_/X vssd1 vssd1 vccd1 vccd1 _11653_/X sky130_fd_sc_hd__or3b_1
XFILLER_30_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14441_ _18708_/Q _14440_/C _14427_/X vssd1 vssd1 vccd1 vccd1 _14441_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16663__S _16663_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14972__A _15458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ _09562_/A _10599_/Y _10603_/Y _09875_/A vssd1 vssd1 vccd1 vccd1 _10604_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_11_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12397__A2 _12012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17160_ _17697_/A vssd1 vssd1 vccd1 vccd1 _17160_/X sky130_fd_sc_hd__clkbuf_2
X_14372_ _14399_/A _14372_/B _14378_/C vssd1 vssd1 vccd1 vccd1 _18687_/D sky130_fd_sc_hd__nor3_1
XFILLER_155_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11584_ _11582_/A _11526_/Y _11583_/X vssd1 vssd1 vccd1 vccd1 _11584_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_168_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13323_ _17704_/A vssd1 vssd1 vccd1 vccd1 _13323_/X sky130_fd_sc_hd__clkbuf_1
X_16111_ _13202_/X _19078_/Q _16111_/S vssd1 vssd1 vccd1 vccd1 _16112_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10535_ _10520_/A _10532_/X _10534_/X vssd1 vssd1 vccd1 vccd1 _10535_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17091_ _19483_/Q _17090_/X _17094_/S vssd1 vssd1 vccd1 vccd1 _17092_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16042_ _13365_/X _19050_/Q _16042_/S vssd1 vssd1 vccd1 vccd1 _16043_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_8_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13254_ _18883_/Q vssd1 vssd1 vccd1 vccd1 _13256_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10466_ _09849_/A _10456_/X _10465_/X _09539_/A _18852_/Q vssd1 vssd1 vccd1 vccd1
+ _15958_/C sky130_fd_sc_hd__a32o_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17494__S _17496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ _12205_/A vssd1 vssd1 vccd1 vccd1 _12205_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13185_ _13630_/A _13183_/B _12897_/X vssd1 vssd1 vccd1 vccd1 _13186_/B sky130_fd_sc_hd__o21ai_1
X_10397_ _15962_/C _12853_/B vssd1 vssd1 vccd1 vccd1 _11629_/A sky130_fd_sc_hd__or2_1
XFILLER_151_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19801_ _19864_/CLK _19801_/D vssd1 vssd1 vccd1 vccd1 _19801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12136_ _12059_/X _12135_/X _12165_/A vssd1 vssd1 vccd1 vccd1 _12136_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17993_ _17993_/A vssd1 vssd1 vccd1 vccd1 _19863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19732_ _19732_/CLK _19732_/D vssd1 vssd1 vccd1 vccd1 _19732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18037__A1 _12956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16944_ _16990_/S vssd1 vssd1 vccd1 vccd1 _16953_/S sky130_fd_sc_hd__clkbuf_4
X_12067_ _18711_/Q _12061_/A _12163_/C _12066_/Y vssd1 vssd1 vccd1 vccd1 _12067_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__11204__S0 _11063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11018_ _10962_/X _10979_/Y _11017_/Y _11157_/A vssd1 vssd1 vccd1 vccd1 _11018_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19663_ _20015_/CLK _19663_/D vssd1 vssd1 vccd1 vccd1 _19663_/Q sky130_fd_sc_hd__dfxtp_1
X_16875_ _16336_/X _19400_/Q _16881_/S vssd1 vssd1 vccd1 vccd1 _16876_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18614_ _18745_/CLK _18614_/D vssd1 vssd1 vccd1 vccd1 _18614_/Q sky130_fd_sc_hd__dfxtp_1
X_15826_ _15826_/A vssd1 vssd1 vccd1 vccd1 _18970_/D sky130_fd_sc_hd__clkbuf_1
X_19594_ _19947_/CLK _19594_/D vssd1 vssd1 vccd1 vccd1 _19594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10139__A1_N _18860_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18545_ _18547_/CLK _18545_/D vssd1 vssd1 vccd1 vccd1 _18545_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _12082_/X _15752_/X _15755_/X _15756_/X vssd1 vssd1 vccd1 vccd1 _18948_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _19488_/Q vssd1 vssd1 vccd1 vccd1 _13245_/A sky130_fd_sc_hd__inv_2
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14708_ _18805_/Q _13629_/X _14716_/S vssd1 vssd1 vccd1 vccd1 _14709_/A sky130_fd_sc_hd__mux2_1
X_18476_ _18547_/CLK _18476_/D vssd1 vssd1 vccd1 vccd1 _18476_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__B2 _19005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15688_ _18921_/Q _18542_/Q _15688_/S vssd1 vssd1 vccd1 vccd1 _15689_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17427_ _17483_/A vssd1 vssd1 vccd1 vccd1 _17496_/S sky130_fd_sc_hd__buf_6
XFILLER_33_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15978__A _15978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13034__B1 _11855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14639_ _18780_/Q _11879_/X _14649_/S vssd1 vssd1 vccd1 vccd1 _14640_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18354__A _18422_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17358_ _17358_/A vssd1 vssd1 vccd1 vccd1 _19591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16309_ _16309_/A vssd1 vssd1 vccd1 vccd1 _19162_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09695__B _18939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17289_ _17106_/X _19561_/Q _17293_/S vssd1 vssd1 vccd1 vccd1 _17290_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19028_ _19720_/CLK _19028_/D vssd1 vssd1 vccd1 vccd1 _19028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18028__A1 _11845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09614_ _09614_/A vssd1 vssd1 vccd1 vccd1 _09614_/X sky130_fd_sc_hd__buf_4
XFILLER_84_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09545_ _11291_/A vssd1 vssd1 vccd1 vccd1 _09546_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09476_ _15139_/A _15942_/A _15899_/B _14766_/A vssd1 vssd1 vccd1 vccd1 _09476_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_51_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16762__A1 _13857_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14792__A _14792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12379__A2 _12843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13201__A _17039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10320_ _10492_/A vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_137_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_162_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10251_ _19375_/Q _19710_/Q _10251_/S vssd1 vssd1 vccd1 vccd1 _10251_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17608__A _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11434__S0 _11154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09825__S _09903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ _10185_/A vssd1 vssd1 vccd1 vccd1 _10182_/X sky130_fd_sc_hd__buf_2
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14990_ _14990_/A _15004_/A _14990_/C vssd1 vssd1 vccd1 vccd1 _15099_/A sky130_fd_sc_hd__nor3_1
XFILLER_59_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13941_ _18554_/Q _13937_/C _13940_/Y vssd1 vssd1 vccd1 vccd1 _18554_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17778__A0 _17691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16660_ _16660_/A vssd1 vssd1 vccd1 vccd1 _19305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13872_ _12113_/A _12113_/B _13870_/X vssd1 vssd1 vccd1 vccd1 _18522_/D sky130_fd_sc_hd__a21o_1
XFILLER_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15611_ _18887_/Q _18919_/Q _15611_/S vssd1 vssd1 vccd1 vccd1 _15612_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12067__A1 _18711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ _15899_/A _12823_/B vssd1 vssd1 vccd1 vccd1 _12824_/A sky130_fd_sc_hd__and2_4
X_16591_ _19275_/Q _13819_/X _16591_/S vssd1 vssd1 vccd1 vccd1 _16592_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18330_ _18330_/A vssd1 vssd1 vccd1 vccd1 _19998_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_87_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _15542_/A _15542_/B vssd1 vssd1 vccd1 vccd1 _15542_/Y sky130_fd_sc_hd__nor2_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _14750_/B _12657_/X _12778_/A _12753_/Y vssd1 vssd1 vccd1 vccd1 _12755_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _19968_/Q _17710_/A _18263_/S vssd1 vssd1 vccd1 vccd1 _18262_/A sky130_fd_sc_hd__mux2_1
X_11705_ _11705_/A _14227_/B vssd1 vssd1 vccd1 vccd1 _11706_/A sky130_fd_sc_hd__nor2_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15473_ _15099_/X _15470_/Y _15472_/X _15268_/A vssd1 vssd1 vccd1 vccd1 _15476_/B
+ sky130_fd_sc_hd__a211o_1
X_12685_ _12756_/A _15487_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _12686_/B sky130_fd_sc_hd__a21o_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17212_ _17280_/S vssd1 vssd1 vccd1 vccd1 _17221_/S sky130_fd_sc_hd__buf_4
X_11636_ _10248_/X _11585_/X _11633_/X _11635_/Y vssd1 vssd1 vccd1 vccd1 _11636_/X
+ sky130_fd_sc_hd__a211o_1
X_14424_ _14472_/A _14431_/C vssd1 vssd1 vccd1 vccd1 _14424_/Y sky130_fd_sc_hd__nor2_1
X_18192_ _18192_/A vssd1 vssd1 vccd1 vccd1 _19937_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12934__B _12956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17143_ _17143_/A vssd1 vssd1 vccd1 vccd1 _19503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _09833_/X _11566_/X _11558_/A vssd1 vssd1 vccd1 vccd1 _11567_/X sky130_fd_sc_hd__a21o_1
X_14355_ _18683_/Q _14355_/B _14355_/C vssd1 vssd1 vccd1 vccd1 _14356_/C sky130_fd_sc_hd__and3_1
XANTENNA__10735__A _18847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10518_ _10567_/A _10517_/X _10162_/A vssd1 vssd1 vccd1 vccd1 _10518_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_144_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13306_ _18886_/Q vssd1 vssd1 vccd1 vccd1 _13306_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14516__B1 _14507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17074_ _17074_/A vssd1 vssd1 vccd1 vccd1 _17074_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14286_ _18661_/Q _14290_/D _14285_/Y vssd1 vssd1 vccd1 vccd1 _18661_/D sky130_fd_sc_hd__o21a_1
X_11498_ _11502_/A _11498_/B vssd1 vssd1 vccd1 vccd1 _11498_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16025_ _13238_/X _19042_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16026_/A sky130_fd_sc_hd__mux2_1
X_13237_ _17046_/A vssd1 vssd1 vccd1 vccd1 _17688_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10449_ _19371_/Q _19706_/Q _10449_/S vssd1 vssd1 vccd1 vccd1 _10449_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13168_ _14062_/A _13120_/A _12887_/A _18627_/Q vssd1 vssd1 vccd1 vccd1 _13168_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17952__S _17952_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12119_ _12118_/Y _18902_/Q _12179_/S vssd1 vssd1 vccd1 vccd1 _14912_/A sky130_fd_sc_hd__mux2_1
X_17976_ _19856_/Q _17023_/X _17976_/S vssd1 vssd1 vccd1 vccd1 _17977_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13099_ _13098_/X _18432_/Q _13116_/S vssd1 vssd1 vccd1 vccd1 _13100_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19715_ _19873_/CLK _19715_/D vssd1 vssd1 vccd1 vccd1 _19715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16927_ _16307_/X _19423_/Q _16931_/S vssd1 vssd1 vccd1 vccd1 _16928_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15980__B _15980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13781__A _17017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19646_ _20003_/CLK _19646_/D vssd1 vssd1 vccd1 vccd1 _19646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16858_ _16858_/A vssd1 vssd1 vccd1 vccd1 _19392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15809_ _09436_/B _11860_/A _15798_/X input61/X vssd1 vssd1 vccd1 vccd1 _15810_/B
+ sky130_fd_sc_hd__a22o_1
X_19577_ _19865_/CLK _19577_/D vssd1 vssd1 vccd1 vccd1 _19577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16789_ _16332_/X _19362_/Q _16797_/S vssd1 vssd1 vccd1 vccd1 _16790_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09330_ _18985_/Q _18940_/Q vssd1 vssd1 vccd1 vccd1 _09698_/C sky130_fd_sc_hd__or2b_1
XFILLER_80_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18528_ _18867_/CLK _18528_/D vssd1 vssd1 vccd1 vccd1 _18528_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11266__C1 _09873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10164__S0 _10141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09261_ _09261_/A _09261_/B vssd1 vssd1 vccd1 vccd1 _09264_/B sky130_fd_sc_hd__or2_1
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18459_ _19885_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11018__C1 _11157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09192_ _09272_/A vssd1 vssd1 vccd1 vccd1 _11667_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12844__B _12844_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10467__S1 _10223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10219__S1 _10223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17428__A _17496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11416__S0 _10980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12860__A _12866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16332__A _17668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10544__A1 _10822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__B1 _14672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10380__A _10380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16478__S _16486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13494__B1 _12890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_109_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _12084_/S _09498_/Y _09510_/X _09527_/X vssd1 vssd1 vccd1 vccd1 _09528_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_71_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10539__B _12849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _18971_/Q hold2/A _09459_/C vssd1 vssd1 vccd1 vccd1 _12004_/B sky130_fd_sc_hd__or3_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12470_ _12470_/A vssd1 vssd1 vccd1 vccd1 _12470_/Y sky130_fd_sc_hd__clkinv_8
X_11421_ _11421_/A _11421_/B vssd1 vssd1 vccd1 vccd1 _11421_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14140_ _14142_/B _14142_/C _14139_/Y vssd1 vssd1 vccd1 vccd1 _18619_/D sky130_fd_sc_hd__o21a_1
XANTENNA__11575__A3 _09702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11352_ _19657_/Q _19423_/Q _18488_/Q _19753_/Q _11230_/X _11021_/A vssd1 vssd1 vccd1
+ vccd1 _11352_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ _10411_/A _10303_/B vssd1 vssd1 vccd1 vccd1 _10303_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14071_ _14070_/B _14070_/C _18599_/Q vssd1 vssd1 vccd1 vccd1 _14072_/C sky130_fd_sc_hd__a21oi_1
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11283_ _11283_/A _11283_/B vssd1 vssd1 vccd1 vccd1 _11283_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_7_0_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_7_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13022_ _17010_/A vssd1 vssd1 vccd1 vccd1 _17652_/A sky130_fd_sc_hd__clkbuf_2
X_10234_ _19218_/Q _19809_/Q _19971_/Q _19186_/Q _10005_/A _10207_/A vssd1 vssd1 vccd1
+ vccd1 _10235_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input51_A io_ibus_inst[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13721__A1 _18481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17830_ _19791_/Q _17020_/X _17832_/S vssd1 vssd1 vccd1 vccd1 _17831_/A sky130_fd_sc_hd__mux2_1
X_10165_ _10392_/A _10165_/B vssd1 vssd1 vccd1 vccd1 _10165_/X sky130_fd_sc_hd__or2_1
XFILLER_79_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17761_ _17761_/A vssd1 vssd1 vccd1 vccd1 _19760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16388__S _16394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ _09833_/X _10095_/X _10292_/A vssd1 vssd1 vccd1 vccd1 _10096_/X sky130_fd_sc_hd__a21o_1
X_14973_ _14973_/A _14973_/B vssd1 vssd1 vccd1 vccd1 _15482_/B sky130_fd_sc_hd__or2_4
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19500_ _19664_/CLK _19500_/D vssd1 vssd1 vccd1 vccd1 _19500_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output138_A _12831_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10299__B1 _09884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16712_ _19328_/Q _13784_/X _16714_/S vssd1 vssd1 vccd1 vccd1 _16713_/A sky130_fd_sc_hd__mux2_1
X_13924_ _18550_/Q _13924_/B _14108_/B vssd1 vssd1 vccd1 vccd1 _13925_/C sky130_fd_sc_hd__and3_1
X_17692_ _17691_/X _19736_/Q _17698_/S vssd1 vssd1 vccd1 vccd1 _17693_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19431_ _19731_/CLK _19431_/D vssd1 vssd1 vccd1 vccd1 _19431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16643_ _16689_/S vssd1 vssd1 vccd1 vccd1 _16652_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13855_ _18516_/Q _13854_/X _13858_/S vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13788__A1 _13787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19362_ _19957_/CLK _19362_/D vssd1 vssd1 vccd1 vccd1 _19362_/Q sky130_fd_sc_hd__dfxtp_1
X_12806_ _15553_/B _12807_/B vssd1 vssd1 vccd1 vccd1 _15552_/A sky130_fd_sc_hd__and2_1
XFILLER_76_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18176__A0 _17691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16574_ _19267_/Q _13794_/X _16580_/S vssd1 vssd1 vccd1 vccd1 _16575_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12010__A _12722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13786_ _13786_/A vssd1 vssd1 vccd1 vccd1 _18494_/D sky130_fd_sc_hd__clkbuf_1
X_10998_ _11137_/A _10997_/X _09683_/A vssd1 vssd1 vccd1 vccd1 _10998_/Y sky130_fd_sc_hd__o21ai_1
X_18313_ _17681_/X _19991_/Q _18313_/S vssd1 vssd1 vccd1 vccd1 _18314_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _12743_/Y _15458_/X _15524_/X _15454_/X vssd1 vssd1 vccd1 vccd1 _15525_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19293_ _19758_/CLK _19293_/D vssd1 vssd1 vccd1 vccd1 _19293_/Q sky130_fd_sc_hd__dfxtp_1
X_12737_ _15976_/C _18925_/Q _12782_/S vssd1 vssd1 vccd1 vccd1 _12738_/A sky130_fd_sc_hd__mux2_4
XANTENNA__12460__A1 _12514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09861__C1 _09690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17012__S _17024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18244_ _19960_/Q _17684_/A _18252_/S vssd1 vssd1 vccd1 vccd1 _18245_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15456_ _18855_/Q _15363_/X _15455_/X vssd1 vssd1 vccd1 vccd1 _18855_/D sky130_fd_sc_hd__o21a_1
X_12668_ _12668_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _12670_/A sky130_fd_sc_hd__nor2_2
X_14407_ _14407_/A vssd1 vssd1 vccd1 vccd1 _14452_/A sky130_fd_sc_hd__buf_2
X_18175_ _18175_/A vssd1 vssd1 vccd1 vccd1 _19929_/D sky130_fd_sc_hd__clkbuf_1
X_11619_ _11615_/Y _11616_/X _11618_/Y vssd1 vssd1 vccd1 vccd1 _11622_/C sky130_fd_sc_hd__a21oi_1
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12212__A1 _18905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16851__S _16859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15387_ _15399_/A _15387_/B _15387_/C vssd1 vssd1 vccd1 vccd1 _15387_/X sky130_fd_sc_hd__and3_1
X_12599_ _12599_/A vssd1 vssd1 vccd1 vccd1 _12599_/Y sky130_fd_sc_hd__clkinv_4
X_17126_ _17125_/X _19498_/Q _17129_/S vssd1 vssd1 vccd1 vccd1 _17127_/A sky130_fd_sc_hd__mux2_1
X_14338_ _18677_/Q _18676_/Q _18675_/Q _14338_/D vssd1 vssd1 vccd1 vccd1 _14373_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17057_ _17057_/A vssd1 vssd1 vccd1 vccd1 _19472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14269_ _14280_/A _14275_/D vssd1 vssd1 vccd1 vccd1 _14270_/B sky130_fd_sc_hd__and2_1
XANTENNA__16152__A _16208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16008_ _16008_/A vssd1 vssd1 vccd1 vccd1 _19034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17682__S _17682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11296__A _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_191_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19947_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17959_ _19848_/Q _16998_/X _17965_/S vssd1 vssd1 vccd1 vccd1 _17960_/A sky130_fd_sc_hd__mux2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10385__S0 _10209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_110_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11314__A1_N _18836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__B _12839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19629_ _19757_/CLK _19629_/D vssd1 vssd1 vccd1 vccd1 _19629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13779__A1 _13778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11462__C _11462_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09313_ _09313_/A _11919_/C vssd1 vssd1 vccd1 vccd1 _09516_/B sky130_fd_sc_hd__or2_2
XFILLER_81_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10688__S1 _10638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12855__A _12857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18018__S _18020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09244_ _18975_/Q _18974_/Q vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__or2b_1
XFILLER_167_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17857__S _17865_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ _14756_/A _09282_/D vssd1 vssd1 vccd1 vccd1 _12866_/B sky130_fd_sc_hd__nor2_8
XANTENNA__12203__A1 _12188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10375__A _10380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_144_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19912_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_35_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11714__B1 _11713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10314__S _10314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_159_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19885_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15456__A1 _18855_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13467__B1 _09410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11970_ _12871_/A vssd1 vssd1 vccd1 vccd1 _11971_/B sky130_fd_sc_hd__inv_2
XFILLER_56_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16001__S _16009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09404__A _14227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ _19361_/Q _19696_/Q _10921_/S vssd1 vssd1 vccd1 vccd1 _10921_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16936__S _16942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10852_ _11172_/A vssd1 vssd1 vccd1 vccd1 _11015_/A sky130_fd_sc_hd__buf_2
X_13640_ _18470_/Q _13639_/X _13670_/S vssd1 vssd1 vccd1 vccd1 _13641_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10774_/Y _10778_/Y _10780_/Y _10782_/Y _09550_/A vssd1 vssd1 vccd1 vccd1
+ _10784_/A sky130_fd_sc_hd__o221a_1
X_13571_ _13589_/A _19002_/Q vssd1 vssd1 vccd1 vccd1 _13571_/Y sky130_fd_sc_hd__nand2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16708__A1 _13778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _15243_/X _15299_/X _15309_/X _15258_/X vssd1 vssd1 vccd1 vccd1 _15310_/X
+ sky130_fd_sc_hd__o211a_1
X_12522_ _12522_/A vssd1 vssd1 vccd1 vccd1 _12522_/X sky130_fd_sc_hd__clkbuf_2
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16290_/A vssd1 vssd1 vccd1 vccd1 _19156_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17381__A1 _17030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17767__S _17771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15241_ _12221_/Y _15146_/X _15240_/X _15951_/A vssd1 vssd1 vccd1 vccd1 _15241_/X
+ sky130_fd_sc_hd__a211o_1
X_12453_ _12347_/X _12451_/X _12452_/Y _12350_/X vssd1 vssd1 vccd1 vccd1 _12453_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_166_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11404_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11404_/X sky130_fd_sc_hd__or2_1
X_15172_ _15478_/A _15172_/B vssd1 vssd1 vccd1 vccd1 _15172_/X sky130_fd_sc_hd__or2_1
X_12384_ _12385_/A _14879_/A vssd1 vssd1 vccd1 vccd1 _12386_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17068__A _17068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11335_ _11335_/A _11335_/B vssd1 vssd1 vccd1 vccd1 _11335_/X sky130_fd_sc_hd__or2_1
X_14123_ _14124_/B _14529_/B _18614_/Q vssd1 vssd1 vccd1 vccd1 _14125_/B sky130_fd_sc_hd__a21oi_1
XFILLER_153_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19980_ _19980_/CLK _19980_/D vssd1 vssd1 vccd1 vccd1 _19980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18931_ _18967_/CLK _18931_/D vssd1 vssd1 vccd1 vccd1 _18931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14054_ _14745_/A vssd1 vssd1 vccd1 vccd1 _14245_/A sky130_fd_sc_hd__buf_2
X_11266_ _11058_/X _11257_/Y _11261_/Y _11265_/Y _09873_/A vssd1 vssd1 vccd1 vccd1
+ _11266_/X sky130_fd_sc_hd__o311a_1
XANTENNA__11828__B _11828_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10217_ _10522_/A vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13170__A2 _13081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13005_ _13297_/A vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__buf_4
X_18862_ _19010_/CLK _18862_/D vssd1 vssd1 vccd1 vccd1 _18862_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12005__A _18520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ _19659_/Q _19425_/Q _18490_/Q _19755_/Q _11125_/S _11077_/X vssd1 vssd1 vccd1
+ vccd1 _11197_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17813_ _19783_/Q _16992_/X _17821_/S vssd1 vssd1 vccd1 vccd1 _17814_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10148_ _10630_/A vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__buf_2
X_18793_ _19062_/CLK _18793_/D vssd1 vssd1 vccd1 vccd1 _18793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17744_ _17744_/A vssd1 vssd1 vccd1 vccd1 _19752_/D sky130_fd_sc_hd__clkbuf_1
X_10079_ _18857_/Q vssd1 vssd1 vccd1 vccd1 _10079_/Y sky130_fd_sc_hd__inv_2
X_14956_ _12738_/A _15100_/B _14956_/S vssd1 vssd1 vccd1 vccd1 _14956_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12659__B _12857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ _12745_/A _12820_/A _12748_/Y _12751_/Y _13904_/X vssd1 vssd1 vccd1 vccd1
+ _18546_/D sky130_fd_sc_hd__o221a_1
X_17675_ _17675_/A vssd1 vssd1 vccd1 vccd1 _17675_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14887_ _15306_/B _15410_/B _14908_/S vssd1 vssd1 vccd1 vccd1 _14887_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19414_ _19873_/CLK _19414_/D vssd1 vssd1 vccd1 vccd1 _19414_/Q sky130_fd_sc_hd__dfxtp_1
X_16626_ _16307_/X _19290_/Q _16630_/S vssd1 vssd1 vccd1 vccd1 _16627_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13838_ _17074_/A vssd1 vssd1 vccd1 vccd1 _13838_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19345_ _19587_/CLK _19345_/D vssd1 vssd1 vccd1 vccd1 _19345_/Q sky130_fd_sc_hd__dfxtp_1
X_16557_ _16557_/A vssd1 vssd1 vccd1 vccd1 _19259_/D sky130_fd_sc_hd__clkbuf_1
X_13769_ _18489_/Q _13768_/X _13772_/S vssd1 vssd1 vccd1 vccd1 _13770_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15508_ _14991_/X _15505_/Y _15507_/X _14998_/X vssd1 vssd1 vccd1 vccd1 _15511_/B
+ sky130_fd_sc_hd__a211o_1
X_19276_ _19997_/CLK _19276_/D vssd1 vssd1 vccd1 vccd1 _19276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16488_ _16545_/S vssd1 vssd1 vccd1 vccd1 _16497_/S sky130_fd_sc_hd__clkbuf_4
X_18227_ _18227_/A vssd1 vssd1 vccd1 vccd1 _19952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19963_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15986__A _16150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15439_ _15151_/X _15263_/X _15438_/X _15413_/X vssd1 vssd1 vccd1 vccd1 _15439_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18158_ _17665_/X _19922_/Q _18158_/S vssd1 vssd1 vccd1 vccd1 _18159_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11944__B1 _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17109_ _17646_/A vssd1 vssd1 vccd1 vccd1 _17109_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18089_ _18088_/X _19898_/Q _18095_/S vssd1 vssd1 vccd1 vccd1 _18090_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_76_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19842_/CLK sky130_fd_sc_hd__clkbuf_16
X_09931_ _09933_/A _09930_/X _09568_/A vssd1 vssd1 vccd1 vccd1 _09931_/X sky130_fd_sc_hd__o21a_1
XFILLER_171_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13697__B1 _13695_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09862_ _09862_/A _09862_/B _09862_/C vssd1 vssd1 vccd1 vccd1 _09862_/X sky130_fd_sc_hd__or3_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09793_ _09793_/A vssd1 vssd1 vccd1 vccd1 _09794_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10132__C1 _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16756__S _16758_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19693_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11268__A1_N _18838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10817__B _12841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17587__S _17595_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _20017_/CLK sky130_fd_sc_hd__clkbuf_16
X_09227_ _18962_/Q vssd1 vssd1 vccd1 vccd1 _09481_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__16491__S _16497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11935__B1 _09458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10833__S1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15677__A1 _18537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11120_ _09881_/A _11101_/X _11118_/X _09911_/A _11119_/Y vssd1 vssd1 vccd1 vccd1
+ _12831_/B sky130_fd_sc_hd__o32a_2
XFILLER_122_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11051_ _11122_/A _11048_/X _11050_/X _11137_/A vssd1 vssd1 vccd1 vccd1 _11051_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18211__S _18219_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10002_ _10342_/A vssd1 vssd1 vccd1 vccd1 _10007_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13355__S _13366_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14810_ _15004_/A vssd1 vssd1 vccd1 vccd1 _14973_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15790_ _15785_/Y _15788_/X _15789_/X _09481_/D vssd1 vssd1 vccd1 vccd1 _15791_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_91_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input14_A io_dbus_rdata[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ _14741_/A vssd1 vssd1 vccd1 vccd1 _18820_/D sky130_fd_sc_hd__clkbuf_1
X_11953_ _12859_/A _09525_/A _14807_/B _12290_/B vssd1 vssd1 vccd1 vccd1 _12432_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16666__S _16674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17460_ _17460_/A vssd1 vssd1 vccd1 vccd1 _19637_/D sky130_fd_sc_hd__clkbuf_1
X_10904_ _19665_/Q _19431_/Q _18496_/Q _19761_/Q _10892_/X _10893_/X vssd1 vssd1 vccd1
+ vccd1 _10905_/B sky130_fd_sc_hd__mux4_1
X_14672_ _14672_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14729_/A sky130_fd_sc_hd__and2_1
XFILLER_60_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11884_ _14102_/A vssd1 vssd1 vccd1 vccd1 _11884_/X sky130_fd_sc_hd__buf_4
XFILLER_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16411_ _19195_/Q _13768_/X _16413_/S vssd1 vssd1 vccd1 vccd1 _16412_/A sky130_fd_sc_hd__mux2_1
X_13623_ _13621_/X _13622_/Y _13623_/S vssd1 vssd1 vccd1 vccd1 _13623_/X sky130_fd_sc_hd__mux2_1
X_10835_ _19203_/Q _19794_/Q _19956_/Q _19171_/Q _11467_/S _10820_/A vssd1 vssd1 vccd1
+ vccd1 _10836_/B sky130_fd_sc_hd__mux4_1
X_17391_ _17391_/A vssd1 vssd1 vccd1 vccd1 _19606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19130_ _19979_/CLK _19130_/D vssd1 vssd1 vccd1 vccd1 _19130_/Q sky130_fd_sc_hd__dfxtp_1
X_16342_ _17678_/A vssd1 vssd1 vccd1 vccd1 _16342_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13554_ _13554_/A _18871_/Q _13554_/C vssd1 vssd1 vccd1 vccd1 _13565_/B sky130_fd_sc_hd__or3_1
X_10766_ _09664_/A _10765_/X _10727_/A vssd1 vssd1 vccd1 vccd1 _10766_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19061_ _19062_/CLK _19061_/D vssd1 vssd1 vccd1 vccd1 _19061_/Q sky130_fd_sc_hd__dfxtp_1
X_12505_ _18472_/Q _12343_/X _12344_/X vssd1 vssd1 vccd1 vccd1 _12505_/Y sky130_fd_sc_hd__o21ai_1
X_16273_ _16273_/A vssd1 vssd1 vccd1 vccd1 _19148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10697_ _10680_/A _10696_/X _10579_/X vssd1 vssd1 vccd1 vccd1 _10697_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12179__A0 _15925_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13485_ _18896_/Q _13486_/B vssd1 vssd1 vccd1 vccd1 _13485_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18182__A _18193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18012_ _19872_/Q _17074_/X _18020_/S vssd1 vssd1 vccd1 vccd1 _18013_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15224_ _12186_/Y _15146_/X _15223_/X _15951_/A vssd1 vssd1 vccd1 vccd1 _15224_/X
+ sky130_fd_sc_hd__a211o_1
X_12436_ _10652_/A _18913_/Q _12517_/S vssd1 vssd1 vccd1 vccd1 _12467_/A sky130_fd_sc_hd__mux2_2
XANTENNA__10729__A1 _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15155_ _15368_/A vssd1 vssd1 vccd1 vccd1 _15155_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12367_ _12368_/A _12416_/D vssd1 vssd1 vccd1 vccd1 _12369_/A sky130_fd_sc_hd__or2_1
XFILLER_154_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output82_A _11971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14106_ _14105_/B _14105_/C _18611_/Q vssd1 vssd1 vccd1 vccd1 _14107_/C sky130_fd_sc_hd__a21oi_1
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _19226_/Q _19721_/Q _11367_/S vssd1 vssd1 vccd1 vccd1 _11318_/X sky130_fd_sc_hd__mux2_1
X_19963_ _19963_/CLK _19963_/D vssd1 vssd1 vccd1 vccd1 _19963_/Q sky130_fd_sc_hd__dfxtp_1
X_12298_ _12298_/A vssd1 vssd1 vccd1 vccd1 _15270_/B sky130_fd_sc_hd__buf_2
X_15086_ _15165_/S _15078_/B _15084_/X _15085_/Y vssd1 vssd1 vccd1 vccd1 _15086_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13679__B1 _13674_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14037_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14042_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11249_ _20014_/Q _19852_/Q _19261_/Q _19031_/Q _11212_/X _11208_/X vssd1 vssd1 vccd1
+ vccd1 _11250_/B sky130_fd_sc_hd__mux4_1
X_18914_ _19350_/CLK _18914_/D vssd1 vssd1 vccd1 vccd1 _18914_/Q sky130_fd_sc_hd__dfxtp_1
X_19894_ _19896_/CLK _19894_/D vssd1 vssd1 vccd1 vccd1 _19894_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15972__C _15972_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18845_ _19792_/CLK _18845_/D vssd1 vssd1 vccd1 vccd1 _18845_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11574__A _11574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18776_ _19900_/CLK _18776_/D vssd1 vssd1 vccd1 vccd1 _18776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15988_ _16044_/A vssd1 vssd1 vccd1 vccd1 _16057_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_48_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12389__B _12389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17727_ _17726_/X _19747_/Q _17730_/S vssd1 vssd1 vccd1 vccd1 _17728_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14939_ _14935_/X _14938_/X _15020_/A vssd1 vssd1 vccd1 vccd1 _14939_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16576__S _16580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15480__S _15480_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17658_ _17658_/A vssd1 vssd1 vccd1 vccd1 _19725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16609_ _19283_/Q _13845_/X _16613_/S vssd1 vssd1 vccd1 vccd1 _16610_/A sky130_fd_sc_hd__mux2_1
X_17589_ _17135_/X _19698_/Q _17595_/S vssd1 vssd1 vccd1 vccd1 _17590_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10417__B1 _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19328_ _19824_/CLK _19328_/D vssd1 vssd1 vccd1 vccd1 _19328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19259_ _19485_/CLK _19259_/D vssd1 vssd1 vccd1 vccd1 _19259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09918__S _09918_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11749__A _14665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14125__A _14143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09914_ _18862_/Q vssd1 vssd1 vccd1 vccd1 _09914_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14331__A1 _18674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20034_ _20034_/CLK _20034_/D vssd1 vssd1 vccd1 vccd1 _20034_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input6_A io_dbus_rdata[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _15980_/B _12864_/C vssd1 vssd1 vccd1 vccd1 _11529_/A sky130_fd_sc_hd__or2_2
XFILLER_100_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17870__S _17876_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09776_ _09776_/A vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12299__B _15270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16486__S _16486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ _10892_/A vssd1 vssd1 vccd1 vccd1 _10907_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10503__S0 _10125_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10551_ _10668_/A _10551_/B _10551_/C vssd1 vssd1 vccd1 vccd1 _10551_/X sky130_fd_sc_hd__or3_1
XANTENNA__18206__S _18206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17110__S _17113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10482_ _10001_/A _10481_/X _10162_/A vssd1 vssd1 vccd1 vccd1 _10482_/Y sky130_fd_sc_hd__o21ai_1
X_13270_ _19900_/Q _13290_/B vssd1 vssd1 vccd1 vccd1 _13270_/X sky130_fd_sc_hd__and2_1
XANTENNA__14570__A1 _11801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12221_ _12221_/A vssd1 vssd1 vccd1 vccd1 _12221_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_136_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10563__A _10572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ _12191_/A _12477_/C vssd1 vssd1 vccd1 vccd1 _12153_/D sky130_fd_sc_hd__xor2_1
XFILLER_135_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11103_ _19662_/Q _19428_/Q _18493_/Q _19758_/Q _11293_/A _09737_/A vssd1 vssd1 vccd1
+ vccd1 _11103_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13125__A2 _12889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16960_ _16355_/X _19438_/Q _16964_/S vssd1 vssd1 vccd1 vccd1 _16961_/A sky130_fd_sc_hd__mux2_1
X_12083_ _09466_/A _12082_/X _15899_/B vssd1 vssd1 vccd1 vccd1 _12083_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11034_ _11149_/A _11033_/X _09791_/A vssd1 vssd1 vccd1 vccd1 _11034_/Y sky130_fd_sc_hd__o21ai_1
X_15911_ _18997_/Q _15910_/X _15914_/S vssd1 vssd1 vccd1 vccd1 _15912_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16891_ _16891_/A vssd1 vssd1 vccd1 vccd1 _19407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11231__S1 _11108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13085__S _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17780__S _17782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18630_ _19683_/CLK _18630_/D vssd1 vssd1 vccd1 vccd1 _18630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15842_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15842_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18561_ _18741_/CLK _18561_/D vssd1 vssd1 vccd1 vccd1 _18561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _15773_/A _15773_/B vssd1 vssd1 vccd1 vccd1 _15773_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12985_ _19058_/Q _12878_/A _13269_/A _18794_/Q vssd1 vssd1 vccd1 vccd1 _12985_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _19662_/Q vssd1 vssd1 vccd1 vccd1 _17513_/A sky130_fd_sc_hd__clkbuf_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_157_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14724_ _14724_/A vssd1 vssd1 vccd1 vccd1 _18812_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _15899_/A _12033_/S _11935_/X vssd1 vssd1 vccd1 vccd1 _11936_/X sky130_fd_sc_hd__o21a_1
X_18492_ _19757_/CLK _18492_/D vssd1 vssd1 vccd1 vccd1 _18492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__S0 _09725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17443_ _17443_/A vssd1 vssd1 vccd1 vccd1 _19629_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ _14655_/A vssd1 vssd1 vccd1 vccd1 _18784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _15765_/A vssd1 vssd1 vccd1 vccd1 _11867_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13114__A _17023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13606_ _11860_/D _13605_/Y _13623_/S vssd1 vssd1 vccd1 vccd1 _13606_/X sky130_fd_sc_hd__mux2_1
X_10818_ _10818_/A _10818_/B vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__and2_1
X_17374_ _19599_/Q _17020_/X _17376_/S vssd1 vssd1 vccd1 vccd1 _17375_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13061__A1 _13560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14586_ _14595_/A _14586_/B vssd1 vssd1 vccd1 vccd1 _14587_/A sky130_fd_sc_hd__and2_1
X_11798_ _11831_/A _11798_/B vssd1 vssd1 vccd1 vccd1 _11798_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19113_ _19641_/CLK _19113_/D vssd1 vssd1 vccd1 vccd1 _19113_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11072__B1 _11003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16325_ _16325_/A vssd1 vssd1 vccd1 vccd1 _19167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13537_ _13595_/A vssd1 vssd1 vccd1 vccd1 _13583_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_158_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10749_ _19366_/Q _19701_/Q _10749_/S vssd1 vssd1 vccd1 vccd1 _10749_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19044_ _19865_/CLK _19044_/D vssd1 vssd1 vccd1 vccd1 _19044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16256_ _13180_/X _19141_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _16257_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13468_ _18484_/Q _13511_/A _11847_/X _18708_/Q _13467_/Y vssd1 vssd1 vccd1 vccd1
+ _13468_/X sky130_fd_sc_hd__a221o_1
X_15207_ _14978_/X _15206_/X _15097_/X vssd1 vssd1 vccd1 vccd1 _15478_/B sky130_fd_sc_hd__o21a_1
XANTENNA__14561__A1 _18995_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ _12791_/A _12413_/Y _12154_/X vssd1 vssd1 vccd1 vccd1 _12419_/Y sky130_fd_sc_hd__a21oi_1
X_16187_ _13219_/X _19111_/Q _16195_/S vssd1 vssd1 vccd1 vccd1 _16188_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10473__A _10473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13399_ _14327_/B _12889_/X _12887_/X _18640_/Q vssd1 vssd1 vccd1 vccd1 _13399_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15138_ _15247_/A _15138_/B vssd1 vssd1 vccd1 vccd1 _15142_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13784__A _17020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17256__A _17267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19946_ _19946_/CLK _19946_/D vssd1 vssd1 vccd1 vccd1 _19946_/Q sky130_fd_sc_hd__dfxtp_1
X_15069_ _15061_/X _15067_/X _15171_/S vssd1 vssd1 vccd1 vccd1 _15069_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19877_ _19877_/CLK _19877_/D vssd1 vssd1 vccd1 vccd1 _19877_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16066__A1 _14562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09630_ _09973_/A vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18828_ _18960_/CLK _18828_/D vssd1 vssd1 vccd1 vccd1 _18828_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_96_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09561_ _10712_/A vssd1 vssd1 vccd1 vccd1 _09562_/A sky130_fd_sc_hd__clkbuf_2
X_18759_ _18762_/CLK _18759_/D vssd1 vssd1 vccd1 vccd1 _18759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18087__A _18104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09492_ _09492_/A _12845_/A vssd1 vssd1 vccd1 vccd1 _15899_/A sky130_fd_sc_hd__nand2_4
XFILLER_64_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12847__B _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13024__A _13502_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_4_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13959__A _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12863__A _12863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17865__S _17865_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13107__A2 _13070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11213__S1 _11208_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20017_ _20017_/CLK _20017_/D vssd1 vssd1 vccd1 vccd1 _20017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09828_ _09828_/A vssd1 vssd1 vccd1 vccd1 _11237_/A sky130_fd_sc_hd__buf_4
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09759_ _09759_/A vssd1 vssd1 vccd1 vccd1 _10680_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13633__S _13689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13291__A1 _18474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12766_/A _12769_/X _12770_/S vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__mux2_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11721_ _11897_/A _19010_/Q vssd1 vssd1 vccd1 vccd1 _11721_/Y sky130_fd_sc_hd__nand2_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14440_ _14452_/A _14440_/B _14440_/C vssd1 vssd1 vccd1 vccd1 _18707_/D sky130_fd_sc_hd__nor3_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11652_ _11659_/B vssd1 vssd1 vccd1 vccd1 _11975_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10603_ _10836_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _10603_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14371_ _18687_/Q _14371_/B _14371_/C vssd1 vssd1 vccd1 vccd1 _14378_/C sky130_fd_sc_hd__and3_1
XANTENNA__12251__C1 _12154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11583_ _11644_/A _10247_/Y _11524_/Y _11643_/A vssd1 vssd1 vccd1 vccd1 _11583_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16110_ _16110_/A vssd1 vssd1 vccd1 vccd1 _19077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13322_ _17062_/A vssd1 vssd1 vccd1 vccd1 _17704_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10534_ _10149_/A _10533_/X _09796_/A vssd1 vssd1 vccd1 vccd1 _10534_/X sky130_fd_sc_hd__o21a_1
X_17090_ _17090_/A vssd1 vssd1 vccd1 vccd1 _17090_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13588__B _13588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16041_ _16041_/A vssd1 vssd1 vccd1 vccd1 _19049_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14543__A1 _18753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ _10458_/X _10460_/X _10462_/X _10464_/X _09875_/A vssd1 vssd1 vccd1 vccd1
+ _10465_/X sky130_fd_sc_hd__a221o_1
XFILLER_129_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13253_ input10/X _13231_/X _13234_/X vssd1 vssd1 vccd1 vccd1 _13261_/A sky130_fd_sc_hd__a21oi_1
XFILLER_171_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12204_ _12204_/A _12204_/B vssd1 vssd1 vccd1 vccd1 _12205_/A sky130_fd_sc_hd__and2_4
XFILLER_108_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10396_ _09702_/X _10384_/X _10395_/X _09843_/A _18854_/Q vssd1 vssd1 vccd1 vccd1
+ _12853_/B sky130_fd_sc_hd__a32oi_4
XFILLER_108_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13184_ _18879_/Q vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__buf_2
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13808__S _13820_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19800_ _19864_/CLK _19800_/D vssd1 vssd1 vccd1 vccd1 _19800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12135_ _12108_/A _12107_/A _12134_/X vssd1 vssd1 vccd1 vccd1 _12135_/X sky130_fd_sc_hd__a21o_1
X_17992_ _19863_/Q _17046_/X _17998_/S vssd1 vssd1 vccd1 vccd1 _17993_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11109__A1 _09721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19731_ _19731_/CLK _19731_/D vssd1 vssd1 vccd1 vccd1 _19731_/Q sky130_fd_sc_hd__dfxtp_1
X_16943_ _16943_/A vssd1 vssd1 vccd1 vccd1 _19430_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18037__A2 _13648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ _12066_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12066_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11204__S1 _11065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10868__B1 _09843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _11017_/A _19232_/Q vssd1 vssd1 vccd1 vccd1 _11017_/Y sky130_fd_sc_hd__nor2_1
X_16874_ _16874_/A vssd1 vssd1 vccd1 vccd1 _19399_/D sky130_fd_sc_hd__clkbuf_1
X_19662_ _19758_/CLK _19662_/D vssd1 vssd1 vccd1 vccd1 _19662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15825_ _15831_/A _15825_/B vssd1 vssd1 vccd1 vccd1 _15826_/A sky130_fd_sc_hd__and2_1
X_18613_ _18745_/CLK _18613_/D vssd1 vssd1 vccd1 vccd1 _18613_/Q sky130_fd_sc_hd__dfxtp_1
X_19593_ _19947_/CLK _19593_/D vssd1 vssd1 vccd1 vccd1 _19593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17015__S _17024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _15769_/A vssd1 vssd1 vccd1 vccd1 _15756_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18544_ _18544_/CLK _18544_/D vssd1 vssd1 vccd1 vccd1 _18544_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12968_ _13226_/A vssd1 vssd1 vccd1 vccd1 _13360_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10096__A1 _09833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12667__B _15487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ _14729_/A vssd1 vssd1 vccd1 vccd1 _14716_/S sky130_fd_sc_hd__buf_2
X_11919_ _11919_/A _11919_/B _11919_/C vssd1 vssd1 vccd1 vccd1 _11920_/D sky130_fd_sc_hd__or3_1
X_18475_ _19900_/CLK _18475_/D vssd1 vssd1 vccd1 vccd1 _18475_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10468__A _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ _15687_/A vssd1 vssd1 vccd1 vccd1 _18920_/D sky130_fd_sc_hd__clkbuf_1
X_12899_ _19486_/Q vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__inv_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _17426_/A _17426_/B vssd1 vssd1 vccd1 vccd1 _17483_/A sky130_fd_sc_hd__or2_4
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ _14638_/A vssd1 vssd1 vccd1 vccd1 _18779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15978__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17357_ _19591_/Q _16992_/X _17365_/S vssd1 vssd1 vccd1 vccd1 _17358_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14569_ _14569_/A vssd1 vssd1 vccd1 vccd1 _18759_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12683__A _12753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16308_ _16307_/X _19162_/Q _16314_/S vssd1 vssd1 vccd1 vccd1 _16309_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17288_ _17288_/A vssd1 vssd1 vccd1 vccd1 _19560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19027_ _20010_/CLK _19027_/D vssd1 vssd1 vccd1 vccd1 _19027_/Q sky130_fd_sc_hd__dfxtp_1
X_16239_ _13023_/X _19133_/Q _16247_/S vssd1 vssd1 vccd1 vccd1 _16240_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13337__A2 _11776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11899__A2 _11898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17484__A0 _17179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19929_ _19993_/CLK _19929_/D vssd1 vssd1 vccd1 vccd1 _19929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11238__S _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13019__A _13359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09613_ _09646_/A vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__buf_2
XFILLER_56_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12858__A _12863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _09544_/A vssd1 vssd1 vccd1 vccd1 _11291_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09477__B1 _09476_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09475_ _15633_/B _09475_/B vssd1 vssd1 vccd1 vccd1 _14766_/A sky130_fd_sc_hd__nand2_4
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17595__S _17595_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_105_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_clock_A clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10250_ _10248_/X _11635_/A vssd1 vssd1 vccd1 vccd1 _11524_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11434__S1 _11107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10181_ _10355_/A _10181_/B vssd1 vssd1 vccd1 vccd1 _10181_/X sky130_fd_sc_hd__and2_1
XFILLER_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _13967_/A _13945_/C vssd1 vssd1 vccd1 vccd1 _13940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13871_ _12076_/A _12076_/B _13870_/X vssd1 vssd1 vccd1 vccd1 _18521_/D sky130_fd_sc_hd__a21o_1
XFILLER_75_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15610_ _15610_/A vssd1 vssd1 vccd1 vccd1 _18886_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11672__A _11772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12822_ _12827_/A _12822_/B vssd1 vssd1 vccd1 vccd1 _12822_/Y sky130_fd_sc_hd__nor2_8
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16590_ _16590_/A vssd1 vssd1 vccd1 vccd1 _19274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_3_0_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _15366_/A _15538_/Y _15540_/X _15268_/A vssd1 vssd1 vccd1 vccd1 _15544_/B
+ sky130_fd_sc_hd__a211o_1
X_12753_ _12753_/A _12863_/B vssd1 vssd1 vccd1 vccd1 _12753_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16674__S _16674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14983__A _15103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18260_ _18260_/A vssd1 vssd1 vccd1 vccd1 _19967_/D sky130_fd_sc_hd__clkbuf_1
X_11704_ _11870_/A vssd1 vssd1 vccd1 vccd1 _12943_/A sky130_fd_sc_hd__buf_2
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _15155_/X _15474_/B _15102_/X _15471_/X vssd1 vssd1 vccd1 vccd1 _15472_/X
+ sky130_fd_sc_hd__o211a_1
X_12684_ _09261_/A _12657_/X _12778_/A _12683_/Y vssd1 vssd1 vccd1 vccd1 _15498_/A
+ sky130_fd_sc_hd__a211o_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17267_/A vssd1 vssd1 vccd1 vccd1 _17280_/S sky130_fd_sc_hd__buf_4
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14433_/D vssd1 vssd1 vccd1 vccd1 _14431_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18191_ _17713_/X _19937_/Q _18191_/S vssd1 vssd1 vccd1 vccd1 _18192_/A sky130_fd_sc_hd__mux2_1
X_11635_ _11635_/A _11635_/B vssd1 vssd1 vccd1 vccd1 _11635_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__13567__A2 _14548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15961__B1 _15955_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17142_ _17141_/X _19503_/Q _17145_/S vssd1 vssd1 vccd1 vccd1 _17143_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14354_ _14355_/B _14355_/C _18683_/Q vssd1 vssd1 vccd1 vccd1 _14356_/B sky130_fd_sc_hd__a21oi_1
X_11566_ _19255_/Q _19750_/Q _11566_/S vssd1 vssd1 vccd1 vccd1 _11566_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13305_ _13305_/A vssd1 vssd1 vccd1 vccd1 _18444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10517_ _18442_/Q _19471_/Q _19508_/Q _19082_/Q _10529_/S _10011_/A vssd1 vssd1 vccd1
+ vccd1 _10517_/X sky130_fd_sc_hd__mux4_1
X_17073_ _17073_/A vssd1 vssd1 vccd1 vccd1 _19477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14285_ _14288_/A _14285_/B vssd1 vssd1 vccd1 vccd1 _14285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11497_ _18437_/Q _19466_/Q _19503_/Q _19077_/Q _11486_/S _10856_/X vssd1 vssd1 vccd1
+ vccd1 _11498_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12008__A _12393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16024_ _16024_/A vssd1 vssd1 vccd1 vccd1 _19041_/D sky130_fd_sc_hd__clkbuf_1
X_13236_ _13223_/X _13230_/X _13235_/Y vssd1 vssd1 vccd1 vccd1 _17046_/A sky130_fd_sc_hd__a21oi_4
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10448_ _10448_/A _10448_/B vssd1 vssd1 vccd1 vccd1 _10448_/X sky130_fd_sc_hd__and2_1
XFILLER_156_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _18595_/Q vssd1 vssd1 vccd1 vccd1 _14062_/A sky130_fd_sc_hd__clkbuf_2
X_10379_ _20030_/Q _19868_/Q _19277_/Q _19047_/Q _10209_/S _09745_/A vssd1 vssd1 vccd1
+ vccd1 _10380_/B sky130_fd_sc_hd__mux4_1
XFILLER_112_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12118_ _12118_/A vssd1 vssd1 vccd1 vccd1 _12118_/Y sky130_fd_sc_hd__inv_2
X_17975_ _17975_/A vssd1 vssd1 vccd1 vccd1 _19855_/D sky130_fd_sc_hd__clkbuf_1
X_13098_ _17662_/A vssd1 vssd1 vccd1 vccd1 _13098_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19714_ _19972_/CLK _19714_/D vssd1 vssd1 vccd1 vccd1 _19714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16926_ _16926_/A vssd1 vssd1 vccd1 vccd1 _19422_/D sky130_fd_sc_hd__clkbuf_1
X_12049_ _18053_/A vssd1 vssd1 vccd1 vccd1 _13508_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19645_ _19999_/CLK _19645_/D vssd1 vssd1 vccd1 vccd1 _19645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16857_ _16310_/X _19392_/Q _16859_/S vssd1 vssd1 vccd1 vccd1 _16858_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15808_ _15808_/A vssd1 vssd1 vccd1 vccd1 _18965_/D sky130_fd_sc_hd__clkbuf_1
X_19576_ _20026_/CLK _19576_/D vssd1 vssd1 vccd1 vccd1 _19576_/Q sky130_fd_sc_hd__dfxtp_1
X_16788_ _16834_/S vssd1 vssd1 vccd1 vccd1 _16797_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15989__A _16057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15739_ _18941_/Q _15738_/B _15738_/Y _15730_/X vssd1 vssd1 vccd1 vccd1 _18941_/D
+ sky130_fd_sc_hd__o211a_1
X_18527_ _18997_/CLK _18527_/D vssd1 vssd1 vccd1 vccd1 _18527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14893__A _15016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18365__A _18422_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10164__S1 _10163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ _18986_/Q vssd1 vssd1 vccd1 vccd1 _09261_/B sky130_fd_sc_hd__buf_4
X_18458_ _18526_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17409_ _19615_/Q _17071_/X _17409_/S vssd1 vssd1 vccd1 vccd1 _17410_/A sky130_fd_sc_hd__mux2_1
X_09191_ _11919_/A vssd1 vssd1 vccd1 vccd1 _09272_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18389_ _18389_/A vssd1 vssd1 vccd1 vccd1 _20024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11416__S1 _10972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12860__B _12866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17457__A0 _17141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11741__A1 _18471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13246__A1 _12875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_31_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09527_ _14804_/D _14765_/B _09527_/C _09527_/D vssd1 vssd1 vccd1 vccd1 _09527_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__15899__A _15899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11352__S0 _11230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09897__A _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09458_/A hold4/A _18970_/Q vssd1 vssd1 vccd1 vccd1 _09459_/C sky130_fd_sc_hd__or3_1
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09870__B1 _09690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10836__A _10836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ _11697_/A _11697_/B _09399_/A _15775_/A vssd1 vssd1 vccd1 vccd1 _11869_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_40_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11420_ _19913_/Q _19527_/Q _19977_/Q _19096_/Q _09586_/A _11208_/A vssd1 vssd1 vccd1
+ vccd1 _11421_/B sky130_fd_sc_hd__mux4_2
XFILLER_165_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17619__A _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ _10854_/A _11348_/X _11350_/X vssd1 vssd1 vccd1 vccd1 _11351_/X sky130_fd_sc_hd__a21o_1
XFILLER_126_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14742__S _14742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ _20031_/Q _19869_/Q _19278_/Q _19048_/Q _09595_/A _10260_/A vssd1 vssd1 vccd1
+ vccd1 _10303_/B sky130_fd_sc_hd__mux4_1
XFILLER_137_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14070_ _18599_/Q _14070_/B _14070_/C vssd1 vssd1 vccd1 vccd1 _14072_/B sky130_fd_sc_hd__and3_1
XFILLER_141_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11282_ _19916_/Q _19530_/Q _19980_/Q _19099_/Q _11063_/X _11065_/X vssd1 vssd1 vccd1
+ vccd1 _11283_/B sky130_fd_sc_hd__mux4_2
XFILLER_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13021_ _13005_/X _13020_/X _12906_/A input28/X vssd1 vssd1 vccd1 vccd1 _17010_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_10233_ _10438_/A _10232_/X _09779_/A vssd1 vssd1 vccd1 vccd1 _10233_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__15139__A _15139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10164_ _19682_/Q _19448_/Q _18513_/Q _19778_/Q _10141_/X _10163_/X vssd1 vssd1 vccd1
+ vccd1 _10165_/B sky130_fd_sc_hd__mux4_1
XFILLER_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input44_A io_ibus_inst[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10095_ _19248_/Q _19743_/Q _10095_/S vssd1 vssd1 vccd1 vccd1 _10095_/X sky130_fd_sc_hd__mux2_1
X_17760_ _17665_/X _19760_/Q _17760_/S vssd1 vssd1 vccd1 vccd1 _17761_/A sky130_fd_sc_hd__mux2_1
X_14972_ _15458_/A _14972_/B _14972_/C vssd1 vssd1 vccd1 vccd1 _14972_/X sky130_fd_sc_hd__or3_1
XFILLER_75_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13923_ _13924_/B _14108_/B _18550_/Q vssd1 vssd1 vccd1 vccd1 _13925_/B sky130_fd_sc_hd__a21oi_1
XFILLER_48_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16711_ _16711_/A vssd1 vssd1 vccd1 vccd1 _19327_/D sky130_fd_sc_hd__clkbuf_1
X_17691_ _17691_/A vssd1 vssd1 vccd1 vccd1 _17691_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11496__B1 _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10299__B2 _10298_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12498__A _12498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17620__A0 _17179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19430_ _19664_/CLK _19430_/D vssd1 vssd1 vccd1 vccd1 _19430_/Q sky130_fd_sc_hd__dfxtp_1
X_16642_ _16642_/A vssd1 vssd1 vccd1 vccd1 _19297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13854_ _17090_/A vssd1 vssd1 vccd1 vccd1 _13854_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12805_ _12804_/Y _18928_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12807_/B sky130_fd_sc_hd__mux2_4
X_16573_ _16573_/A vssd1 vssd1 vccd1 vccd1 _19266_/D sky130_fd_sc_hd__clkbuf_1
X_19361_ _19664_/CLK _19361_/D vssd1 vssd1 vccd1 vccd1 _19361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ _18494_/Q _13784_/X _13788_/S vssd1 vssd1 vccd1 vccd1 _13786_/A sky130_fd_sc_hd__mux2_1
X_10997_ _19328_/Q _19599_/Q _19823_/Q _19567_/Q _10995_/X _10996_/X vssd1 vssd1 vccd1
+ vccd1 _10997_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11343__S0 _10618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16187__A0 _13219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18312_ _18312_/A vssd1 vssd1 vccd1 vccd1 _19990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15524_ _15243_/A _15098_/X _15523_/X _15093_/X vssd1 vssd1 vccd1 vccd1 _15524_/X
+ sky130_fd_sc_hd__o211a_2
XANTENNA__15602__A _15602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ _19981_/CLK _19292_/D vssd1 vssd1 vccd1 vccd1 _19292_/Q sky130_fd_sc_hd__dfxtp_1
X_12736_ _15520_/A _12736_/B vssd1 vssd1 vccd1 vccd1 _12740_/A sky130_fd_sc_hd__xnor2_1
XFILLER_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10471__A1 _10424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18243_ _18265_/A vssd1 vssd1 vccd1 vccd1 _18252_/S sky130_fd_sc_hd__buf_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09600__A _10972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15455_ _12599_/Y _15364_/X _15453_/X _15454_/X vssd1 vssd1 vccd1 vccd1 _15455_/X
+ sky130_fd_sc_hd__a211o_1
X_12667_ _12667_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _12668_/B sky130_fd_sc_hd__nor2_1
XFILLER_169_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14406_ _14411_/C _14409_/C _14405_/Y vssd1 vssd1 vccd1 vccd1 _18697_/D sky130_fd_sc_hd__o21a_1
X_18174_ _17688_/X _19929_/Q _18180_/S vssd1 vssd1 vccd1 vccd1 _18175_/A sky130_fd_sc_hd__mux2_1
X_11618_ _10818_/A _11621_/A _11510_/X vssd1 vssd1 vccd1 vccd1 _11618_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15386_ _15384_/X _15380_/Y _15385_/Y vssd1 vssd1 vccd1 vccd1 _15387_/C sky130_fd_sc_hd__a21oi_1
X_12598_ _12598_/A _12598_/B vssd1 vssd1 vccd1 vccd1 _12599_/A sky130_fd_sc_hd__xnor2_4
XFILLER_144_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17125_ _17662_/A vssd1 vssd1 vccd1 vccd1 _17125_/X sky130_fd_sc_hd__clkbuf_2
X_14337_ _14356_/A _14337_/B _14369_/B vssd1 vssd1 vccd1 vccd1 _18676_/D sky130_fd_sc_hd__nor3_1
X_11549_ _11543_/A _11548_/X _09568_/A vssd1 vssd1 vccd1 vccd1 _11549_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17056_ _19472_/Q _17055_/X _17056_/S vssd1 vssd1 vccd1 vccd1 _17057_/A sky130_fd_sc_hd__mux2_1
X_14268_ _14479_/A vssd1 vssd1 vccd1 vccd1 _14288_/A sky130_fd_sc_hd__clkbuf_2
X_16007_ _13098_/X _19034_/Q _16009_/S vssd1 vssd1 vccd1 vccd1 _16008_/A sky130_fd_sc_hd__mux2_1
X_13219_ _17684_/A vssd1 vssd1 vccd1 vccd1 _13219_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11577__A _15982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17963__S _17965_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _14245_/A vssd1 vssd1 vccd1 vccd1 _14239_/A sky130_fd_sc_hd__buf_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _17958_/A vssd1 vssd1 vccd1 vccd1 _19847_/D sky130_fd_sc_hd__clkbuf_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16909_ _16909_/A vssd1 vssd1 vccd1 vccd1 _19415_/D sky130_fd_sc_hd__clkbuf_1
X_17889_ _19817_/Q _17001_/X _17893_/S vssd1 vssd1 vccd1 vccd1 _17890_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19628_ _19757_/CLK _19628_/D vssd1 vssd1 vccd1 vccd1 _19628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11239__B1 _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14976__A1 _09347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19559_ _20010_/CLK _19559_/D vssd1 vssd1 vccd1 vccd1 _19559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11334__S0 _10980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09312_ _14813_/B _14811_/B _14811_/C vssd1 vssd1 vccd1 vccd1 _14765_/A sky130_fd_sc_hd__or3_2
XFILLER_34_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12855__B _12855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ _09247_/C vssd1 vssd1 vccd1 vccd1 _11919_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15231__B _15234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09174_ _18975_/Q _18973_/Q vssd1 vssd1 vccd1 vccd1 _09282_/D sky130_fd_sc_hd__or2_4
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13967__A _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17439__A _17496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16489__S _16497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15406__B _15410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10920_ _11122_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _10920_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09404__B _11869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14416__B1 _14366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ _10953_/S vssd1 vssd1 vccd1 vccd1 _11488_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_147_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17113__S _17113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _19002_/Q _13570_/B vssd1 vssd1 vccd1 vccd1 _13570_/X sky130_fd_sc_hd__or2_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _11473_/A _10781_/X _09685_/A vssd1 vssd1 vccd1 vccd1 _10782_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12546_/A _12521_/B vssd1 vssd1 vccd1 vccd1 _12521_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__14719__A1 _13667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15240_ _14830_/X _15228_/X _15239_/X _15089_/X vssd1 vssd1 vccd1 vccd1 _15240_/X
+ sky130_fd_sc_hd__o211a_1
X_12452_ _12452_/A _12483_/C vssd1 vssd1 vccd1 vccd1 _12452_/Y sky130_fd_sc_hd__nand2_1
X_11403_ _19193_/Q _19784_/Q _19946_/Q _19161_/Q _19384_/Q _19385_/Q vssd1 vssd1 vccd1
+ vccd1 _11404_/B sky130_fd_sc_hd__mux4_1
X_15171_ _15167_/X _15170_/X _15171_/S vssd1 vssd1 vccd1 vccd1 _15172_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12781__A _15980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ _10760_/A _18911_/Q _12409_/A vssd1 vssd1 vccd1 vccd1 _14879_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10756__A2 _10753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14122_ _14126_/D vssd1 vssd1 vccd1 vccd1 _14529_/B sky130_fd_sc_hd__clkbuf_2
X_11334_ _19194_/Q _19785_/Q _19947_/Q _19162_/Q _10980_/A _11322_/A vssd1 vssd1 vccd1
+ vccd1 _11335_/B sky130_fd_sc_hd__mux4_1
XFILLER_4_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18930_ _18967_/CLK _18930_/D vssd1 vssd1 vccd1 vccd1 _18930_/Q sky130_fd_sc_hd__dfxtp_1
X_14053_ _14088_/A _14053_/B _14053_/C vssd1 vssd1 vccd1 vccd1 _18593_/D sky130_fd_sc_hd__nor3_1
X_11265_ _11252_/A _11262_/X _11264_/X vssd1 vssd1 vccd1 vccd1 _11265_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ _13004_/A vssd1 vssd1 vccd1 vccd1 _18428_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18094__A0 _18852_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ _10216_/A vssd1 vssd1 vccd1 vccd1 _10388_/S sky130_fd_sc_hd__buf_4
X_18861_ _19025_/CLK _18861_/D vssd1 vssd1 vccd1 vccd1 _18861_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_output150_A _12485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11196_ _09880_/A _11183_/X _11194_/X _09911_/A _11195_/Y vssd1 vssd1 vccd1 vccd1
+ _12827_/B sky130_fd_sc_hd__o32a_2
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15447__A2 _15449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17812_ _17880_/S vssd1 vssd1 vccd1 vccd1 _17821_/S sky130_fd_sc_hd__clkbuf_4
X_10147_ _10843_/A vssd1 vssd1 vccd1 vccd1 _10630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18792_ _19062_/CLK _18792_/D vssd1 vssd1 vccd1 vccd1 _18792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17743_ _17640_/X _19752_/Q _17749_/S vssd1 vssd1 vccd1 vccd1 _17744_/A sky130_fd_sc_hd__mux2_1
X_14955_ _12760_/A _15078_/B _14955_/S vssd1 vssd1 vccd1 vccd1 _14955_/X sky130_fd_sc_hd__mux2_1
X_10078_ _10078_/A vssd1 vssd1 vccd1 vccd1 _10078_/X sky130_fd_sc_hd__buf_4
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_0_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17812__A _17880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13906_ _18545_/Q _13900_/X _12723_/X _12727_/X _13904_/X vssd1 vssd1 vccd1 vccd1
+ _18545_/D sky130_fd_sc_hd__o221a_1
XFILLER_63_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17674_ _17674_/A vssd1 vssd1 vccd1 vccd1 _19730_/D sky130_fd_sc_hd__clkbuf_1
X_14886_ _14886_/A vssd1 vssd1 vccd1 vccd1 _15410_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19413_ _20035_/CLK _19413_/D vssd1 vssd1 vccd1 vccd1 _19413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10692__A1 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ _13837_/A vssd1 vssd1 vccd1 vccd1 _18510_/D sky130_fd_sc_hd__clkbuf_1
X_16625_ _16625_/A vssd1 vssd1 vccd1 vccd1 _19289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12956__A _12956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11316__S0 _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__A _11860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19344_ _19839_/CLK _19344_/D vssd1 vssd1 vccd1 vccd1 _19344_/Q sky130_fd_sc_hd__dfxtp_1
X_16556_ _19259_/Q _13768_/X _16558_/S vssd1 vssd1 vccd1 vccd1 _16557_/A sky130_fd_sc_hd__mux2_1
X_13768_ _17004_/A vssd1 vssd1 vccd1 vccd1 _13768_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15907__A0 _11982_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ _18545_/Q _12719_/B vssd1 vssd1 vccd1 vccd1 _12768_/C sky130_fd_sc_hd__and2_1
X_15507_ _15101_/X _15509_/B _14994_/X _15506_/X vssd1 vssd1 vccd1 vccd1 _15507_/X
+ sky130_fd_sc_hd__o211a_1
X_19275_ _20028_/CLK _19275_/D vssd1 vssd1 vccd1 vccd1 _19275_/Q sky130_fd_sc_hd__dfxtp_1
X_16487_ _16487_/A vssd1 vssd1 vccd1 vccd1 _19228_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13699_ _13699_/A _13699_/B vssd1 vssd1 vccd1 vccd1 _13699_/Y sky130_fd_sc_hd__nand2_1
X_18226_ _19952_/Q _17659_/A _18230_/S vssd1 vssd1 vccd1 vccd1 _18227_/A sky130_fd_sc_hd__mux2_1
X_15438_ _15438_/A _15438_/B _15438_/C vssd1 vssd1 vccd1 vccd1 _15438_/X sky130_fd_sc_hd__and3_1
XANTENNA__15986__B _16691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13787__A _17023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18157_ _18157_/A vssd1 vssd1 vccd1 vccd1 _19921_/D sky130_fd_sc_hd__clkbuf_1
X_15369_ _15369_/A vssd1 vssd1 vccd1 vccd1 _15369_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11944__A1 _09702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17108_ _17108_/A vssd1 vssd1 vccd1 vccd1 _19492_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11944__B2 _09347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18088_ _18850_/Q _11748_/X _18101_/S vssd1 vssd1 vccd1 vccd1 _18088_/X sky130_fd_sc_hd__mux2_2
XFILLER_172_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17039_ _17039_/A vssd1 vssd1 vccd1 vccd1 _17039_/X sky130_fd_sc_hd__buf_2
X_09930_ _18452_/Q _19481_/Q _19518_/Q _19092_/Q _09668_/S _09614_/A vssd1 vssd1 vccd1
+ vccd1 _09930_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10055__S0 _10254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09996__S0 _10356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09861_ _11543_/A _09858_/X _09860_/X _09690_/X vssd1 vssd1 vccd1 vccd1 _09862_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _09792_/A vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__clkbuf_2
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11555__S0 _11553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12866__A _12866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14557__S _14601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11770__A _12060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17868__S _17876_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09226_ _18963_/Q vssd1 vssd1 vccd1 vccd1 _09481_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15126__B2 _12046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11050_ _11050_/A _11050_/B vssd1 vssd1 vccd1 vccd1 _11050_/X sky130_fd_sc_hd__and2_1
XFILLER_89_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10001_ _10001_/A vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__buf_2
XFILLER_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11945__A _11945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16012__S _16020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10371__B1 _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16947__S _16953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11546__S0 _11532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11156__S _11156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14740_ _18820_/Q _13742_/X _14742_/S vssd1 vssd1 vccd1 vccd1 _14741_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11952_ _09522_/A _15740_/A _09275_/A _14812_/C vssd1 vssd1 vccd1 vccd1 _14807_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _10895_/X _10898_/X _10900_/X _10902_/X _09804_/A vssd1 vssd1 vccd1 vccd1
+ _10903_/X sky130_fd_sc_hd__a221o_1
XFILLER_72_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14671_ _14671_/A vssd1 vssd1 vccd1 vccd1 _18789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11883_ _14159_/A vssd1 vssd1 vccd1 vccd1 _14102_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_33_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16410_ _16410_/A vssd1 vssd1 vccd1 vccd1 _19194_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13622_ _13630_/A _13630_/C vssd1 vssd1 vccd1 vccd1 _13622_/Y sky130_fd_sc_hd__xnor2_4
X_10834_ _09624_/A _10833_/X _10712_/X vssd1 vssd1 vccd1 vccd1 _10834_/Y sky130_fd_sc_hd__o21ai_1
X_17390_ _19606_/Q _17042_/X _17398_/S vssd1 vssd1 vccd1 vccd1 _17391_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13612__B2 _19007_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17778__S _17782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16341_ _16341_/A vssd1 vssd1 vccd1 vccd1 _19172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13553_ _13528_/X _13551_/X _13552_/Y _13532_/X _19000_/Q vssd1 vssd1 vccd1 vccd1
+ _13553_/X sky130_fd_sc_hd__a32o_4
XFILLER_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10765_ _19236_/Q _19731_/Q _10872_/S vssd1 vssd1 vccd1 vccd1 _10765_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19060_ _19882_/CLK _19060_/D vssd1 vssd1 vccd1 vccd1 _19060_/Q sky130_fd_sc_hd__dfxtp_1
X_12504_ _12498_/A _12502_/X _12697_/S vssd1 vssd1 vccd1 vccd1 _12504_/X sky130_fd_sc_hd__mux2_1
X_16272_ _13302_/X _19148_/Q _16280_/S vssd1 vssd1 vccd1 vccd1 _16273_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_190_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19485_/CLK sky130_fd_sc_hd__clkbuf_16
X_13484_ input25/X _13340_/X _13368_/X vssd1 vssd1 vccd1 vccd1 _13484_/Y sky130_fd_sc_hd__a21oi_1
X_10696_ _19335_/Q _19606_/Q _19830_/Q _19574_/Q _10637_/S _10010_/A vssd1 vssd1 vccd1
+ vccd1 _10696_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18011_ _18011_/A vssd1 vssd1 vccd1 vccd1 _18020_/S sky130_fd_sc_hd__buf_4
XANTENNA__13376__B1 _11852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15223_ _14830_/X _15204_/X _15222_/X _15089_/X vssd1 vssd1 vccd1 vccd1 _15223_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12435_ _15373_/A _12435_/B vssd1 vssd1 vccd1 vccd1 _12437_/A sky130_fd_sc_hd__xor2_4
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_0_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15154_ _15160_/A _15160_/B vssd1 vssd1 vccd1 vccd1 _15154_/Y sky130_fd_sc_hd__nand2_1
X_12366_ _12368_/A _12366_/B vssd1 vssd1 vccd1 vccd1 _12377_/A sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_153_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14105_ _18611_/Q _14105_/B _14105_/C vssd1 vssd1 vccd1 vccd1 _14107_/B sky130_fd_sc_hd__and3_1
XANTENNA__13128__B1 _13124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11317_ _11414_/A _11317_/B vssd1 vssd1 vccd1 vccd1 _11317_/X sky130_fd_sc_hd__or2_1
X_19962_ _20026_/CLK _19962_/D vssd1 vssd1 vccd1 vccd1 _19962_/Q sky130_fd_sc_hd__dfxtp_1
X_15085_ _15142_/A _15078_/Y _15365_/A vssd1 vssd1 vccd1 vccd1 _15085_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12297_ _12297_/A _14859_/A vssd1 vssd1 vccd1 vccd1 _12301_/A sky130_fd_sc_hd__xor2_4
XFILLER_4_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18067__A0 _18844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output75_A _12364_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14036_ _14044_/A _14036_/B _14036_/C vssd1 vssd1 vccd1 vccd1 _18587_/D sky130_fd_sc_hd__nor3_1
X_18913_ _18918_/CLK _18913_/D vssd1 vssd1 vccd1 vccd1 _18913_/Q sky130_fd_sc_hd__dfxtp_1
X_11248_ _11287_/A _11248_/B vssd1 vssd1 vccd1 vccd1 _11248_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19893_ _19896_/CLK _19893_/D vssd1 vssd1 vccd1 vccd1 _19893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16617__A1 _13857_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17018__S _17024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18844_ _19792_/CLK _18844_/D vssd1 vssd1 vccd1 vccd1 _18844_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10362__B1 _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14231__A _14385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ _11225_/A _11179_/B vssd1 vssd1 vccd1 vccd1 _11179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18775_ _19900_/CLK _18775_/D vssd1 vssd1 vccd1 vccd1 _18775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15987_ _17426_/A _18352_/C vssd1 vssd1 vccd1 vccd1 _16044_/A sky130_fd_sc_hd__or2_4
XANTENNA__16857__S _16859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__S0 _09635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17726_ _17726_/A vssd1 vssd1 vccd1 vccd1 _17726_/X sky130_fd_sc_hd__clkbuf_2
X_14938_ _14936_/X _14937_/X _14938_/S vssd1 vssd1 vccd1 vccd1 _14938_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_143_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18744_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17657_ _17656_/X _19725_/Q _17666_/S vssd1 vssd1 vccd1 vccd1 _17658_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14869_ _14869_/A vssd1 vssd1 vccd1 vccd1 _14908_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_91_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16608_ _16608_/A vssd1 vssd1 vccd1 vccd1 _19282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_78_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17588_ _17588_/A vssd1 vssd1 vccd1 vccd1 _19697_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10417__A1 _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19327_ _19951_/CLK _19327_/D vssd1 vssd1 vccd1 vccd1 _19327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16539_ _19252_/Q _13848_/X _16541_/S vssd1 vssd1 vccd1 vccd1 _16540_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_158_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19899_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09995__A _09995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19258_ _19485_/CLK _19258_/D vssd1 vssd1 vccd1 vccd1 _19258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18209_ _18265_/A vssd1 vssd1 vccd1 vccd1 _18278_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_129_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19189_ _20006_/CLK _19189_/D vssd1 vssd1 vccd1 vccd1 _19189_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12625__S _12814_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12590__A1 _09454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17717__A _17717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16621__A _16689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ _09913_/A vssd1 vssd1 vccd1 vccd1 _09913_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_160_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20033_ _20033_/CLK _20033_/D vssd1 vssd1 vccd1 vccd1 _20033_/Q sky130_fd_sc_hd__dfxtp_1
X_09844_ _09702_/X _09808_/X _09839_/X _09843_/X _18863_/Q vssd1 vssd1 vccd1 vccd1
+ _12864_/C sky130_fd_sc_hd__a32o_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14619__A0 _18774_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09775_ _09775_/A vssd1 vssd1 vccd1 vccd1 _09776_/A sky130_fd_sc_hd__buf_2
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16767__S _16775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11853__B1 _11852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17598__S _17606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10550_ _09988_/A _10547_/X _10549_/X _09687_/A vssd1 vssd1 vccd1 vccd1 _10551_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ _19488_/Q vssd1 vssd1 vccd1 vccd1 _13226_/A sky130_fd_sc_hd__buf_2
XFILLER_167_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10481_ _18443_/Q _19472_/Q _19509_/Q _19083_/Q _10388_/S _10223_/A vssd1 vssd1 vccd1
+ vccd1 _10481_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16007__S _16009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14316__A _18670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13220__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ _12220_/A _12220_/B vssd1 vssd1 vccd1 vccd1 _12221_/A sky130_fd_sc_hd__xnor2_4
XFILLER_170_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09982__C1 _09876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ _18524_/Q vssd1 vssd1 vccd1 vccd1 _12191_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18222__S _18230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11102_ _11441_/S vssd1 vssd1 vccd1 vccd1 _11293_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_151_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ _18980_/Q vssd1 vssd1 vccd1 vccd1 _12082_/X sky130_fd_sc_hd__buf_4
XANTENNA__15986__C_N _15735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13366__S _13366_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11033_ _20017_/Q _19855_/Q _19264_/Q _19034_/Q _10892_/A _11022_/X vssd1 vssd1 vccd1
+ vccd1 _11033_/X sky130_fd_sc_hd__mux4_1
X_15910_ _12032_/X _11292_/X _15946_/A vssd1 vssd1 vccd1 vccd1 _15910_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15147__A _15147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16890_ _16358_/X _19407_/Q _16892_/S vssd1 vssd1 vccd1 vccd1 _16891_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11541__C1 _09876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15841_ _15883_/A vssd1 vssd1 vccd1 vccd1 _15861_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16677__S _16685_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _20027_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13890__A _14385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12097__B1 _12094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18560_ _18741_/CLK _18560_/D vssd1 vssd1 vccd1 vccd1 _18560_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _12984_/A vssd1 vssd1 vccd1 vccd1 _12984_/X sky130_fd_sc_hd__buf_2
X_15772_ _09261_/B _15765_/X _15771_/X _15769_/X vssd1 vssd1 vccd1 vccd1 _18954_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17511_ _17511_/A vssd1 vssd1 vccd1 vccd1 _19661_/D sky130_fd_sc_hd__clkbuf_1
X_11935_ _12290_/B _12317_/A _12315_/A _09458_/A vssd1 vssd1 vccd1 vccd1 _11935_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14723_ _18812_/Q _13685_/X _14727_/S vssd1 vssd1 vccd1 vccd1 _14724_/A sky130_fd_sc_hd__mux2_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output113_A _12842_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18491_ _20016_/CLK _18491_/D vssd1 vssd1 vccd1 vccd1 _18491_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _14663_/A _14654_/B vssd1 vssd1 vccd1 vccd1 _14655_/A sky130_fd_sc_hd__and2_1
XFILLER_72_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17442_ _17119_/X _19629_/Q _17448_/S vssd1 vssd1 vccd1 vccd1 _17443_/A sky130_fd_sc_hd__mux2_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _15719_/A vssd1 vssd1 vccd1 vccd1 _15765_/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_75_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19974_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13597__A0 _18464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13605_ _13614_/B _13605_/B vssd1 vssd1 vccd1 vccd1 _13605_/Y sky130_fd_sc_hd__nand2_1
X_10817_ _15938_/C _12841_/A vssd1 vssd1 vccd1 vccd1 _10818_/B sky130_fd_sc_hd__or2_1
XFILLER_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14585_ _18764_/Q _13563_/A _14598_/S vssd1 vssd1 vccd1 vccd1 _14586_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17373_ _17373_/A vssd1 vssd1 vccd1 vccd1 _19598_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18193__A _18193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11797_ _18717_/Q _11776_/X _11796_/X vssd1 vssd1 vccd1 vccd1 _11798_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19112_ _20024_/CLK _19112_/D vssd1 vssd1 vccd1 vccd1 _19112_/Q sky130_fd_sc_hd__dfxtp_1
X_13536_ _13554_/C _13536_/B vssd1 vssd1 vccd1 vccd1 _13536_/Y sky130_fd_sc_hd__nand2_1
X_16324_ _16323_/X _19167_/Q _16330_/S vssd1 vssd1 vccd1 vccd1 _16325_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10748_ _10748_/A _10748_/B vssd1 vssd1 vccd1 vccd1 _10748_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13349__A0 _18856_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19043_ _19864_/CLK _19043_/D vssd1 vssd1 vccd1 vccd1 _19043_/Q sky130_fd_sc_hd__dfxtp_1
X_16255_ _16255_/A vssd1 vssd1 vccd1 vccd1 _19140_/D sky130_fd_sc_hd__clkbuf_1
X_13467_ _13466_/Y _13373_/B _09410_/A vssd1 vssd1 vccd1 vccd1 _13467_/Y sky130_fd_sc_hd__a21oi_1
X_10679_ _19207_/Q _19798_/Q _19960_/Q _19175_/Q _10637_/S _10638_/X vssd1 vssd1 vccd1
+ vccd1 _10680_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _14922_/S _14919_/X _14984_/X vssd1 vssd1 vccd1 vccd1 _15206_/X sky130_fd_sc_hd__o21a_1
XFILLER_173_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10258__S0 _09657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__B1 _12020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12418_ _12446_/B _12791_/A _12417_/X vssd1 vssd1 vccd1 vccd1 _12418_/X sky130_fd_sc_hd__or3b_1
X_16186_ _16208_/A vssd1 vssd1 vccd1 vccd1 _16195_/S sky130_fd_sc_hd__buf_2
XANTENNA__14561__A2 _12933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13398_ _18672_/Q vssd1 vssd1 vccd1 vccd1 _14327_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15137_ _14858_/X _15136_/X _15074_/X vssd1 vssd1 vccd1 vccd1 _15137_/X sky130_fd_sc_hd__o21a_1
XFILLER_153_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12349_ _12349_/A _12374_/C vssd1 vssd1 vccd1 vccd1 _12349_/Y sky130_fd_sc_hd__nand2_1
XFILLER_153_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19726_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14313__A2 _14314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19945_ _19946_/CLK _19945_/D vssd1 vssd1 vccd1 vccd1 _19945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15068_ _15068_/A vssd1 vssd1 vccd1 vccd1 _15171_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14019_ _14102_/A vssd1 vssd1 vccd1 vccd1 _14019_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19876_ _19876_/CLK _19876_/D vssd1 vssd1 vccd1 vccd1 _19876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10430__S0 _10209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18827_ _18975_/CLK _18827_/D vssd1 vssd1 vccd1 vccd1 _18827_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_28_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19567_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16587__S _16591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14896__A _14927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ _09560_/A vssd1 vssd1 vccd1 vccd1 _10712_/A sky130_fd_sc_hd__buf_2
X_18758_ _19062_/CLK _18758_/D vssd1 vssd1 vccd1 vccd1 _18758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17709_ _17709_/A vssd1 vssd1 vccd1 vccd1 _19741_/D sky130_fd_sc_hd__clkbuf_1
X_09491_ _09491_/A vssd1 vssd1 vccd1 vccd1 _12845_/A sky130_fd_sc_hd__buf_2
X_18689_ _19882_/CLK _18689_/D vssd1 vssd1 vccd1 vccd1 _18689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13052__A2 _13164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18307__S _18313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12863__B _12863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10664__A _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14570__S _14601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10326__B1 _09547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09827_ _11019_/A vssd1 vssd1 vccd1 vccd1 _09828_/A sky130_fd_sc_hd__inv_2
X_20016_ _20016_/CLK _20016_/D vssd1 vssd1 vccd1 vccd1 _20016_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16497__S _16497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09758_ _11502_/A vssd1 vssd1 vccd1 vccd1 _09759_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_101_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _09980_/A vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13291__A2 _11755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11720_ _14552_/A vssd1 vssd1 vccd1 vccd1 _11897_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11659_/B _14756_/B vssd1 vssd1 vccd1 vccd1 _14758_/B sky130_fd_sc_hd__or2_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18217__S _18219_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10602_ _19336_/Q _19607_/Q _19831_/Q _19575_/Q _10655_/S _10654_/A vssd1 vssd1 vccd1
+ vccd1 _10603_/B sky130_fd_sc_hd__mux4_1
X_14370_ _14371_/B _14371_/C _18687_/Q vssd1 vssd1 vccd1 vccd1 _14372_/B sky130_fd_sc_hd__a21oi_1
X_11582_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11582_/X sky130_fd_sc_hd__or2_1
X_13321_ _13309_/X _13317_/Y _13320_/Y vssd1 vssd1 vccd1 vccd1 _17062_/A sky130_fd_sc_hd__a21oi_4
X_10533_ _19338_/Q _19609_/Q _19833_/Q _19577_/Q _10574_/S _10011_/A vssd1 vssd1 vccd1
+ vccd1 _10533_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10801__A1 _10843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16960__S _16964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17190__A0 _17189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16040_ _13354_/X _19049_/Q _16042_/S vssd1 vssd1 vccd1 vccd1 _16041_/A sky130_fd_sc_hd__mux2_1
X_13252_ _13252_/A vssd1 vssd1 vccd1 vccd1 _18441_/D sky130_fd_sc_hd__clkbuf_1
X_10464_ _10411_/A _10463_/X _10192_/X vssd1 vssd1 vccd1 vccd1 _10464_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12203_ _12188_/X _12195_/X _12197_/X _12202_/Y vssd1 vssd1 vccd1 vccd1 _12204_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_136_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13751__B1 _16075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _18879_/Q _13183_/B vssd1 vssd1 vccd1 vccd1 _13224_/C sky130_fd_sc_hd__and2_1
XFILLER_151_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10565__B1 _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10395_ _10162_/X _10390_/X _10392_/X _10394_/X _09822_/A vssd1 vssd1 vccd1 vccd1
+ _10395_/X sky130_fd_sc_hd__a221o_4
XFILLER_135_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_26_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12134_ _16069_/A _12134_/B vssd1 vssd1 vccd1 vccd1 _12134_/X sky130_fd_sc_hd__and2b_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17991_ _17991_/A vssd1 vssd1 vccd1 vccd1 _19862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17791__S _17793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19730_ _20023_/CLK _19730_/D vssd1 vssd1 vccd1 vccd1 _19730_/Q sky130_fd_sc_hd__dfxtp_1
X_16942_ _16329_/X _19430_/Q _16942_/S vssd1 vssd1 vccd1 vccd1 _16943_/A sky130_fd_sc_hd__mux2_1
X_12065_ _15758_/A _12065_/B vssd1 vssd1 vccd1 vccd1 _12163_/C sky130_fd_sc_hd__nand2_1
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10868__A1 _09702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ _19663_/Q _19429_/Q _18494_/Q _19759_/Q _11017_/A _11015_/X vssd1 vssd1 vccd1
+ vccd1 _11016_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10412__S0 _10319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19661_ _19757_/CLK _19661_/D vssd1 vssd1 vccd1 vccd1 _19661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10868__B2 _18844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16873_ _16332_/X _19399_/Q _16881_/S vssd1 vssd1 vccd1 vccd1 _16874_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13824__S _13836_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10963__S1 _10893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18612_ _18744_/CLK _18612_/D vssd1 vssd1 vccd1 vccd1 _18612_/Q sky130_fd_sc_hd__dfxtp_1
X_15824_ _18970_/Q _15816_/X _15820_/X input65/X vssd1 vssd1 vccd1 vccd1 _15825_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16200__S _16206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19592_ _19816_/CLK _19592_/D vssd1 vssd1 vccd1 vccd1 _19592_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12609__A2 _15449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12948__B _13373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18543_ _18928_/CLK _18543_/D vssd1 vssd1 vccd1 vccd1 _18543_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15755_ _18948_/Q _15760_/B vssd1 vssd1 vccd1 vccd1 _15755_/X sky130_fd_sc_hd__or2_1
X_12967_ _13297_/A vssd1 vssd1 vccd1 vccd1 _12967_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11918_ _11918_/A vssd1 vssd1 vccd1 vccd1 _11918_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _14706_/A vssd1 vssd1 vccd1 vccd1 _18804_/D sky130_fd_sc_hd__clkbuf_1
X_18474_ _18544_/CLK _18474_/D vssd1 vssd1 vccd1 vccd1 _18474_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ _12875_/X _12892_/X _12895_/Y _12897_/X vssd1 vssd1 vccd1 vccd1 _12898_/X
+ sky130_fd_sc_hd__a211o_1
X_15686_ _18920_/Q _18541_/Q _15688_/S vssd1 vssd1 vccd1 vccd1 _15687_/A sky130_fd_sc_hd__mux2_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _17425_/A vssd1 vssd1 vccd1 vccd1 _19622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11849_ _19893_/Q _11845_/X _11847_/X _18690_/Q _11848_/X vssd1 vssd1 vccd1 vccd1
+ _11849_/X sky130_fd_sc_hd__a221o_1
X_14637_ _14646_/A _14637_/B vssd1 vssd1 vccd1 vccd1 _14638_/A sky130_fd_sc_hd__and2_1
XFILLER_159_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15978__C _15978_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17031__S _17040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17356_ _17424_/S vssd1 vssd1 vccd1 vccd1 _17365_/S sky130_fd_sc_hd__buf_4
XFILLER_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14568_ _14577_/A _14568_/B vssd1 vssd1 vccd1 vccd1 _14569_/A sky130_fd_sc_hd__and2_1
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12683__B _12858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16307_ _17643_/A vssd1 vssd1 vccd1 vccd1 _16307_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17181__A0 _17179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13519_ _13689_/S _13519_/B vssd1 vssd1 vccd1 vccd1 _16072_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10484__A _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17287_ _17103_/X _19560_/Q _17293_/S vssd1 vssd1 vccd1 vccd1 _17288_/A sky130_fd_sc_hd__mux2_1
X_14499_ _14501_/A _14501_/C _14465_/X vssd1 vssd1 vccd1 vccd1 _14499_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19026_ _20010_/CLK _19026_/D vssd1 vssd1 vccd1 vccd1 _19026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15731__A1 _18970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16238_ _16295_/S vssd1 vssd1 vccd1 vccd1 _16247_/S sky130_fd_sc_hd__buf_2
XFILLER_86_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17267__A _17267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16169_ _13065_/X _19103_/Q _16173_/S vssd1 vssd1 vccd1 vccd1 _16170_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19928_ _19993_/CLK _19928_/D vssd1 vssd1 vccd1 vccd1 _19928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10423__S _10470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10403__S0 _10319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19859_ _20021_/CLK _19859_/D vssd1 vssd1 vccd1 vccd1 _19859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18098__A _18115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09612_ _09612_/A vssd1 vssd1 vccd1 vccd1 _09646_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__13734__S _16066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12858__B _12858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09543_ _18976_/Q _09465_/C _10077_/A vssd1 vssd1 vccd1 vccd1 _09544_/A sky130_fd_sc_hd__o21ai_1
XFILLER_37_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15234__B _15234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09477__A1 _13439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09474_ _14749_/B _12055_/A _12055_/B _12004_/C vssd1 vssd1 vccd1 vccd1 _09475_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__12481__B1 _12522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09659__S _09659_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17876__S _17876_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16780__S _16786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10642__S0 _09726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ _19250_/Q _19745_/Q _10180_/S vssd1 vssd1 vccd1 vccd1 _10181_/B sky130_fd_sc_hd__mux2_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12114__A _12114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13870_ _14529_/A vssd1 vssd1 vccd1 vccd1 _13870_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16020__S _16020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12768__B _18547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12821_ _18549_/Q _12790_/X _12816_/X _12820_/Y vssd1 vssd1 vccd1 vccd1 _12821_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ _15155_/X _15542_/B _15369_/A _15539_/X vssd1 vssd1 vccd1 vccd1 _15540_/X
+ sky130_fd_sc_hd__o211a_1
X_12752_ _12745_/A _12673_/X _12748_/Y _12751_/Y vssd1 vssd1 vccd1 vccd1 _12752_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11703_/A vssd1 vssd1 vccd1 vccd1 _11870_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _15539_/A _15474_/A vssd1 vssd1 vccd1 vccd1 _15471_/X sky130_fd_sc_hd__or2_1
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12753_/A _12858_/B vssd1 vssd1 vccd1 vccd1 _12683_/Y sky130_fd_sc_hd__nor2_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _18280_/B _17635_/B vssd1 vssd1 vccd1 vccd1 _17267_/A sky130_fd_sc_hd__or2_4
X_14422_ _18702_/Q _18701_/Q _14422_/C _14422_/D vssd1 vssd1 vccd1 vccd1 _14433_/D
+ sky130_fd_sc_hd__and4_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11634_/A _11634_/B vssd1 vssd1 vccd1 vccd1 _11635_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18190_ _18190_/A vssd1 vssd1 vccd1 vccd1 _19936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17141_ _17678_/A vssd1 vssd1 vccd1 vccd1 _17141_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14353_ _14355_/B _14355_/C _14352_/Y vssd1 vssd1 vccd1 vccd1 _18682_/D sky130_fd_sc_hd__o21a_1
X_11565_ _11565_/A _11565_/B vssd1 vssd1 vccd1 vccd1 _11565_/X sky130_fd_sc_hd__and2_1
XFILLER_11_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _13302_/X _18444_/Q _13366_/S vssd1 vssd1 vccd1 vccd1 _13305_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10516_ _10520_/A _10516_/B vssd1 vssd1 vccd1 vccd1 _10516_/Y sky130_fd_sc_hd__nor2_1
X_17072_ _19477_/Q _17071_/X _17072_/S vssd1 vssd1 vccd1 vccd1 _17073_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10881__S0 _10704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14284_ _18661_/Q _18660_/Q _14287_/D vssd1 vssd1 vccd1 vccd1 _14285_/B sky130_fd_sc_hd__and3_1
X_11496_ _09794_/A _11493_/X _11495_/X _09819_/A vssd1 vssd1 vccd1 vccd1 _11496_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16023_ _13219_/X _19041_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16024_/A sky130_fd_sc_hd__mux2_1
X_13235_ input8/X _13231_/X _13234_/X vssd1 vssd1 vccd1 vccd1 _13235_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13724__B1 _13700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10447_ _19243_/Q _19738_/Q _10447_/S vssd1 vssd1 vccd1 vccd1 _10448_/B sky130_fd_sc_hd__mux2_1
XFILLER_136_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13166_ _18803_/Q _11841_/A _12879_/A _18770_/Q _13165_/X vssd1 vssd1 vccd1 vccd1
+ _13166_/X sky130_fd_sc_hd__a221o_2
X_10378_ _10484_/A _10377_/X _10162_/A vssd1 vssd1 vccd1 vccd1 _10378_/X sky130_fd_sc_hd__o21a_1
XFILLER_112_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12117_ _15160_/A _12117_/B vssd1 vssd1 vccd1 vccd1 _12121_/A sky130_fd_sc_hd__xnor2_1
XFILLER_69_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18410__S _18418_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17974_ _19855_/Q _17020_/X _17976_/S vssd1 vssd1 vccd1 vccd1 _17975_/A sky130_fd_sc_hd__mux2_1
X_13097_ _17020_/A vssd1 vssd1 vccd1 vccd1 _17662_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19713_ _19942_/CLK _19713_/D vssd1 vssd1 vccd1 vccd1 _19713_/Q sky130_fd_sc_hd__dfxtp_1
X_16925_ _16304_/X _19422_/Q _16931_/S vssd1 vssd1 vccd1 vccd1 _16926_/A sky130_fd_sc_hd__mux2_1
X_12048_ _13511_/B vssd1 vssd1 vccd1 vccd1 _18053_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11863__A _15715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19644_ _19644_/CLK _19644_/D vssd1 vssd1 vccd1 vccd1 _19644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16856_ _16856_/A vssd1 vssd1 vccd1 vccd1 _19391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15807_ _15807_/A _15807_/B vssd1 vssd1 vccd1 vccd1 _15808_/A sky130_fd_sc_hd__or2_1
X_19575_ _19828_/CLK _19575_/D vssd1 vssd1 vccd1 vccd1 _19575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16787_ _16787_/A vssd1 vssd1 vccd1 vccd1 _19361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13999_ _18574_/Q _18573_/Q _13999_/C vssd1 vssd1 vccd1 vccd1 _14001_/B sky130_fd_sc_hd__and3_1
XFILLER_46_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18526_ _18526_/CLK _18526_/D vssd1 vssd1 vccd1 vccd1 _18526_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11266__A1 _11058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ _15738_/A _15738_/B vssd1 vssd1 vccd1 vccd1 _15738_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18457_ _19885_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15669_ _18912_/Q _12416_/C _15677_/S vssd1 vssd1 vccd1 vccd1 _15670_/A sky130_fd_sc_hd__mux2_1
X_17408_ _17408_/A vssd1 vssd1 vccd1 vccd1 _19614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09190_ _09306_/A _12003_/B vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__or2_2
XFILLER_159_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18388_ _17684_/X _20024_/Q _18396_/S vssd1 vssd1 vccd1 vccd1 _18389_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17339_ _17339_/A vssd1 vssd1 vccd1 vccd1 _17348_/S sky130_fd_sc_hd__buf_4
XFILLER_119_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16901__A0 _16374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19009_ _19010_/CLK _19009_/D vssd1 vssd1 vccd1 vccd1 _19009_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_146_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16105__S _16111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12860__C _12860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15468__B1 _15467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18320__S _18324_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13494__A2 _11815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13464__S _13464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16775__S _16775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13246__A2 _18850_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09526_ _14805_/A _14804_/B _11948_/A _09525_/X vssd1 vssd1 vccd1 vccd1 _09527_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10465__C1 _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09457_ _18976_/Q vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__buf_4
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09870__A1 _11538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09388_ _15779_/A _18957_/Q _18960_/Q _18959_/Q vssd1 vssd1 vccd1 vccd1 _09399_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_8_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12757__A1 _14993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17145__A0 _17144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__S _10328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11013__A _15930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ _09828_/A _11349_/X _11111_/A vssd1 vssd1 vccd1 vccd1 _11350_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10863__S0 _10787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10301_ _10301_/A vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13639__S _13689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11281_ _11003_/X _11276_/X _11278_/X _11280_/X _11133_/A vssd1 vssd1 vccd1 vccd1
+ _11281_/X sky130_fd_sc_hd__a221o_1
X_13020_ _12936_/A _13014_/X _13046_/C _13019_/Y vssd1 vssd1 vccd1 vccd1 _13020_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_10232_ _18450_/Q _19479_/Q _19516_/Q _19090_/Q _10330_/S _10013_/A vssd1 vssd1 vccd1
+ vccd1 _10232_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15139__B _15183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10163_ _10473_/A vssd1 vssd1 vccd1 vccd1 _10163_/X sky130_fd_sc_hd__buf_4
XFILLER_126_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18230__S _18230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input37_A io_ibus_inst[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10094_ _19376_/Q _19711_/Q _10094_/S vssd1 vssd1 vccd1 vccd1 _10094_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14971_ _12811_/A _12812_/Y _15007_/B _14970_/X vssd1 vssd1 vccd1 vccd1 _14972_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15155__A _15368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16710_ _19327_/Q _13781_/X _16714_/S vssd1 vssd1 vccd1 vccd1 _16711_/A sky130_fd_sc_hd__mux2_1
X_13922_ _13929_/D vssd1 vssd1 vccd1 vccd1 _14108_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17690_ _17690_/A vssd1 vssd1 vccd1 vccd1 _19735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16641_ _16329_/X _19297_/Q _16641_/S vssd1 vssd1 vccd1 vccd1 _16642_/A sky130_fd_sc_hd__mux2_1
X_13853_ _13853_/A vssd1 vssd1 vccd1 vccd1 _18515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16685__S _16685_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11833__D _11833_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12804_ _15982_/B vssd1 vssd1 vccd1 vccd1 _12804_/Y sky130_fd_sc_hd__inv_2
X_19360_ _19985_/CLK _19360_/D vssd1 vssd1 vccd1 vccd1 _19360_/Q sky130_fd_sc_hd__dfxtp_1
X_16572_ _19266_/Q _13790_/X _16580_/S vssd1 vssd1 vccd1 vccd1 _16573_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10996_ _10996_/A vssd1 vssd1 vccd1 vccd1 _10996_/X sky130_fd_sc_hd__buf_2
X_13784_ _17020_/A vssd1 vssd1 vccd1 vccd1 _13784_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18311_ _17678_/X _19990_/Q _18313_/S vssd1 vssd1 vccd1 vccd1 _18312_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11343__S1 _11086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11799__A2 _18997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10456__C1 _10194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ _14977_/X _15125_/B _15522_/X _15005_/X vssd1 vssd1 vccd1 vccd1 _15523_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19291_ _19981_/CLK _19291_/D vssd1 vssd1 vccd1 vccd1 _19291_/Q sky130_fd_sc_hd__dfxtp_1
X_12735_ _12756_/A _15509_/A _12708_/B vssd1 vssd1 vccd1 vccd1 _12736_/B sky130_fd_sc_hd__a21boi_1
XFILLER_16_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _18242_/A vssd1 vssd1 vccd1 vccd1 _19959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12666_ _12666_/A vssd1 vssd1 vccd1 vccd1 _12668_/A sky130_fd_sc_hd__inv_2
X_15454_ _15920_/A vssd1 vssd1 vccd1 vccd1 _15454_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12748__A1 _12338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17136__A0 _17135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11617_ _11617_/A _11617_/B _11617_/C vssd1 vssd1 vccd1 vccd1 _11621_/A sky130_fd_sc_hd__nand3_1
X_14405_ _14411_/C _14409_/C _14366_/X vssd1 vssd1 vccd1 vccd1 _14405_/Y sky130_fd_sc_hd__a21oi_1
X_18173_ _18173_/A vssd1 vssd1 vccd1 vccd1 _19928_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13122__B _13451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15385_ _15385_/A _15385_/B vssd1 vssd1 vccd1 vccd1 _15385_/Y sky130_fd_sc_hd__nor2_1
X_12597_ _12550_/A _12550_/B _12574_/A _12596_/Y vssd1 vssd1 vccd1 vccd1 _12598_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__18405__S _18407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17124_ _17124_/A vssd1 vssd1 vccd1 vccd1 _19497_/D sky130_fd_sc_hd__clkbuf_1
X_11548_ _18455_/Q _19484_/Q _19521_/Q _19095_/Q _11534_/S _09660_/A vssd1 vssd1 vccd1
+ vccd1 _11548_/X sky130_fd_sc_hd__mux4_2
X_14336_ _18676_/Q _14336_/B _18674_/Q _14336_/D vssd1 vssd1 vccd1 vccd1 _14369_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17055_ _17055_/A vssd1 vssd1 vccd1 vccd1 _17055_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14267_ _14745_/A vssd1 vssd1 vccd1 vccd1 _14479_/A sky130_fd_sc_hd__clkbuf_2
X_11479_ _09624_/A _11478_/X _10712_/X vssd1 vssd1 vccd1 vccd1 _11479_/X sky130_fd_sc_hd__o21a_1
XFILLER_143_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13218_ _17042_/A vssd1 vssd1 vccd1 vccd1 _17684_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16006_ _16006_/A vssd1 vssd1 vccd1 vccd1 _19033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11577__B _12866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14198_ _14315_/A _14198_/B _14200_/B vssd1 vssd1 vccd1 vccd1 _18638_/D sky130_fd_sc_hd__nor3_1
XFILLER_152_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13149_ _17030_/A vssd1 vssd1 vccd1 vccd1 _17672_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17957_ _19847_/Q _16992_/X _17965_/S vssd1 vssd1 vccd1 vccd1 _17958_/A sky130_fd_sc_hd__mux2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15870__B1 _15789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16908_ _16384_/X _19415_/Q _16914_/S vssd1 vssd1 vccd1 vccd1 _16909_/A sky130_fd_sc_hd__mux2_1
X_17888_ _17888_/A vssd1 vssd1 vccd1 vccd1 _19816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19627_ _19981_/CLK _19627_/D vssd1 vssd1 vccd1 vccd1 _19627_/Q sky130_fd_sc_hd__dfxtp_1
X_16839_ _17201_/A _16839_/B vssd1 vssd1 vccd1 vccd1 _16840_/A sky130_fd_sc_hd__and2_1
XFILLER_53_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18376__A _18422_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11239__A1 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19558_ _19846_/CLK _19558_/D vssd1 vssd1 vccd1 vccd1 _19558_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_148_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10002__A _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14976__A2 _14803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09311_ _09311_/A _11920_/B _11920_/C _09316_/B vssd1 vssd1 vccd1 vccd1 _14811_/C
+ sky130_fd_sc_hd__nor4_2
X_18509_ _20032_/CLK _18509_/D vssd1 vssd1 vccd1 vccd1 _18509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19489_ _19885_/CLK _19489_/D vssd1 vssd1 vccd1 vccd1 _19489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11532__S _11532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09242_ _09499_/B _09310_/C vssd1 vssd1 vccd1 vccd1 _11932_/A sky130_fd_sc_hd__or2_1
XFILLER_61_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09173_ _11961_/A _09282_/C vssd1 vssd1 vccd1 vccd1 _14756_/A sky130_fd_sc_hd__or2_2
XFILLER_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11411__A1 _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11768__A _15875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11714__A2 _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13983__A _13991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13467__A2 _13373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12599__A _12599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12675__A0 _15482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _10843_/X _10845_/X _09805_/A _10849_/X vssd1 vssd1 vccd1 vccd1 _10850_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _14782_/B _14766_/A _14782_/D vssd1 vssd1 vccd1 vccd1 _09510_/B sky130_fd_sc_hd__nor3_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10781_ _20021_/Q _19859_/Q _19268_/Q _19038_/Q _10776_/X _10710_/A vssd1 vssd1 vccd1
+ vccd1 _10781_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14319__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12493_/A _15397_/B _12497_/A _12497_/B vssd1 vssd1 vccd1 vccd1 _12521_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12452_/A _12483_/C vssd1 vssd1 vccd1 vccd1 _12451_/X sky130_fd_sc_hd__or2_1
XFILLER_40_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11402_ _20010_/Q _19848_/Q _19257_/Q _19027_/Q _11356_/X _11357_/X vssd1 vssd1 vccd1
+ vccd1 _11402_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15170_ _15168_/X _15072_/X _15298_/S vssd1 vssd1 vccd1 vccd1 _15170_/X sky130_fd_sc_hd__mux2_1
X_12382_ _15338_/A _12382_/B vssd1 vssd1 vccd1 vccd1 _12385_/A sky130_fd_sc_hd__xor2_2
XFILLER_166_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14121_ _18743_/Q _18742_/Q _18744_/Q _14521_/A vssd1 vssd1 vccd1 vccd1 _14126_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_153_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11333_ _20011_/Q _19849_/Q _19258_/Q _19028_/Q _11409_/S _11208_/A vssd1 vssd1 vccd1
+ vccd1 _11333_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14054__A _14745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ _14051_/B _14051_/C _18593_/Q vssd1 vssd1 vccd1 vccd1 _14053_/C sky130_fd_sc_hd__a21oi_1
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11264_ _11140_/A _11263_/X _09682_/A vssd1 vssd1 vccd1 vccd1 _11264_/X sky130_fd_sc_hd__o21a_1
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13003_ _13002_/X _18428_/Q _13003_/S vssd1 vssd1 vccd1 vccd1 _13004_/A sky130_fd_sc_hd__mux2_1
X_10215_ _10521_/A vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__buf_2
XFILLER_122_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18094__A1 _13661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18860_ _19025_/CLK _18860_/D vssd1 vssd1 vccd1 vccd1 _18860_/Q sky130_fd_sc_hd__dfxtp_4
X_11195_ _18837_/Q vssd1 vssd1 vccd1 vccd1 _11195_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17811_ _17867_/A vssd1 vssd1 vccd1 vccd1 _17880_/S sky130_fd_sc_hd__clkbuf_8
X_10146_ _11493_/A vssd1 vssd1 vccd1 vccd1 _10843_/A sky130_fd_sc_hd__buf_2
XANTENNA__17841__A1 _17036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ _19062_/CLK _18791_/D vssd1 vssd1 vccd1 vccd1 _18791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output143_A _12288_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11469__A1 _09664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17742_ _17742_/A vssd1 vssd1 vccd1 vccd1 _19751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10077_ _10077_/A vssd1 vssd1 vccd1 vccd1 _10078_/A sky130_fd_sc_hd__buf_4
X_14954_ _14952_/X _14953_/X _14957_/S vssd1 vssd1 vccd1 vccd1 _14954_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10677__C1 _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13905_ _18544_/Q _13900_/X _12699_/Y _12702_/Y _13904_/X vssd1 vssd1 vccd1 vccd1
+ _18544_/D sky130_fd_sc_hd__o221a_1
X_17673_ _17672_/X _19730_/Q _17682_/S vssd1 vssd1 vccd1 vccd1 _17674_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14885_ _14885_/A vssd1 vssd1 vccd1 vccd1 _15306_/B sky130_fd_sc_hd__clkbuf_2
X_19412_ _20003_/CLK _19412_/D vssd1 vssd1 vccd1 vccd1 _19412_/Q sky130_fd_sc_hd__dfxtp_1
X_16624_ _16304_/X _19289_/Q _16630_/S vssd1 vssd1 vccd1 vccd1 _16625_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15613__A _15624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ _18510_/Q _13835_/X _13836_/S vssd1 vssd1 vccd1 vccd1 _13837_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11316__S1 _11073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12956__B _12956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19343_ _20030_/CLK _19343_/D vssd1 vssd1 vccd1 vccd1 _19343_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09611__A _09636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16555_ _16555_/A vssd1 vssd1 vccd1 vccd1 _19258_/D sky130_fd_sc_hd__clkbuf_1
X_13767_ _13767_/A vssd1 vssd1 vccd1 vccd1 _18488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10979_ _19727_/Q vssd1 vssd1 vccd1 vccd1 _10979_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15506_ _15506_/A _15509_/A vssd1 vssd1 vccd1 vccd1 _15506_/X sky130_fd_sc_hd__or2_1
X_19274_ _19865_/CLK _19274_/D vssd1 vssd1 vccd1 vccd1 _19274_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15907__A1 _11452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ _18545_/Q _12719_/B vssd1 vssd1 vccd1 vccd1 _12720_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16486_ _19228_/Q _13771_/X _16486_/S vssd1 vssd1 vccd1 vccd1 _16487_/A sky130_fd_sc_hd__mux2_1
X_13698_ _13699_/A _13699_/B vssd1 vssd1 vccd1 vccd1 _13714_/C sky130_fd_sc_hd__or2_1
X_18225_ _18225_/A vssd1 vssd1 vccd1 vccd1 _19951_/D sky130_fd_sc_hd__clkbuf_1
X_15437_ _15159_/X _15432_/Y _15436_/Y vssd1 vssd1 vccd1 vccd1 _15438_/C sky130_fd_sc_hd__a21oi_1
XFILLER_129_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12649_ _12645_/X _12648_/Y _12770_/S vssd1 vssd1 vccd1 vccd1 _12649_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18156_ _17662_/X _19921_/Q _18158_/S vssd1 vssd1 vccd1 vccd1 _18157_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15368_ _15368_/A vssd1 vssd1 vccd1 vccd1 _15368_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17974__S _17976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17107_ _17106_/X _19492_/Q _17113_/S vssd1 vssd1 vccd1 vccd1 _17108_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11944__A2 _11438_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14319_ _14319_/A _14327_/C vssd1 vssd1 vccd1 vccd1 _14319_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10492__A _10492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18087_ _18104_/A vssd1 vssd1 vccd1 vccd1 _18101_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15299_ _15096_/X _15298_/X _15348_/S vssd1 vssd1 vccd1 vccd1 _15299_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17038_ _17038_/A vssd1 vssd1 vccd1 vccd1 _19466_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13146__B2 _13289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_74_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ _09929_/A _09860_/B vssd1 vssd1 vccd1 vccd1 _09860_/X sky130_fd_sc_hd__or2_1
XFILLER_124_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09996__S1 _09636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _09791_/A vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__clkbuf_2
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _18992_/CLK _18989_/D vssd1 vssd1 vccd1 vccd1 _18989_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12866__B _12866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09225_ _18964_/Q vssd1 vssd1 vccd1 vccd1 _09481_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14573__S _14581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11243__S0 _11158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10000_ _09849_/X _09982_/X _09999_/X _09540_/A _18858_/Q vssd1 vssd1 vccd1 vccd1
+ _15970_/C sky130_fd_sc_hd__a32o_4
XFILLER_49_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09989_ _10112_/A vssd1 vssd1 vccd1 vccd1 _10305_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18998__CLK _18998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13218__A _17042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11546__S1 _09614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11951_ _11951_/A _11951_/B vssd1 vssd1 vccd1 vccd1 _14812_/C sky130_fd_sc_hd__nor2_1
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10902_ _10905_/A _10901_/X _09792_/A vssd1 vssd1 vccd1 vccd1 _10902_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11882_ _12060_/B _14528_/A _11865_/X _11867_/X _11881_/X vssd1 vssd1 vccd1 vccd1
+ _18710_/D sky130_fd_sc_hd__o32a_1
X_14670_ _11801_/A _18789_/Q _14670_/S vssd1 vssd1 vccd1 vccd1 _14671_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09431__A _15624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10833_ _18435_/Q _19464_/Q _19501_/Q _19075_/Q _09650_/A _10049_/A vssd1 vssd1 vccd1
+ vccd1 _10833_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13621_ _13587_/X _13619_/X _13620_/Y _13590_/X _19008_/Q vssd1 vssd1 vccd1 vccd1
+ _13621_/X sky130_fd_sc_hd__a32o_4
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16340_ _16339_/X _19172_/Q _16346_/S vssd1 vssd1 vccd1 vccd1 _16341_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10764_ _19364_/Q _19699_/Q _10764_/S vssd1 vssd1 vccd1 vccd1 _10764_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13552_ _13589_/A _19000_/Q vssd1 vssd1 vccd1 vccd1 _13552_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12503_ _12503_/A vssd1 vssd1 vccd1 vccd1 _12697_/S sky130_fd_sc_hd__buf_2
X_16271_ _16282_/A vssd1 vssd1 vccd1 vccd1 _16280_/S sky130_fd_sc_hd__buf_4
X_13483_ _13483_/A vssd1 vssd1 vccd1 vccd1 _18454_/D sky130_fd_sc_hd__clkbuf_1
X_10695_ _10695_/A _10695_/B vssd1 vssd1 vccd1 vccd1 _10695_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18010_ _18010_/A vssd1 vssd1 vccd1 vccd1 _19871_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14573__A0 _12134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15222_ _15205_/X _15478_/B _15221_/X _15491_/A vssd1 vssd1 vccd1 vccd1 _15222_/X
+ sky130_fd_sc_hd__a211o_1
X_12434_ _14966_/A _12458_/A vssd1 vssd1 vccd1 vccd1 _12435_/B sky130_fd_sc_hd__nor2_2
XANTENNA__10809__S0 _10797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13099__S _13116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12365_ _18531_/Q vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__clkbuf_2
X_15153_ _15171_/S _15152_/X _15097_/X vssd1 vssd1 vccd1 vccd1 _15153_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11316_ _19657_/Q _19423_/Q _18488_/Q _19753_/Q _11124_/A _11073_/A vssd1 vssd1 vccd1
+ vccd1 _11317_/B sky130_fd_sc_hd__mux4_1
X_14104_ _14105_/B _14105_/C _14103_/Y vssd1 vssd1 vccd1 vccd1 _18610_/D sky130_fd_sc_hd__o21a_1
XFILLER_153_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19961_ _20025_/CLK _19961_/D vssd1 vssd1 vccd1 vccd1 _19961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15084_ _15077_/X _15078_/Y _15083_/X _14855_/A vssd1 vssd1 vccd1 vccd1 _15084_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_141_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12296_ _12295_/Y _18908_/Q _12409_/A vssd1 vssd1 vccd1 vccd1 _14859_/A sky130_fd_sc_hd__mux2_4
XFILLER_141_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13679__A2 _13517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13827__S _13836_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18067__A1 _11833_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14035_ _14034_/B _14034_/C _18587_/Q vssd1 vssd1 vccd1 vccd1 _14036_/C sky130_fd_sc_hd__a21oi_1
X_18912_ _19010_/CLK _18912_/D vssd1 vssd1 vccd1 vccd1 _18912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11247_ _19197_/Q _19788_/Q _19950_/Q _19165_/Q _11273_/A _11073_/X vssd1 vssd1 vccd1
+ vccd1 _11248_/B sky130_fd_sc_hd__mux4_1
X_19892_ _19896_/CLK _19892_/D vssd1 vssd1 vccd1 vccd1 _19892_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14512__A _14528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18843_ _19324_/CLK _18843_/D vssd1 vssd1 vccd1 vccd1 _18843_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11855__B _11855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _19917_/Q _19531_/Q _19981_/Q _19100_/Q _11171_/X _11172_/X vssd1 vssd1 vccd1
+ vccd1 _11179_/B sky130_fd_sc_hd__mux4_1
XANTENNA__14628__A1 _13667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10129_ _19379_/Q _19714_/Q _10129_/S vssd1 vssd1 vccd1 vccd1 _10129_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10251__S _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17823__A _17880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18774_ _19900_/CLK _18774_/D vssd1 vssd1 vccd1 vccd1 _18774_/Q sky130_fd_sc_hd__dfxtp_2
X_15986_ _16150_/B _16691_/B _15735_/A vssd1 vssd1 vccd1 vccd1 _18352_/C sky130_fd_sc_hd__or3b_4
X_17725_ _17725_/A vssd1 vssd1 vccd1 vccd1 _19746_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11537__S1 _09639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14937_ _15424_/B _15291_/B _14937_/S vssd1 vssd1 vccd1 vccd1 _14937_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17034__S _17040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11862__A1 _18711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17656_ _17656_/A vssd1 vssd1 vccd1 vccd1 _17656_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14868_ _14868_/A vssd1 vssd1 vccd1 vccd1 _15254_/B sky130_fd_sc_hd__buf_2
X_16607_ _19282_/Q _13842_/X _16613_/S vssd1 vssd1 vccd1 vccd1 _16608_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13819_ _17055_/A vssd1 vssd1 vccd1 vccd1 _13819_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16873__S _16881_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17587_ _17131_/X _19697_/Q _17595_/S vssd1 vssd1 vccd1 vccd1 _17588_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14799_ _14813_/A _15747_/A _14778_/A _18832_/Q vssd1 vssd1 vccd1 vccd1 _14800_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19326_ _19951_/CLK _19326_/D vssd1 vssd1 vccd1 vccd1 _19326_/Q sky130_fd_sc_hd__dfxtp_1
X_16538_ _16538_/A vssd1 vssd1 vccd1 vccd1 _19251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19257_ _19946_/CLK _19257_/D vssd1 vssd1 vccd1 vccd1 _19257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16469_ _16469_/A vssd1 vssd1 vccd1 vccd1 _19221_/D sky130_fd_sc_hd__clkbuf_1
X_18208_ _18208_/A _18208_/B vssd1 vssd1 vccd1 vccd1 _18265_/A sky130_fd_sc_hd__nor2_4
XFILLER_164_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19188_ _19973_/CLK _19188_/D vssd1 vssd1 vccd1 vccd1 _19188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18139_ _17634_/X _19913_/Q _18147_/S vssd1 vssd1 vccd1 vccd1 _18140_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13310__B _13451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15108__A2 _15100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09912_ _09912_/A vssd1 vssd1 vccd1 vccd1 _09913_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20032_ _20032_/CLK _20032_/D vssd1 vssd1 vccd1 vccd1 _20032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09843_ _09843_/A vssd1 vssd1 vccd1 vccd1 _09843_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10889__C1 _09550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11765__B _13910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14619__A1 _11748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _09774_/A vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__buf_2
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12877__A _13070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10397__A _15962_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13055__B1 _13053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10813__C1 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09208_ _14804_/A vssd1 vssd1 vccd1 vccd1 _14782_/A sky130_fd_sc_hd__buf_6
X_10480_ _10480_/A _10480_/B vssd1 vssd1 vccd1 vccd1 _10480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12150_ _12150_/A _12184_/A vssd1 vssd1 vccd1 vccd1 _12150_/Y sky130_fd_sc_hd__xnor2_4
X_11101_ _11088_/Y _11096_/Y _11098_/Y _11100_/Y _09817_/A vssd1 vssd1 vccd1 vccd1
+ _11101_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11956__A _11956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _12085_/A vssd1 vssd1 vccd1 vccd1 _12537_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16023__S _16031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14332__A _14427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11032_ _11032_/A _11032_/B vssd1 vssd1 vccd1 vccd1 _11032_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16958__S _16964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15840_ _15871_/A _15840_/B vssd1 vssd1 vccd1 vccd1 _18975_/D sky130_fd_sc_hd__nor2_1
XFILLER_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _20016_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _18954_/Q _15775_/B vssd1 vssd1 vccd1 vccd1 _15771_/X sky130_fd_sc_hd__or2_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12983_ _19885_/Q _11845_/X _13511_/A _18458_/Q vssd1 vssd1 vccd1 vccd1 _12983_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13294__B1 _13082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11691__A _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17510_ _19661_/Q vssd1 vssd1 vccd1 vccd1 _17511_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _14722_/A vssd1 vssd1 vccd1 vccd1 _18811_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _15740_/A _11663_/A _09437_/A _09280_/Y vssd1 vssd1 vccd1 vccd1 _12315_/A
+ sky130_fd_sc_hd__a211o_1
X_18490_ _19949_/CLK _18490_/D vssd1 vssd1 vccd1 vccd1 _18490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17789__S _17793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17441_ _17441_/A vssd1 vssd1 vccd1 vccd1 _19628_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ _12750_/B _13719_/X _14667_/S vssd1 vssd1 vccd1 vccd1 _14654_/B sky130_fd_sc_hd__mux2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _11865_/A vssd1 vssd1 vccd1 vccd1 _11865_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output106_A _14782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _13603_/A _13603_/C _13174_/A vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__o21ai_1
X_10816_ _15938_/C _12841_/A vssd1 vssd1 vccd1 vccd1 _10818_/A sky130_fd_sc_hd__nand2_1
X_17372_ _19598_/Q _17017_/X _17376_/S vssd1 vssd1 vccd1 vccd1 _17373_/A sky130_fd_sc_hd__mux2_1
X_14584_ _14601_/A vssd1 vssd1 vccd1 vccd1 _14598_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_14_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11796_ _11796_/A _11796_/B _11796_/C vssd1 vssd1 vccd1 vccd1 _11796_/X sky130_fd_sc_hd__or3_4
XFILLER_41_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19111_ _20024_/CLK _19111_/D vssd1 vssd1 vccd1 vccd1 _19111_/Q sky130_fd_sc_hd__dfxtp_1
X_16323_ _17659_/A vssd1 vssd1 vccd1 vccd1 _16323_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13535_ _13535_/A _13535_/B vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__nand2_1
X_10747_ _19669_/Q _19435_/Q _18500_/Q _19765_/Q _09725_/A _10626_/A vssd1 vssd1 vccd1
+ vccd1 _10748_/B sky130_fd_sc_hd__mux4_1
XFILLER_13_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19042_ _20026_/CLK _19042_/D vssd1 vssd1 vccd1 vccd1 _19042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16254_ _13161_/X _19140_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _16255_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ _09849_/A _10668_/X _10677_/X _09539_/A _18848_/Q vssd1 vssd1 vccd1 vccd1
+ _15947_/C sky130_fd_sc_hd__a32o_4
X_13466_ _19911_/Q vssd1 vssd1 vccd1 vccd1 _13466_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15205_ _15365_/A vssd1 vssd1 vccd1 vccd1 _15205_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12417_ _12368_/A _12416_/B _12416_/D _12416_/C vssd1 vssd1 vccd1 vccd1 _12417_/X
+ sky130_fd_sc_hd__a31o_1
X_16185_ _16185_/A vssd1 vssd1 vccd1 vccd1 _19110_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10258__S1 _09637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12027__A _18520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13397_ _18816_/Q _13269_/X _12879_/X _18783_/Q _13396_/X vssd1 vssd1 vccd1 vccd1
+ _13397_/X sky130_fd_sc_hd__a221o_1
XFILLER_154_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15136_ _14923_/X _15122_/X _14984_/X vssd1 vssd1 vccd1 vccd1 _15136_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12348_ _12349_/A _12374_/C vssd1 vssd1 vccd1 vccd1 _12348_/X sky130_fd_sc_hd__or2_1
XFILLER_142_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11866__A _15719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15338__A _15338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19944_ _20040_/CLK _19944_/D vssd1 vssd1 vccd1 vccd1 _19944_/Q sky130_fd_sc_hd__dfxtp_1
X_12279_ _12279_/A _12279_/B _12279_/C _12279_/D vssd1 vssd1 vccd1 vccd1 _12279_/X
+ sky130_fd_sc_hd__or4_1
X_15067_ _15064_/X _15066_/X _15280_/S vssd1 vssd1 vccd1 vccd1 _15067_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14018_ _18580_/Q _14016_/B _14017_/Y vssd1 vssd1 vccd1 vccd1 _18580_/D sky130_fd_sc_hd__o21a_1
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19875_ _20037_/CLK _19875_/D vssd1 vssd1 vccd1 vccd1 _19875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18826_ _18960_/CLK _18826_/D vssd1 vssd1 vccd1 vccd1 _18826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10430__S1 _10163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18757_ _19063_/CLK _18757_/D vssd1 vssd1 vccd1 vccd1 _18757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15969_ _19018_/Q _15954_/X _15955_/X _15968_/Y vssd1 vssd1 vccd1 vccd1 _19018_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17708_ _17707_/X _19741_/Q _17714_/S vssd1 vssd1 vccd1 vccd1 _17709_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09490_ _19485_/Q vssd1 vssd1 vccd1 vccd1 _09909_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18688_ _18688_/CLK _18688_/D vssd1 vssd1 vccd1 vccd1 _18688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13037__A0 _18839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17639_ _17639_/A vssd1 vssd1 vccd1 vccd1 _19719_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11106__A _19385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10010__A _10010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19309_ _19644_/CLK _19309_/D vssd1 vssd1 vccd1 vccd1 _19309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11446__S0 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16632__A _16689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09811__S0 _09898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16778__S _16786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20015_ _20015_/CLK _20015_/D vssd1 vssd1 vccd1 vccd1 _20015_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13991__A _13991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09826_ _09826_/A _09826_/B vssd1 vssd1 vccd1 vccd1 _09826_/X sky130_fd_sc_hd__and2_1
XFILLER_24_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09757_ _10947_/A vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13276__B1 _12890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16079__A _16135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _10192_/A vssd1 vssd1 vccd1 vccd1 _09980_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11650_ _11578_/X _11579_/Y _11580_/Y _11530_/X _11649_/X vssd1 vssd1 vccd1 vccd1
+ _11650_/X sky130_fd_sc_hd__a221o_4
XANTENNA__11039__C1 _11166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13579__B2 _19003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10601_ _10727_/A vssd1 vssd1 vccd1 vccd1 _10836_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11581_ _11581_/A vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__inv_2
XFILLER_167_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16018__S _16020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10855__A _10893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13231__A _13340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10532_ _19146_/Q _19407_/Q _19306_/Q _19641_/Q _10216_/A _10218_/A vssd1 vssd1 vccd1
+ vccd1 _10532_/X sky130_fd_sc_hd__mux4_1
X_13320_ input14/X _13318_/X _13319_/X vssd1 vssd1 vccd1 vccd1 _13320_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10463_ _20028_/Q _19866_/Q _19275_/Q _19045_/Q _10314_/S _10400_/A vssd1 vssd1 vccd1
+ vccd1 _10463_/X sky130_fd_sc_hd__mux4_1
X_13251_ _13250_/X _18441_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _13252_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18233__S _18241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09955__B1 _09837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ _12255_/C _12201_/Y _12366_/B vssd1 vssd1 vccd1 vccd1 _12202_/Y sky130_fd_sc_hd__o21ai_1
X_13182_ _13182_/A vssd1 vssd1 vccd1 vccd1 _18437_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11211__C1 _11133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10394_ _10335_/A _10393_/X _10382_/X vssd1 vssd1 vccd1 vccd1 _10394_/X sky130_fd_sc_hd__o21a_1
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input67_A io_irq_motor_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_142_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18719_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12133_ _18762_/Q vssd1 vssd1 vccd1 vccd1 _12165_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11686__A _11686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _19862_/Q _17042_/X _17998_/S vssd1 vssd1 vccd1 vccd1 _17991_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12064_ _12064_/A _12064_/B vssd1 vssd1 vccd1 vccd1 _12161_/B sky130_fd_sc_hd__nor2_2
X_16941_ _16941_/A vssd1 vssd1 vccd1 vccd1 _19429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11015_ _11015_/A vssd1 vssd1 vccd1 vccd1 _11015_/X sky130_fd_sc_hd__buf_2
X_19660_ _20016_/CLK _19660_/D vssd1 vssd1 vccd1 vccd1 _19660_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10412__S1 _10320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16872_ _16918_/S vssd1 vssd1 vccd1 vccd1 _16881_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10868__A2 _10850_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_157_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19896_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18611_ _18724_/CLK _18611_/D vssd1 vssd1 vccd1 vccd1 _18611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15823_ _15823_/A vssd1 vssd1 vccd1 vccd1 _18969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19591_ _19816_/CLK _19591_/D vssd1 vssd1 vccd1 vccd1 _19591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18542_ _18548_/CLK _18542_/D vssd1 vssd1 vccd1 vccd1 _18542_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _12032_/X _15752_/X _15753_/X _15743_/X vssd1 vssd1 vccd1 vccd1 _18947_/D
+ sky130_fd_sc_hd__o211a_1
X_12966_ _19487_/Q vssd1 vssd1 vccd1 vccd1 _13297_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14705_ _18804_/Q _13621_/X _14705_/S vssd1 vssd1 vccd1 vccd1 _14706_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _18518_/Q _13861_/C vssd1 vssd1 vccd1 vccd1 _11918_/A sky130_fd_sc_hd__and2_4
X_18473_ _18547_/CLK _18473_/D vssd1 vssd1 vccd1 vccd1 _18473_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _15685_/A vssd1 vssd1 vccd1 vccd1 _18919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12897_ _12957_/A vssd1 vssd1 vccd1 vccd1 _12897_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13840__S _13852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ _19622_/Q _17093_/X _17424_/S vssd1 vssd1 vccd1 vccd1 _17425_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14636_ _18779_/Q _13685_/X _14649_/S vssd1 vssd1 vccd1 vccd1 _14637_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11848_ _18466_/Q _12943_/A _11772_/A _18713_/Q vssd1 vssd1 vccd1 vccd1 _11848_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09869__S0 _09635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17355_ _17411_/A vssd1 vssd1 vccd1 vccd1 _17424_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14567_ _12020_/X _13508_/B _14581_/S vssd1 vssd1 vccd1 vccd1 _14568_/B sky130_fd_sc_hd__mux2_1
X_11779_ _12060_/A _11705_/A _11783_/C _15760_/A vssd1 vssd1 vccd1 vccd1 _12878_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16306_ _16306_/A vssd1 vssd1 vccd1 vccd1 _19161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13518_ _13518_/A vssd1 vssd1 vccd1 vccd1 _13689_/S sky130_fd_sc_hd__clkbuf_4
X_17286_ _17286_/A vssd1 vssd1 vccd1 vccd1 _19559_/D sky130_fd_sc_hd__clkbuf_1
X_14498_ _18732_/Q _14495_/B _14497_/Y vssd1 vssd1 vccd1 vccd1 _18732_/D sky130_fd_sc_hd__o21a_1
XFILLER_174_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19025_ _19025_/CLK _19025_/D vssd1 vssd1 vccd1 vccd1 _19025_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__17548__A _19680_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16237_ _16237_/A vssd1 vssd1 vccd1 vccd1 _19132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13449_ _18894_/Q _13449_/B vssd1 vssd1 vccd1 vccd1 _13476_/B sky130_fd_sc_hd__and2_1
XANTENNA__18143__S _18147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13742__A1 _13531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18130__A0 _18863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16168_ _16168_/A vssd1 vssd1 vccd1 vccd1 _19102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11753__B1 _11687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15119_ _15117_/X _15118_/X _15189_/S vssd1 vssd1 vccd1 vccd1 _15119_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16099_ _16099_/A vssd1 vssd1 vccd1 vccd1 _19072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19927_ _20023_/CLK _19927_/D vssd1 vssd1 vccd1 vccd1 _19927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16598__S _16602_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17283__A _17339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10403__S1 _10320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19858_ _19990_/CLK _19858_/D vssd1 vssd1 vccd1 vccd1 _19858_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10005__A _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ _09636_/A vssd1 vssd1 vccd1 vccd1 _09612_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18809_ _19900_/CLK _18809_/D vssd1 vssd1 vccd1 vccd1 _18809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19789_ _19855_/CLK _19789_/D vssd1 vssd1 vccd1 vccd1 _19789_/Q sky130_fd_sc_hd__dfxtp_1
X_09542_ _09542_/A _09542_/B _09542_/C _09303_/X vssd1 vssd1 vccd1 vccd1 _10077_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_110_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09477__A2 _09433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09473_ _09514_/A _12055_/C vssd1 vssd1 vccd1 vccd1 _12004_/C sky130_fd_sc_hd__or2_1
XANTENNA__12481__A1 _18471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18318__S _18324_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15250__B _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11270__S _11270_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14581__S _14581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12890__A _12890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09937__B1 _09540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18121__A0 _18860_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10642__S1 _10626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _20039_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09809_ _09809_/A vssd1 vssd1 vccd1 vccd1 _09809_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_89_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 _19581_/CLK sky130_fd_sc_hd__clkbuf_16
X_12820_ _12820_/A _12820_/B vssd1 vssd1 vccd1 vccd1 _12820_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10158__S0 _10328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12530_/X _12749_/Y _12774_/B _12583_/X vssd1 vssd1 vccd1 vccd1 _12751_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_15_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18228__S _18230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _18773_/Q vssd1 vssd1 vccd1 vccd1 _12452_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19757_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15474_/A _15474_/B vssd1 vssd1 vccd1 vccd1 _15470_/Y sky130_fd_sc_hd__nand2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12682_/A vssd1 vssd1 vccd1 vccd1 _12778_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _14479_/A vssd1 vssd1 vccd1 vccd1 _14472_/A sky130_fd_sc_hd__buf_2
XFILLER_70_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11633_ _11633_/A _11633_/B _11633_/C vssd1 vssd1 vccd1 vccd1 _11633_/X sky130_fd_sc_hd__or3_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15160__B _15160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16971__S _16975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13421__B1 _13420_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__A _15952_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17140_ _17140_/A vssd1 vssd1 vccd1 vccd1 _19502_/D sky130_fd_sc_hd__clkbuf_1
X_14352_ _14355_/B _14355_/C _14332_/X vssd1 vssd1 vccd1 vccd1 _14352_/Y sky130_fd_sc_hd__a21oi_1
X_11564_ _19383_/Q _19718_/Q _11566_/S vssd1 vssd1 vccd1 vccd1 _11565_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ _13386_/A vssd1 vssd1 vccd1 vccd1 _13366_/S sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_27_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19853_/CLK sky130_fd_sc_hd__clkbuf_16
X_10515_ _19931_/Q _19545_/Q _19995_/Q _19114_/Q _10216_/A _10218_/A vssd1 vssd1 vccd1
+ vccd1 _10516_/B sky130_fd_sc_hd__mux4_1
X_17071_ _17071_/A vssd1 vssd1 vccd1 vccd1 _17071_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11495_ _11500_/A _11495_/B vssd1 vssd1 vccd1 vccd1 _11495_/X sky130_fd_sc_hd__or2_1
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14283_ _14290_/D _14283_/B vssd1 vssd1 vccd1 vccd1 _18660_/D sky130_fd_sc_hd__nor2_1
XFILLER_109_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16022_ _16044_/A vssd1 vssd1 vccd1 vccd1 _16031_/S sky130_fd_sc_hd__clkbuf_4
X_10446_ _19674_/Q _19440_/Q _18505_/Q _19770_/Q _10319_/X _10320_/X vssd1 vssd1 vccd1
+ vccd1 _10446_/X sky130_fd_sc_hd__mux4_1
X_13234_ _13319_/A vssd1 vssd1 vccd1 vccd1 _13234_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output173_A _12259_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10377_ _18445_/Q _19474_/Q _19511_/Q _19085_/Q _10209_/S _10163_/X vssd1 vssd1 vccd1
+ vccd1 _10377_/X sky130_fd_sc_hd__mux4_2
X_13165_ _18467_/Q _12982_/A _11847_/A _18691_/Q _13164_/X vssd1 vssd1 vccd1 vccd1
+ _13165_/X sky130_fd_sc_hd__a221o_1
XFILLER_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14223__C _18940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12116_ _12080_/B _12143_/A _12029_/A vssd1 vssd1 vccd1 vccd1 _12117_/B sky130_fd_sc_hd__o21ai_1
XFILLER_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17973_ _17973_/A vssd1 vssd1 vccd1 vccd1 _19854_/D sky130_fd_sc_hd__clkbuf_1
X_13096_ _09532_/X _13090_/X _13095_/X vssd1 vssd1 vccd1 vccd1 _17020_/A sky130_fd_sc_hd__o21a_4
XFILLER_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19712_ _19971_/CLK _19712_/D vssd1 vssd1 vccd1 vccd1 _19712_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17307__S _17315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16924_ _16924_/A vssd1 vssd1 vccd1 vccd1 _19421_/D sky130_fd_sc_hd__clkbuf_1
X_12047_ _18521_/Q _12583_/A vssd1 vssd1 vccd1 vccd1 _12076_/A sky130_fd_sc_hd__or2_1
XANTENNA__16211__S _16217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14520__A _14528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09614__A _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19643_ _19996_/CLK _19643_/D vssd1 vssd1 vccd1 vccd1 _19643_/Q sky130_fd_sc_hd__dfxtp_1
X_16855_ _16307_/X _19391_/Q _16859_/S vssd1 vssd1 vccd1 vccd1 _16856_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15335__B _15338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13136__A _17026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15806_ _15805_/Y _15834_/A _15789_/A _09436_/C vssd1 vssd1 vccd1 vccd1 _15807_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19574_ _19828_/CLK _19574_/D vssd1 vssd1 vccd1 vccd1 _19574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16786_ _16329_/X _19361_/Q _16786_/S vssd1 vssd1 vccd1 vccd1 _16787_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13998_ _18573_/Q _13999_/C _18574_/Q vssd1 vssd1 vccd1 vccd1 _14000_/B sky130_fd_sc_hd__a21oi_1
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18525_ _18867_/CLK _18525_/D vssd1 vssd1 vccd1 vccd1 _18525_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15737_ hold4/X _15734_/X _15736_/X _15730_/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__o211a_1
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12949_ _18456_/Q _12943_/X _12944_/X _14350_/B _12948_/X vssd1 vssd1 vccd1 vccd1
+ _12949_/X sky130_fd_sc_hd__a221o_1
XFILLER_34_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18456_ _18994_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15668_ _15690_/A vssd1 vssd1 vccd1 vccd1 _15677_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_60_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17407_ _19614_/Q _17068_/X _17409_/S vssd1 vssd1 vccd1 vccd1 _17408_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14619_ _18774_/Q _11748_/X _14632_/S vssd1 vssd1 vccd1 vccd1 _14620_/B sky130_fd_sc_hd__mux2_1
XANTENNA__16881__S _16881_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18387_ _18409_/A vssd1 vssd1 vccd1 vccd1 _18396_/S sky130_fd_sc_hd__buf_4
XFILLER_33_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15599_ _15599_/A vssd1 vssd1 vccd1 vccd1 _18881_/D sky130_fd_sc_hd__clkbuf_1
X_17338_ _17338_/A vssd1 vssd1 vccd1 vccd1 _19583_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10321__S0 _10319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17269_ _17269_/A vssd1 vssd1 vccd1 vccd1 _19552_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19008_ _19010_/CLK _19008_/D vssd1 vssd1 vccd1 vccd1 _19008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_144_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13191__A2 _13511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15468__A1 _12621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17217__S _17221_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15640__A1 _18520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09525_ _09525_/A _14822_/B _12845_/A _09525_/D vssd1 vssd1 vccd1 vccd1 _09525_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__12454__A1 _12446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14576__S _14581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12454__B2 _12453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_69_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09456_/A vssd1 vssd1 vccd1 vccd1 _14756_/B sky130_fd_sc_hd__clkbuf_2
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17887__S _17893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16791__S _16797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ _18958_/Q vssd1 vssd1 vccd1 vccd1 _15779_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12206__B2 _18989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10863__S1 _10788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10300_ _15966_/C _12855_/B vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__or2_1
XFILLER_4_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11280_ _11070_/X _11279_/X _09682_/A vssd1 vssd1 vccd1 vccd1 _11280_/X sky130_fd_sc_hd__o21a_1
XFILLER_146_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10231_ _10344_/A _10231_/B vssd1 vssd1 vccd1 vccd1 _10231_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11667__C _11667_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10162_ _10162_/A vssd1 vssd1 vccd1 vccd1 _10162_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_126_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10940__B2 _09550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15436__A _15436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16031__S _16031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10093_ _10093_/A _10093_/B vssd1 vssd1 vccd1 vccd1 _10093_/Y sky130_fd_sc_hd__nor2_1
X_14970_ _15552_/A _14970_/B _14970_/C _14970_/D vssd1 vssd1 vccd1 vccd1 _14970_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__14340__A _14413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10379__S0 _10209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13921_ _18611_/Q _18610_/Q _18612_/Q _14099_/A vssd1 vssd1 vccd1 vccd1 _13929_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16640_ _16640_/A vssd1 vssd1 vccd1 vccd1 _19296_/D sky130_fd_sc_hd__clkbuf_1
X_13852_ _18515_/Q _13851_/X _13852_/S vssd1 vssd1 vccd1 vccd1 _13853_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12803_ _12316_/A _15916_/A _12866_/C _11904_/X vssd1 vssd1 vccd1 vccd1 _15553_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_56_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16571_ _16617_/S vssd1 vssd1 vccd1 vccd1 _16580_/S sky130_fd_sc_hd__clkbuf_4
X_13783_ _13783_/A vssd1 vssd1 vccd1 vccd1 _18493_/D sky130_fd_sc_hd__clkbuf_1
X_10995_ _11409_/S vssd1 vssd1 vccd1 vccd1 _10995_/X sky130_fd_sc_hd__clkbuf_4
X_18310_ _18310_/A vssd1 vssd1 vccd1 vccd1 _19989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ _15522_/A _15522_/B _15522_/C vssd1 vssd1 vccd1 vccd1 _15522_/X sky130_fd_sc_hd__and3_1
X_19290_ _19979_/CLK _19290_/D vssd1 vssd1 vccd1 vccd1 _19290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12734_ _09471_/C _12657_/X _12778_/A _12733_/Y vssd1 vssd1 vccd1 vccd1 _15520_/A
+ sky130_fd_sc_hd__a211o_2
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _19959_/Q _17681_/A _18241_/S vssd1 vssd1 vccd1 vccd1 _18242_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15419_/X _15248_/X _15452_/X _15428_/X vssd1 vssd1 vccd1 vccd1 _15453_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12665_ _12667_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _12666_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _18697_/Q vssd1 vssd1 vccd1 vccd1 _14411_/C sky130_fd_sc_hd__clkbuf_1
X_18172_ _17684_/X _19928_/Q _18180_/S vssd1 vssd1 vccd1 vccd1 _18173_/A sky130_fd_sc_hd__mux2_1
X_11616_ _11616_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11616_/X sky130_fd_sc_hd__or2_1
XFILLER_129_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15384_ _15384_/A vssd1 vssd1 vccd1 vccd1 _15384_/X sky130_fd_sc_hd__clkbuf_2
X_12596_ _12545_/A _12572_/A _12572_/B vssd1 vssd1 vccd1 vccd1 _12596_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_129_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17123_ _17122_/X _19497_/Q _17129_/S vssd1 vssd1 vccd1 vccd1 _17124_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17098__A _17098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14335_ _14336_/B _14338_/D _18676_/Q vssd1 vssd1 vccd1 vccd1 _14337_/B sky130_fd_sc_hd__a21oi_1
XFILLER_11_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11547_ _11547_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _11547_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16206__S _16206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09609__A _10492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17054_ _17054_/A vssd1 vssd1 vccd1 vccd1 _19471_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output98_A _12124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14266_ _18656_/Q _14262_/B _14265_/Y vssd1 vssd1 vccd1 vccd1 _18656_/D sky130_fd_sc_hd__o21a_1
XANTENNA__11858__B _19006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11478_ _18437_/Q _19466_/Q _19503_/Q _19077_/Q _10708_/X _10710_/X vssd1 vssd1 vccd1
+ vccd1 _11478_/X sky130_fd_sc_hd__mux4_2
XFILLER_125_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16005_ _13065_/X _19033_/Q _16009_/S vssd1 vssd1 vccd1 vccd1 _16006_/A sky130_fd_sc_hd__mux2_1
X_13217_ _13217_/A _13217_/B vssd1 vssd1 vccd1 vccd1 _17042_/A sky130_fd_sc_hd__and2_4
X_10429_ _10434_/A _10429_/B vssd1 vssd1 vccd1 vccd1 _10429_/Y sky130_fd_sc_hd__nor2_1
X_14197_ _18638_/Q _18637_/Q _14197_/C vssd1 vssd1 vccd1 vccd1 _14200_/B sky130_fd_sc_hd__and3_1
XFILLER_124_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12381__B1 _12459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _09532_/X _13146_/X _13147_/X vssd1 vssd1 vccd1 vccd1 _17030_/A sky130_fd_sc_hd__o21a_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17037__S _17040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14250__A _14265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17956_ _18024_/S vssd1 vssd1 vccd1 vccd1 _17965_/S sky130_fd_sc_hd__clkbuf_4
X_13079_ _18590_/Q _13120_/A _11687_/X _14153_/B vssd1 vssd1 vccd1 vccd1 _13079_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12689__B _12715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16907_ _16907_/A vssd1 vssd1 vccd1 vccd1 _19414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17887_ _19816_/Q _16998_/X _17893_/S vssd1 vssd1 vccd1 vccd1 _17888_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12684__A1 _09261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13881__B1 _14447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19626_ _19980_/CLK _19626_/D vssd1 vssd1 vccd1 vccd1 _19626_/Q sky130_fd_sc_hd__dfxtp_1
X_16838_ _16838_/A vssd1 vssd1 vccd1 vccd1 _19384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19557_ _20007_/CLK _19557_/D vssd1 vssd1 vccd1 vccd1 _19557_/Q sky130_fd_sc_hd__dfxtp_1
X_16769_ _16304_/X _19353_/Q _16775_/S vssd1 vssd1 vccd1 vccd1 _16770_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13633__A0 _13629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09310_ _09521_/A _09316_/A _09310_/C vssd1 vssd1 vccd1 vccd1 _14811_/B sky130_fd_sc_hd__nor3_1
X_18508_ _19935_/CLK _18508_/D vssd1 vssd1 vccd1 vccd1 _18508_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_70_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19488_ _19488_/CLK _19488_/D vssd1 vssd1 vccd1 vccd1 _19488_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09241_ _09290_/B vssd1 vssd1 vccd1 vccd1 _09310_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18439_ _20026_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09172_ _09283_/B _09283_/D _09285_/C vssd1 vssd1 vccd1 vccd1 _09282_/C sky130_fd_sc_hd__or3b_1
XFILLER_147_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18331__S _18335_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10922__A1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14160__A _14427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09254__A _18990_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16786__S _16786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10686__B1 _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10781__S0 _10776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12427__A1 _12416_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09508_ _09508_/A _09508_/B _09508_/C vssd1 vssd1 vccd1 vccd1 _14782_/D sky130_fd_sc_hd__nand3_1
XANTENNA__13504__A _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10886_/A _10780_/B vssd1 vssd1 vccd1 vccd1 _10780_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _15393_/A vssd1 vssd1 vccd1 vccd1 _15517_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12450_ _12338_/X _12448_/X _12449_/Y vssd1 vssd1 vccd1 vccd1 _12450_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11401_ _11401_/A _11401_/B vssd1 vssd1 vccd1 vccd1 _11401_/X sky130_fd_sc_hd__or2_1
XANTENNA__11959__A _14931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ _15306_/A _12406_/B _15321_/A _12459_/A vssd1 vssd1 vccd1 vccd1 _12382_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_165_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16877__A0 _16339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ _18739_/Q _18741_/Q _18740_/Q _14513_/A vssd1 vssd1 vccd1 vccd1 _14521_/A
+ sky130_fd_sc_hd__and4_1
X_11332_ _11332_/A _11332_/B vssd1 vssd1 vccd1 vccd1 _11332_/X sky130_fd_sc_hd__or2_1
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14352__A1 _14355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14051_ _18593_/Q _14051_/B _14051_/C vssd1 vssd1 vccd1 vccd1 _14053_/B sky130_fd_sc_hd__and3_1
XFILLER_107_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11263_ _19325_/Q _19596_/Q _19820_/Q _19564_/Q _11367_/S _10996_/A vssd1 vssd1 vccd1
+ vccd1 _11263_/X sky130_fd_sc_hd__mux4_1
XANTENNA__18241__S _18241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13002_ _17649_/A vssd1 vssd1 vccd1 vccd1 _13002_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10214_ _10520_/A vssd1 vssd1 vccd1 vccd1 _10480_/A sky130_fd_sc_hd__buf_2
X_11194_ _11095_/X _11185_/Y _11189_/Y _11193_/Y _09803_/A vssd1 vssd1 vccd1 vccd1
+ _11194_/X sky130_fd_sc_hd__o311a_1
XFILLER_161_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10145_ _10947_/A vssd1 vssd1 vccd1 vccd1 _11493_/A sky130_fd_sc_hd__clkbuf_2
X_17810_ _18208_/B _17954_/B vssd1 vssd1 vccd1 vccd1 _17867_/A sky130_fd_sc_hd__nor2_4
X_18790_ _19062_/CLK _18790_/D vssd1 vssd1 vccd1 vccd1 _18790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17741_ _17634_/X _19751_/Q _17749_/S vssd1 vssd1 vccd1 vccd1 _17742_/A sky130_fd_sc_hd__mux2_1
X_10076_ _10069_/Y _10071_/Y _10073_/Y _10075_/Y _09555_/A vssd1 vssd1 vccd1 vccd1
+ _10076_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14953_ _12783_/A _14996_/B _14955_/S vssd1 vssd1 vccd1 vccd1 _14953_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13904_ _13910_/A vssd1 vssd1 vccd1 vccd1 _13904_/X sky130_fd_sc_hd__buf_2
X_17672_ _17672_/A vssd1 vssd1 vccd1 vccd1 _17672_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14884_ _15321_/B _15397_/B _14908_/S vssd1 vssd1 vccd1 vccd1 _14884_/X sky130_fd_sc_hd__mux2_1
X_19411_ _19999_/CLK _19411_/D vssd1 vssd1 vccd1 vccd1 _19411_/Q sky130_fd_sc_hd__dfxtp_1
X_16623_ _16623_/A vssd1 vssd1 vccd1 vccd1 _19288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13835_ _17071_/A vssd1 vssd1 vccd1 vccd1 _13835_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19342_ _19999_/CLK _19342_/D vssd1 vssd1 vccd1 vccd1 _19342_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16554_ _19258_/Q _13765_/X _16558_/S vssd1 vssd1 vccd1 vccd1 _16555_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13766_ _18488_/Q _13765_/X _13772_/S vssd1 vssd1 vccd1 vccd1 _13767_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ _10978_/A _10978_/B vssd1 vssd1 vccd1 vccd1 _10978_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14229__B _14242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15505_ _15509_/A _15509_/B vssd1 vssd1 vccd1 vccd1 _15505_/Y sky130_fd_sc_hd__nand2_1
X_19273_ _20026_/CLK _19273_/D vssd1 vssd1 vccd1 vccd1 _19273_/Q sky130_fd_sc_hd__dfxtp_1
X_12717_ _12729_/C _12717_/B vssd1 vssd1 vccd1 vccd1 _12717_/X sky130_fd_sc_hd__xor2_4
XFILLER_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16485_ _16485_/A vssd1 vssd1 vccd1 vccd1 _19227_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18416__S _18418_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13697_ _18478_/Q _13526_/A _13695_/Y _13696_/X vssd1 vssd1 vccd1 vccd1 _18478_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17320__S _17326_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18224_ _19951_/Q _17656_/A _18230_/S vssd1 vssd1 vccd1 vccd1 _18225_/A sky130_fd_sc_hd__mux2_1
X_15436_ _15436_/A _15436_/B vssd1 vssd1 vccd1 vccd1 _15436_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12648_ _12648_/A _12695_/C vssd1 vssd1 vccd1 vccd1 _12648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14591__A1 _13579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18155_ _18155_/A vssd1 vssd1 vccd1 vccd1 _19920_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13394__A2 _18859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15367_ _15373_/A _15373_/B vssd1 vssd1 vccd1 vccd1 _15367_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14245__A _14245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12579_ _18475_/Q _12010_/X _12530_/A vssd1 vssd1 vccd1 vccd1 _12579_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17106_ _17643_/A vssd1 vssd1 vccd1 vccd1 _17106_/X sky130_fd_sc_hd__clkbuf_2
X_14318_ _14329_/D vssd1 vssd1 vccd1 vccd1 _14327_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18086_ _18086_/A vssd1 vssd1 vccd1 vccd1 _19897_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11944__A3 _11449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15298_ _15130_/X _15132_/X _15298_/S vssd1 vssd1 vccd1 vccd1 _15298_/X sky130_fd_sc_hd__mux2_1
X_17037_ _19466_/Q _17036_/X _17040_/S vssd1 vssd1 vccd1 vccd1 _17038_/A sky130_fd_sc_hd__mux2_1
X_14249_ _18651_/Q _14278_/D _14279_/C vssd1 vssd1 vccd1 vccd1 _14250_/B sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_17_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17293__A0 _17112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17990__S _17998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09790_ _11095_/A vssd1 vssd1 vccd1 vccd1 _09791_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _18992_/CLK _18988_/D vssd1 vssd1 vccd1 vccd1 _18988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _17939_/A vssd1 vssd1 vccd1 vccd1 _17948_/S sky130_fd_sc_hd__buf_4
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18387__A _18409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__A _10013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19609_ _19864_/CLK _19609_/D vssd1 vssd1 vccd1 vccd1 _19609_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13606__A0 _11860_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__A2 _11879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12866__C _12866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17230__S _17232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ _11659_/B _09306_/C vssd1 vssd1 vccd1 vccd1 _11941_/A sky130_fd_sc_hd__nor2_2
XFILLER_107_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14155__A _14245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14334__A1 _14336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11243__S1 _11022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09988_ _09988_/A vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__buf_2
XFILLER_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09471__A_N _09467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17405__S _17409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ _11950_/A vssd1 vssd1 vccd1 vccd1 _12859_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10754__S0 _10750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10901_ _20019_/Q _19857_/Q _19266_/Q _19036_/Q _10787_/A _10856_/A vssd1 vssd1 vccd1
+ vccd1 _10901_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15433__B _15436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _18712_/Q _17096_/B _11868_/X _11880_/X vssd1 vssd1 vccd1 vccd1 _11881_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11871__A2 _13164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10858__A _10858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13620_ _13709_/A _19008_/Q vssd1 vssd1 vccd1 vccd1 _13620_/Y sky130_fd_sc_hd__nand2_1
X_10832_ _10832_/A _10832_/B vssd1 vssd1 vccd1 vccd1 _10832_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13551_ _19000_/Q _13551_/B vssd1 vssd1 vccd1 vccd1 _13551_/X sky130_fd_sc_hd__or2_1
X_10763_ _10824_/A _10763_/B vssd1 vssd1 vccd1 vccd1 _10763_/X sky130_fd_sc_hd__or2_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12502_ _12502_/A _12523_/B vssd1 vssd1 vccd1 vccd1 _12502_/X sky130_fd_sc_hd__or2_1
X_16270_ _16270_/A vssd1 vssd1 vccd1 vccd1 _19147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13482_ _13481_/X _18454_/Q _13502_/S vssd1 vssd1 vccd1 vccd1 _13483_/A sky130_fd_sc_hd__mux2_1
X_10694_ _19143_/Q _19404_/Q _19303_/Q _19638_/Q _10521_/A _10638_/X vssd1 vssd1 vccd1
+ vccd1 _10695_/B sky130_fd_sc_hd__mux4_1
XFILLER_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15221_ _15236_/A _15221_/B _15221_/C vssd1 vssd1 vccd1 vccd1 _15221_/X sky130_fd_sc_hd__and3_1
XANTENNA__14573__A1 hold7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11689__A _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13376__A2 _12889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ _15355_/A _12433_/B vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__nor2_1
XFILLER_154_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ _14922_/S _15066_/X _14984_/A vssd1 vssd1 vccd1 vccd1 _15152_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ _12364_/A _12364_/B vssd1 vssd1 vccd1 vccd1 _12364_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_5_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14103_ _14105_/B _14105_/C _14102_/X vssd1 vssd1 vccd1 vccd1 _14103_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_153_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11315_ _19524_/Q vssd1 vssd1 vccd1 vccd1 _11414_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13128__A2 _13120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19960_ _19960_/CLK _19960_/D vssd1 vssd1 vccd1 vccd1 _19960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15083_ _15082_/A _15078_/B _15081_/X _15082_/Y vssd1 vssd1 vccd1 vccd1 _15083_/X
+ sky130_fd_sc_hd__o211a_1
X_12295_ _15936_/B vssd1 vssd1 vccd1 vccd1 _12295_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14034_ _18587_/Q _14034_/B _14034_/C vssd1 vssd1 vccd1 vccd1 _14036_/B sky130_fd_sc_hd__and3_1
X_18911_ _18911_/CLK _18911_/D vssd1 vssd1 vccd1 vccd1 _18911_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_141_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11246_ _09702_/A _11234_/X _11245_/X _09842_/A _18838_/Q vssd1 vssd1 vccd1 vccd1
+ _12828_/B sky130_fd_sc_hd__a32o_2
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19891_ _19896_/CLK _19891_/D vssd1 vssd1 vccd1 vccd1 _19891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10898__B1 _09774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18842_ _19324_/CLK _18842_/D vssd1 vssd1 vccd1 vccd1 _18842_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12313__A _12313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ _11309_/A vssd1 vssd1 vccd1 vccd1 _11225_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10128_ _10542_/A vssd1 vssd1 vccd1 vccd1 _10185_/A sky130_fd_sc_hd__buf_2
XFILLER_110_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15985_ _17738_/B vssd1 vssd1 vccd1 vccd1 _17426_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18773_ _18773_/CLK _18773_/D vssd1 vssd1 vccd1 vccd1 _18773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17315__S _17315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13843__S _13852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17724_ _17723_/X _19746_/Q _17730_/S vssd1 vssd1 vccd1 vccd1 _17725_/A sky130_fd_sc_hd__mux2_1
X_10059_ _19248_/Q _19743_/Q _10059_/S vssd1 vssd1 vccd1 vccd1 _10059_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15624__A _15624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14936_ _15436_/B _12298_/A _14937_/S vssd1 vssd1 vccd1 vccd1 _14936_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18000__A _18011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14867_ _14862_/X _14864_/X _14916_/S vssd1 vssd1 vccd1 vccd1 _14867_/X sky130_fd_sc_hd__mux2_1
X_17655_ _17655_/A vssd1 vssd1 vccd1 vccd1 _19724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13818_ _13818_/A vssd1 vssd1 vccd1 vccd1 _18504_/D sky130_fd_sc_hd__clkbuf_1
X_16606_ _16606_/A vssd1 vssd1 vccd1 vccd1 _19281_/D sky130_fd_sc_hd__clkbuf_1
X_17586_ _17632_/S vssd1 vssd1 vccd1 vccd1 _17595_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14798_ _14798_/A vssd1 vssd1 vccd1 vccd1 _18831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16537_ _19251_/Q _13845_/X _16541_/S vssd1 vssd1 vccd1 vccd1 _16538_/A sky130_fd_sc_hd__mux2_1
X_19325_ _19951_/CLK _19325_/D vssd1 vssd1 vccd1 vccd1 _19325_/Q sky130_fd_sc_hd__dfxtp_1
X_13749_ _14560_/A _19025_/Q _09341_/X _13748_/X vssd1 vssd1 vccd1 vccd1 _13750_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_32_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17050__S _17056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16468_ _19221_/Q _13851_/X _16468_/S vssd1 vssd1 vccd1 vccd1 _16469_/A sky130_fd_sc_hd__mux2_1
X_19256_ _19946_/CLK _19256_/D vssd1 vssd1 vccd1 vccd1 _19256_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17985__S _17987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18207_ _18207_/A vssd1 vssd1 vccd1 vccd1 _19944_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14564__A1 _14562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15419_ _15419_/A vssd1 vssd1 vccd1 vccd1 _15419_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19187_ _19972_/CLK _19187_/D vssd1 vssd1 vccd1 vccd1 _19187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16399_ _17735_/A vssd1 vssd1 vccd1 vccd1 _16399_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12575__B1 _18539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18138_ _18206_/S vssd1 vssd1 vccd1 vccd1 _18147_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09991__A1 _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18069_ _18069_/A vssd1 vssd1 vccd1 vccd1 _19892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09911_ _09911_/A vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20031_ _20031_/CLK _20031_/D vssd1 vssd1 vccd1 vccd1 _20031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09842_ _09842_/A vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__buf_4
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11550__A1 _09568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09773_/A vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__buf_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_14_0_clock clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10397__B _12853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12893__A _19488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09207_ _09190_/X _09206_/Y _09188_/A vssd1 vssd1 vccd1 vccd1 _14804_/A sky130_fd_sc_hd__o21ai_1
XFILLER_22_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11369__A1 _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14316__C _14317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11100_ _09755_/A _11099_/X _09773_/A vssd1 vssd1 vccd1 vccd1 _11100_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_192_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12080_ _12208_/A _12080_/B vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11031_ _19200_/Q _19791_/Q _19953_/Q _19168_/Q _10962_/X _11022_/X vssd1 vssd1 vccd1
+ vccd1 _11032_/B sky130_fd_sc_hd__mux4_1
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11541__A1 _09690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11972__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15770_ _09466_/A _15765_/X _15768_/X _15769_/X vssd1 vssd1 vccd1 vccd1 _18953_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _12982_/A vssd1 vssd1 vccd1 vccd1 _13511_/A sky130_fd_sc_hd__buf_2
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A io_dbus_rdata[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14721_ _18811_/Q _13677_/X _14727_/S vssd1 vssd1 vccd1 vccd1 _14722_/A sky130_fd_sc_hd__mux2_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _09499_/B _09248_/X _09265_/D _11931_/X _11932_/X vssd1 vssd1 vccd1 vccd1
+ _11945_/A sky130_fd_sc_hd__o2111ai_4
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17440_ _17115_/X _19628_/Q _17448_/S vssd1 vssd1 vccd1 vccd1 _17441_/A sky130_fd_sc_hd__mux2_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14652_ _14652_/A vssd1 vssd1 vccd1 vccd1 _14667_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _15789_/A vssd1 vssd1 vccd1 vccd1 _11865_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _13603_/A _18877_/Q _13603_/C vssd1 vssd1 vccd1 vccd1 _13614_/B sky130_fd_sc_hd__or3_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _09882_/A _10802_/X _10813_/X _09912_/A _10814_/Y vssd1 vssd1 vccd1 vccd1
+ _12841_/A sky130_fd_sc_hd__o32a_4
XFILLER_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17371_ _17371_/A vssd1 vssd1 vccd1 vccd1 _19597_/D sky130_fd_sc_hd__clkbuf_1
X_14583_ _14583_/A vssd1 vssd1 vccd1 vccd1 _18763_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14794__B2 _11956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11795_ _18585_/Q _11851_/A _11794_/X _18617_/Q vssd1 vssd1 vccd1 vccd1 _11796_/C
+ sky130_fd_sc_hd__a22o_1
X_19110_ _19637_/CLK _19110_/D vssd1 vssd1 vccd1 vccd1 _19110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16322_ _16322_/A vssd1 vssd1 vccd1 vccd1 _19166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13534_ _18869_/Q _13535_/B vssd1 vssd1 vccd1 vccd1 _13554_/C sky130_fd_sc_hd__or2_1
XFILLER_158_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10746_ _10739_/Y _10741_/Y _10743_/Y _10745_/Y _09820_/A vssd1 vssd1 vccd1 vccd1
+ _10746_/X sky130_fd_sc_hd__o221a_2
XFILLER_14_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19041_ _20026_/CLK _19041_/D vssd1 vssd1 vccd1 vccd1 _19041_/Q sky130_fd_sc_hd__dfxtp_1
X_16253_ _16253_/A vssd1 vssd1 vccd1 vccd1 _19139_/D sky130_fd_sc_hd__clkbuf_1
X_13465_ _13465_/A vssd1 vssd1 vccd1 vccd1 _18453_/D sky130_fd_sc_hd__clkbuf_1
X_10677_ _10670_/X _10672_/X _10674_/X _10676_/X _09875_/A vssd1 vssd1 vccd1 vccd1
+ _10677_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11212__A _11212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15204_ _15200_/X _15203_/X _15247_/A vssd1 vssd1 vccd1 vccd1 _15204_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12416_ _18531_/Q _12416_/B _12416_/C _12416_/D vssd1 vssd1 vccd1 vccd1 _12446_/B
+ sky130_fd_sc_hd__and4_1
X_16184_ _13202_/X _19110_/Q _16184_/S vssd1 vssd1 vccd1 vccd1 _16185_/A sky130_fd_sc_hd__mux2_1
X_13396_ _18480_/Q _12943_/X _12944_/X _18704_/Q _13395_/X vssd1 vssd1 vccd1 vccd1
+ _13396_/X sky130_fd_sc_hd__a221o_1
XANTENNA__12027__B _12234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15135_ _15131_/X _15134_/X _15171_/S vssd1 vssd1 vccd1 vccd1 _15135_/X sky130_fd_sc_hd__mux2_1
X_12347_ _12347_/A vssd1 vssd1 vccd1 vccd1 _12347_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output80_A _12498_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19943_ _20007_/CLK _19943_/D vssd1 vssd1 vccd1 vccd1 _19943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15066_ _14980_/X _15065_/X _15202_/S vssd1 vssd1 vccd1 vccd1 _15066_/X sky130_fd_sc_hd__mux2_1
X_12278_ _12278_/A _12340_/C vssd1 vssd1 vccd1 vccd1 _12279_/D sky130_fd_sc_hd__or2_1
XANTENNA__17248__A0 _17151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14017_ _14046_/A _14017_/B vssd1 vssd1 vccd1 vccd1 _14017_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17834__A _17880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _19384_/Q vssd1 vssd1 vccd1 vccd1 _11442_/S sky130_fd_sc_hd__buf_2
XFILLER_136_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19874_ _20006_/CLK _19874_/D vssd1 vssd1 vccd1 vccd1 _19874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18825_ _18960_/CLK _18825_/D vssd1 vssd1 vccd1 vccd1 _18825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18756_ _19063_/CLK _18756_/D vssd1 vssd1 vccd1 vccd1 _18756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15968_ _15982_/A _15968_/B vssd1 vssd1 vccd1 vccd1 _15968_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10718__S0 _10764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17707_ _17707_/A vssd1 vssd1 vccd1 vccd1 _17707_/X sky130_fd_sc_hd__clkbuf_2
X_14919_ _14905_/X _14917_/X _15082_/B vssd1 vssd1 vccd1 vccd1 _14919_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16884__S _16892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18687_ _18687_/CLK _18687_/D vssd1 vssd1 vccd1 vccd1 _18687_/Q sky130_fd_sc_hd__dfxtp_1
X_15899_ _15899_/A _15899_/B vssd1 vssd1 vccd1 vccd1 _15899_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17638_ _17634_/X _19719_/Q _17650_/S vssd1 vssd1 vccd1 vccd1 _17639_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13037__A1 _13551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17569_ _17106_/X _19689_/Q _17573_/S vssd1 vssd1 vccd1 vccd1 _17570_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19308_ _19965_/CLK _19308_/D vssd1 vssd1 vccd1 vccd1 _19308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19239_ _19993_/CLK _19239_/D vssd1 vssd1 vccd1 vccd1 _19239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11122__A _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11446__S1 _19385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11220__B1 _11058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10961__A _11295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17239__A0 _17138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09811__S1 _09895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10957__S0 _10892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20014_ _20016_/CLK _20014_/D vssd1 vssd1 vccd1 vccd1 _20014_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input4_A io_dbus_rdata[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _19382_/Q _19717_/Q _09903_/A vssd1 vssd1 vccd1 vccd1 _09826_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09756_ _11032_/A vssd1 vssd1 vccd1 vccd1 _10947_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _09687_/A vssd1 vssd1 vccd1 vccd1 _10192_/A sky130_fd_sc_hd__buf_2
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11826__A2 _12876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11382__S0 _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_139_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10600_ _11006_/A vssd1 vssd1 vccd1 vccd1 _10727_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11580_ _11581_/A _11582_/B _11580_/C vssd1 vssd1 vccd1 vccd1 _11580_/Y sky130_fd_sc_hd__nand3_1
XFILLER_11_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10531_ _10473_/X _10528_/X _10530_/X vssd1 vssd1 vccd1 vccd1 _10531_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_168_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13250_ _17691_/A vssd1 vssd1 vccd1 vccd1 _13250_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10462_ _10462_/A _10462_/B vssd1 vssd1 vccd1 vccd1 _10462_/X sky130_fd_sc_hd__or2_1
XANTENNA__13200__A1 _13005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ _18764_/Q _12200_/X _13595_/A vssd1 vssd1 vccd1 vccd1 _12201_/Y sky130_fd_sc_hd__o21ai_1
X_13181_ _13180_/X _18437_/Q _13203_/S vssd1 vssd1 vccd1 vccd1 _13182_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13751__A2 _13746_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16034__S _16042_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10393_ _19341_/Q _19612_/Q _19836_/Q _19580_/Q _10141_/X _10283_/A vssd1 vssd1 vccd1
+ vccd1 _10393_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12132_ _18459_/Q _12472_/A vssd1 vssd1 vccd1 vccd1 _12132_/X sky130_fd_sc_hd__or2_1
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16969__S _16975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12063_ _12065_/B _12060_/X _12062_/Y _12016_/X _16075_/A vssd1 vssd1 vccd1 vccd1
+ _12071_/B sky130_fd_sc_hd__a32o_1
X_16940_ _16326_/X _19429_/Q _16942_/S vssd1 vssd1 vccd1 vccd1 _16941_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11014_ _11295_/S vssd1 vssd1 vccd1 vccd1 _11017_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16871_ _16871_/A vssd1 vssd1 vccd1 vccd1 _19398_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10868__A3 _10867_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18610_ _18744_/CLK _18610_/D vssd1 vssd1 vccd1 vccd1 _18610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15822_ _15831_/A _15822_/B vssd1 vssd1 vccd1 vccd1 _15823_/A sky130_fd_sc_hd__and2_1
XFILLER_92_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19590_ _19856_/CLK _19590_/D vssd1 vssd1 vccd1 vccd1 _19590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15753_ _18947_/Q _15760_/B vssd1 vssd1 vccd1 vccd1 _15753_/X sky130_fd_sc_hd__or2_1
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18541_ _18928_/CLK _18541_/D vssd1 vssd1 vccd1 vccd1 _18541_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _12965_/A vssd1 vssd1 vccd1 vccd1 _18426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11916_ _14744_/B _12472_/A _12503_/A _12350_/A vssd1 vssd1 vccd1 vccd1 _13861_/C
+ sky130_fd_sc_hd__a31o_1
X_14704_ _14704_/A vssd1 vssd1 vccd1 vccd1 _18803_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10111__A _10411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15684_ _18919_/Q _12601_/A _15688_/S vssd1 vssd1 vccd1 vccd1 _15685_/A sky130_fd_sc_hd__mux2_1
X_18472_ _18547_/CLK _18472_/D vssd1 vssd1 vccd1 vccd1 _18472_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _19486_/Q vssd1 vssd1 vccd1 vccd1 _12957_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _17423_/A vssd1 vssd1 vccd1 vccd1 _19621_/D sky130_fd_sc_hd__clkbuf_1
X_14635_ _14652_/A vssd1 vssd1 vccd1 vccd1 _14649_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _11847_/A vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16209__S _16217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09869__S1 _09639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _17882_/B _17954_/B vssd1 vssd1 vccd1 vccd1 _17411_/A sky130_fd_sc_hd__nor2_2
X_14566_ _14566_/A vssd1 vssd1 vccd1 vccd1 _18758_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11778_ _12060_/A _11780_/B vssd1 vssd1 vccd1 vccd1 _11778_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16305_ _16304_/X _19161_/Q _16314_/S vssd1 vssd1 vccd1 vccd1 _16306_/A sky130_fd_sc_hd__mux2_1
X_13517_ _13517_/A vssd1 vssd1 vccd1 vccd1 _13517_/X sky130_fd_sc_hd__buf_2
XFILLER_174_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10729_ _10050_/A _10724_/X _10728_/X vssd1 vssd1 vccd1 vccd1 _10729_/Y sky130_fd_sc_hd__a21oi_1
X_17285_ _17097_/X _19559_/Q _17293_/S vssd1 vssd1 vccd1 vccd1 _17286_/A sky130_fd_sc_hd__mux2_1
X_14497_ _14514_/A _14501_/C vssd1 vssd1 vccd1 vccd1 _14497_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16236_ _13002_/X _19132_/Q _16236_/S vssd1 vssd1 vccd1 vccd1 _16237_/A sky130_fd_sc_hd__mux2_1
X_19024_ _19025_/CLK _19024_/D vssd1 vssd1 vccd1 vccd1 _19024_/Q sky130_fd_sc_hd__dfxtp_2
X_13448_ _13737_/A _13449_/B vssd1 vssd1 vccd1 vccd1 _13448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11202__B1 _11425_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13742__A2 _19024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16167_ _13042_/X _19102_/Q _16173_/S vssd1 vssd1 vccd1 vccd1 _16168_/A sky130_fd_sc_hd__mux2_1
X_13379_ _14095_/A _13120_/X _13194_/X _14518_/A vssd1 vssd1 vccd1 vccd1 _13379_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18130__A1 _13742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15118_ _15030_/X _15036_/X _15118_/S vssd1 vssd1 vccd1 vccd1 _15118_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16098_ _13098_/X _19072_/Q _16100_/S vssd1 vssd1 vccd1 vccd1 _16099_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16879__S _16881_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19926_ _19990_/CLK _19926_/D vssd1 vssd1 vccd1 vccd1 _19926_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17564__A _17632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15049_ _15006_/X _15428_/A _15047_/X _15048_/X _11971_/Y vssd1 vssd1 vccd1 vccd1
+ _15049_/X sky130_fd_sc_hd__a32o_1
XFILLER_123_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19857_ _20018_/CLK _19857_/D vssd1 vssd1 vccd1 vccd1 _19857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09610_ _09610_/A vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18808_ _19899_/CLK _18808_/D vssd1 vssd1 vccd1 vccd1 _18808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12501__A _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19788_ _19950_/CLK _19788_/D vssd1 vssd1 vccd1 vccd1 _19788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09541_ _19485_/Q vssd1 vssd1 vccd1 vccd1 _09542_/A sky130_fd_sc_hd__inv_2
X_18739_ _19909_/CLK _18739_/D vssd1 vssd1 vccd1 vccd1 _18739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10021__A _10521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09472_ _12055_/A _12055_/B _12055_/C _09471_/X vssd1 vssd1 vccd1 vccd1 _15633_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_140_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11116__S0 _11186_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10167__S _10279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17739__A _17795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16643__A _16689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19981_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09937__B2 _18861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16789__S _16797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_65_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13497__A1 _12875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09808_ _09750_/X _09781_/X _09783_/X _09800_/X _09807_/X vssd1 vssd1 vccd1 vccd1
+ _09808_/X sky130_fd_sc_hd__a221o_1
XFILLER_101_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09739_ _10624_/A vssd1 vssd1 vccd1 vccd1 _10793_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14997__A1 _15139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _18785_/Q _12750_/B _12750_/C vssd1 vssd1 vccd1 vccd1 _12774_/B sky130_fd_sc_hd__and3_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11701_/A vssd1 vssd1 vccd1 vccd1 _14555_/B sky130_fd_sc_hd__buf_2
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09720__A _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12674_/A _12673_/X _12677_/Y _12680_/Y vssd1 vssd1 vccd1 vccd1 _12681_/X
+ sky130_fd_sc_hd__o22a_4
XANTENNA__16029__S _16031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14420_ _14452_/A _14420_/B _14420_/C vssd1 vssd1 vccd1 vccd1 _18701_/D sky130_fd_sc_hd__nor3_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11634_/A _11522_/A _10352_/A _11588_/A vssd1 vssd1 vccd1 vccd1 _11633_/C
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13421__A1 _13223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__B _12848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14351_ _14356_/A _14351_/B _14355_/C vssd1 vssd1 vccd1 vccd1 _18681_/D sky130_fd_sc_hd__nor3_1
X_11563_ _09837_/X _11556_/X _11558_/X _11562_/X _09807_/X vssd1 vssd1 vccd1 vccd1
+ _11563_/X sky130_fd_sc_hd__a311o_1
XFILLER_7_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18244__S _18252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13302_ _17700_/A vssd1 vssd1 vccd1 vccd1 _13302_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11983__A1 _11982_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17070_ _17070_/A vssd1 vssd1 vccd1 vccd1 _19476_/D sky130_fd_sc_hd__clkbuf_1
X_10514_ _15956_/B vssd1 vssd1 vccd1 vccd1 _10539_/A sky130_fd_sc_hd__inv_2
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14282_ _18660_/Q _14287_/D _14792_/A vssd1 vssd1 vccd1 vccd1 _14283_/B sky130_fd_sc_hd__o21ai_1
X_11494_ _19141_/Q _19402_/Q _19301_/Q _19636_/Q _10906_/S _10625_/A vssd1 vssd1 vccd1
+ vccd1 _11495_/B sky130_fd_sc_hd__mux4_1
XFILLER_6_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16021_ _16021_/A vssd1 vssd1 vccd1 vccd1 _19040_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13185__B1 _12897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ _13233_/A _13368_/A vssd1 vssd1 vccd1 vccd1 _13319_/A sky130_fd_sc_hd__or2_1
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _11589_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10805__S _10859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12932__B1 _12890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164_ _19894_/Q _13164_/B vssd1 vssd1 vccd1 vccd1 _13164_/X sky130_fd_sc_hd__and2_1
X_10376_ _10376_/A vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__buf_2
XANTENNA__16699__S _16703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output166_A _12821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12115_ _11903_/A _12828_/B _12175_/A _09261_/B vssd1 vssd1 vccd1 vccd1 _15160_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_124_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14223__D _16474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17972_ _19854_/Q _17017_/X _17976_/S vssd1 vssd1 vccd1 vccd1 _17973_/A sky130_fd_sc_hd__mux2_1
X_13095_ input31/X _13091_/X _13094_/X vssd1 vssd1 vccd1 vccd1 _13095_/X sky130_fd_sc_hd__a21o_1
XFILLER_78_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19711_ _20035_/CLK _19711_/D vssd1 vssd1 vccd1 vccd1 _19711_/Q sky130_fd_sc_hd__dfxtp_1
X_16923_ _16297_/X _19421_/Q _16931_/S vssd1 vssd1 vccd1 vccd1 _16924_/A sky130_fd_sc_hd__mux2_1
X_12046_ _12046_/A _12046_/B vssd1 vssd1 vccd1 vccd1 _12046_/Y sky130_fd_sc_hd__xnor2_4
X_19642_ _19996_/CLK _19642_/D vssd1 vssd1 vccd1 vccd1 _19642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16854_ _16854_/A vssd1 vssd1 vccd1 vccd1 _19390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ input60/X vssd1 vssd1 vccd1 vccd1 _15805_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19573_ _19829_/CLK _19573_/D vssd1 vssd1 vccd1 vccd1 _19573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13997_ _14094_/A vssd1 vssd1 vccd1 vccd1 _14044_/A sky130_fd_sc_hd__clkbuf_4
X_16785_ _16785_/A vssd1 vssd1 vccd1 vccd1 _19360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18524_ _18526_/CLK _18524_/D vssd1 vssd1 vccd1 vccd1 _18524_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15736_ _16691_/A _15745_/B vssd1 vssd1 vccd1 vccd1 _15736_/X sky130_fd_sc_hd__or2_1
X_12948_ _19883_/Q _13373_/B vssd1 vssd1 vccd1 vccd1 _12948_/X sky130_fd_sc_hd__and2_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18455_ _19856_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _12879_/A vssd1 vssd1 vccd1 vccd1 _12879_/X sky130_fd_sc_hd__clkbuf_4
X_15667_ _15667_/A vssd1 vssd1 vccd1 vccd1 _18911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ _17406_/A vssd1 vssd1 vccd1 vccd1 _19613_/D sky130_fd_sc_hd__clkbuf_1
X_14618_ _14652_/A vssd1 vssd1 vccd1 vccd1 _14632_/S sky130_fd_sc_hd__clkbuf_2
X_18386_ _18386_/A vssd1 vssd1 vccd1 vccd1 _20023_/D sky130_fd_sc_hd__clkbuf_1
X_15598_ _18881_/Q _18913_/Q _15600_/S vssd1 vssd1 vccd1 vccd1 _15599_/A sky130_fd_sc_hd__mux2_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17337_ _17176_/X _19583_/Q _17337_/S vssd1 vssd1 vccd1 vccd1 _17338_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11423__B1 _11003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14549_ _18755_/Q _14547_/X _14548_/X _14540_/X vssd1 vssd1 vccd1 vccd1 _18755_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18154__S _18158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__S1 _10320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11974__A1 _11650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17268_ _17179_/X _19552_/Q _17276_/S vssd1 vssd1 vccd1 vccd1 _17269_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19007_ _19025_/CLK _19007_/D vssd1 vssd1 vccd1 vccd1 _19007_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_161_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16219_ _13481_/X _19126_/Q _16221_/S vssd1 vssd1 vccd1 vccd1 _16220_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17199_ _17198_/X _19521_/Q _17199_/S vssd1 vssd1 vccd1 vccd1 _17200_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16114__A0 _13219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15807__A _15807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19909_ _19909_/CLK _19909_/D vssd1 vssd1 vccd1 vccd1 _19909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18329__S _18335_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09524_ _12536_/A _14819_/B _11937_/B vssd1 vssd1 vccd1 vccd1 _09525_/D sky130_fd_sc_hd__and3_1
XFILLER_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_141_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18655_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _18968_/Q vssd1 vssd1 vccd1 vccd1 _12003_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09386_ _18954_/Q _18953_/Q vssd1 vssd1 vccd1 vccd1 _11697_/B sky130_fd_sc_hd__or2_1
XANTENNA__13997__A _14094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_156_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19888_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11965__A1 _11945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10230_ _19939_/Q _19553_/Q _20003_/Q _19122_/Q _10166_/S _10223_/X vssd1 vssd1 vccd1
+ vccd1 _10231_/B sky130_fd_sc_hd__mux4_1
XFILLER_134_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ _10144_/X _10155_/X _10157_/X _10160_/X _09807_/A vssd1 vssd1 vccd1 vccd1
+ _10161_/X sky130_fd_sc_hd__a221o_1
XFILLER_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14667__A0 _18788_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09769__S0 _09733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10092_ _19679_/Q _19445_/Q _18510_/Q _19775_/Q _09939_/A _10278_/A vssd1 vssd1 vccd1
+ vccd1 _10093_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13237__A _17046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13920_ _18607_/Q _18609_/Q _18608_/Q _14089_/A vssd1 vssd1 vccd1 vccd1 _14099_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13851_ _17087_/A vssd1 vssd1 vccd1 vccd1 _13851_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18239__S _18241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12802_ _12788_/A _12789_/A _12788_/B _12784_/A _15542_/B vssd1 vssd1 vccd1 vccd1
+ _12812_/A sky130_fd_sc_hd__a32o_2
X_16570_ _16570_/A vssd1 vssd1 vccd1 vccd1 _19265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13782_ _18493_/Q _13781_/X _13788_/S vssd1 vssd1 vccd1 vccd1 _13783_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10994_ _11140_/A vssd1 vssd1 vccd1 vccd1 _11137_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_109_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _20034_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10456__A1 _09566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _12753_/A _12862_/B vssd1 vssd1 vccd1 vccd1 _12733_/Y sky130_fd_sc_hd__nor2_1
X_15521_ _15159_/X _15516_/Y _15520_/Y vssd1 vssd1 vccd1 vccd1 _15522_/C sky130_fd_sc_hd__a21oi_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16982__S _16986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10596__A _10596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18240_ _18240_/A vssd1 vssd1 vccd1 vccd1 _19958_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15452_ _15365_/X _15246_/X _15451_/X _15400_/X vssd1 vssd1 vccd1 vccd1 _15452_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12664_/A vssd1 vssd1 vccd1 vccd1 _15487_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _18696_/Q _14399_/C _14402_/Y vssd1 vssd1 vccd1 vccd1 _18696_/D sky130_fd_sc_hd__o21a_1
XFILLER_169_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11615_ _11616_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11615_/Y sky130_fd_sc_hd__nand2_1
X_18171_ _18193_/A vssd1 vssd1 vccd1 vccd1 _18180_/S sky130_fd_sc_hd__buf_2
X_15383_ _15366_/X _15380_/Y _15382_/X _15353_/X vssd1 vssd1 vccd1 vccd1 _15387_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_169_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12595_ _12595_/A vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__clkinv_2
X_14334_ _14336_/B _14338_/D _14333_/Y vssd1 vssd1 vccd1 vccd1 _18675_/D sky130_fd_sc_hd__o21a_1
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17122_ _17659_/A vssd1 vssd1 vccd1 vccd1 _17122_/X sky130_fd_sc_hd__clkbuf_2
X_11546_ _19944_/Q _19558_/Q _20008_/Q _19127_/Q _11532_/S _09614_/X vssd1 vssd1 vccd1
+ vccd1 _11547_/B sky130_fd_sc_hd__mux4_1
XFILLER_7_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17098__B _17098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _19471_/Q _17052_/X _17056_/S vssd1 vssd1 vccd1 vccd1 _17054_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14265_ _14265_/A _14275_/D vssd1 vssd1 vccd1 vccd1 _14265_/Y sky130_fd_sc_hd__nor2_1
X_11477_ _11477_/A _11477_/B vssd1 vssd1 vccd1 vccd1 _11477_/X sky130_fd_sc_hd__or2_1
XFILLER_125_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12316__A _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18097__A0 _18853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16004_ _16004_/A vssd1 vssd1 vccd1 vccd1 _19032_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12905__B1 _19487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13216_ _13207_/Y _13208_/X _13215_/X _13350_/S _13297_/A vssd1 vssd1 vccd1 vccd1
+ _13217_/B sky130_fd_sc_hd__a221o_1
XFILLER_171_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10428_ _19148_/Q _19409_/Q _19308_/Q _19643_/Q _10152_/X _10153_/X vssd1 vssd1 vccd1
+ vccd1 _10429_/B sky130_fd_sc_hd__mux4_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14196_ _18637_/Q _14197_/C _18638_/Q vssd1 vssd1 vccd1 vccd1 _14198_/B sky130_fd_sc_hd__a21oi_1
XFILLER_152_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13846__S _13852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17318__S _17326_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ input3/X _13091_/X _13094_/X vssd1 vssd1 vccd1 vccd1 _13147_/X sky130_fd_sc_hd__a21o_1
X_10359_ _19149_/Q _19410_/Q _19309_/Q _19644_/Q _10356_/S _10261_/A vssd1 vssd1 vccd1
+ vccd1 _10360_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09625__A _10674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _18011_/A vssd1 vssd1 vccd1 vccd1 _18024_/S sky130_fd_sc_hd__buf_6
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _18622_/Q vssd1 vssd1 vccd1 vccd1 _14153_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _16380_/X _19414_/Q _16914_/S vssd1 vssd1 vccd1 vccd1 _16907_/A sky130_fd_sc_hd__mux2_1
X_12029_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12208_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09344__B _09442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__A _18520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17886_ _17886_/A vssd1 vssd1 vccd1 vccd1 _19815_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19625_ _19979_/CLK _19625_/D vssd1 vssd1 vccd1 vccd1 _19625_/Q sky130_fd_sc_hd__dfxtp_1
X_16837_ _17201_/A _16837_/B vssd1 vssd1 vccd1 vccd1 _16838_/A sky130_fd_sc_hd__and2_1
XANTENNA__11892__B1 _11843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17053__S _17056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19556_ _20006_/CLK _19556_/D vssd1 vssd1 vccd1 vccd1 _19556_/Q sky130_fd_sc_hd__dfxtp_1
X_16768_ _16768_/A vssd1 vssd1 vccd1 vccd1 _19352_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13633__A1 _13632_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18507_ _19836_/CLK _18507_/D vssd1 vssd1 vccd1 vccd1 _18507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_13_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09932__S0 _09659_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15719_ _15719_/A vssd1 vssd1 vccd1 vccd1 _15773_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16892__S _16892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19487_ _19487_/CLK _19487_/D vssd1 vssd1 vccd1 vccd1 _19487_/Q sky130_fd_sc_hd__dfxtp_2
X_16699_ _19322_/Q _13765_/X _16703_/S vssd1 vssd1 vccd1 vccd1 _16700_/A sky130_fd_sc_hd__mux2_1
X_09240_ _09284_/A _09247_/B _09247_/C vssd1 vssd1 vccd1 vccd1 _09290_/B sky130_fd_sc_hd__or3_1
XFILLER_62_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18438_ _19636_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_73_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19350_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13397__B1 _12879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09171_ _18966_/Q vssd1 vssd1 vccd1 vccd1 _09285_/C sky130_fd_sc_hd__clkbuf_1
X_18369_ _18369_/A vssd1 vssd1 vccd1 vccd1 _20015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13610__A _14552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_88_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 _19997_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16921__A _16977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14897__A0 _15100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18088__A0 _18850_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17228__S _17232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10383__B1 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19758_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10349__A2_N _09843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10180__S _10180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09254__B _18989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10230__S0 _10166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19824_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09507_ _15139_/A _15899_/B vssd1 vssd1 vccd1 vccd1 _09508_/C sky130_fd_sc_hd__nor2_1
XANTENNA__09923__S0 _09659_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17898__S _17904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10533__S1 _10011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _12003_/C _09309_/A _14761_/C vssd1 vssd1 vccd1 vccd1 _15393_/A sky130_fd_sc_hd__a21oi_4
XFILLER_12_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _18960_/Q _18959_/Q _18958_/Q _18957_/Q vssd1 vssd1 vccd1 vccd1 _09378_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_166_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11400_ _18425_/Q _19454_/Q _19491_/Q _19065_/Q _11442_/S _11019_/A vssd1 vssd1 vccd1
+ vccd1 _11401_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13520__A _13520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12380_ _09522_/A _12428_/A _12379_/Y vssd1 vssd1 vccd1 vccd1 _15338_/A sky130_fd_sc_hd__a21o_2
XFILLER_166_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11331_ _18426_/Q _19455_/Q _19492_/Q _19066_/Q _11328_/X _11322_/X vssd1 vssd1 vccd1
+ vccd1 _11332_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09429__B _12918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14050_ _14094_/A vssd1 vssd1 vccd1 vccd1 _14088_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11262_ _19133_/Q _19394_/Q _19293_/Q _19628_/Q _10977_/S _11045_/X vssd1 vssd1 vccd1
+ vccd1 _11262_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13001_ _17007_/A vssd1 vssd1 vccd1 vccd1 _17649_/A sky130_fd_sc_hd__clkbuf_2
X_10213_ _10695_/A vssd1 vssd1 vccd1 vccd1 _10520_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16042__S _16042_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11193_ _11242_/A _11190_/X _11192_/X vssd1 vssd1 vccd1 vccd1 _11193_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input42_A io_ibus_inst[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _10392_/A _10144_/B vssd1 vssd1 vccd1 vccd1 _10144_/X sky130_fd_sc_hd__or2_1
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11186__S _11186_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12115__B2 _09261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13312__B1 _12984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17662__A _17662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17740_ _17808_/S vssd1 vssd1 vccd1 vccd1 _17749_/S sky130_fd_sc_hd__clkbuf_4
X_10075_ _10270_/A _10074_/X _09690_/A vssd1 vssd1 vccd1 vccd1 _10075_/Y sky130_fd_sc_hd__o21ai_1
X_14952_ _12807_/B _12870_/B _14955_/S vssd1 vssd1 vccd1 vccd1 _14952_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13903_ _12674_/A _13900_/X _12677_/Y _12680_/Y _13897_/X vssd1 vssd1 vccd1 vccd1
+ _18543_/D sky130_fd_sc_hd__o221a_1
XFILLER_130_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17671_ _17671_/A vssd1 vssd1 vccd1 vccd1 _19729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11874__B1 _13335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14883_ _14883_/A vssd1 vssd1 vccd1 vccd1 _15321_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_output129_A _12862_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19410_ _19644_/CLK _19410_/D vssd1 vssd1 vccd1 vccd1 _19410_/Q sky130_fd_sc_hd__dfxtp_1
X_16622_ _16297_/X _19288_/Q _16630_/S vssd1 vssd1 vccd1 vccd1 _16623_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13834_ _13834_/A vssd1 vssd1 vccd1 vccd1 _18509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19341_ _19836_/CLK _19341_/D vssd1 vssd1 vccd1 vccd1 _19341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16553_ _16553_/A vssd1 vssd1 vccd1 vccd1 _19257_/D sky130_fd_sc_hd__clkbuf_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ _17001_/A vssd1 vssd1 vccd1 vccd1 _13765_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11860__D _11860_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10977_ _19360_/Q _19695_/Q _10977_/S vssd1 vssd1 vccd1 vccd1 _10978_/B sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_187_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ _18859_/Q _15457_/X _15503_/X vssd1 vssd1 vccd1 vccd1 _18859_/D sky130_fd_sc_hd__o21a_1
X_19272_ _20025_/CLK _19272_/D vssd1 vssd1 vccd1 vccd1 _19272_/Q sky130_fd_sc_hd__dfxtp_1
X_12716_ _12689_/A _15498_/B _12729_/B _12692_/B vssd1 vssd1 vccd1 vccd1 _12717_/B
+ sky130_fd_sc_hd__a22o_1
X_16484_ _19227_/Q _13768_/X _16486_/S vssd1 vssd1 vccd1 vccd1 _16485_/A sky130_fd_sc_hd__mux2_1
X_13696_ _13650_/X _11898_/X _13514_/S vssd1 vssd1 vccd1 vccd1 _13696_/X sky130_fd_sc_hd__a21bo_1
XFILLER_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18223_ _18223_/A vssd1 vssd1 vccd1 vccd1 _19950_/D sky130_fd_sc_hd__clkbuf_1
X_15435_ _15099_/X _15432_/Y _15434_/X _15105_/X vssd1 vssd1 vccd1 vccd1 _15438_/B
+ sky130_fd_sc_hd__a211o_1
X_12647_ _18542_/Q _12647_/B vssd1 vssd1 vccd1 vccd1 _12695_/C sky130_fd_sc_hd__and2_1
XANTENNA__16217__S _16217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18154_ _17659_/X _19920_/Q _18158_/S vssd1 vssd1 vccd1 vccd1 _18155_/A sky130_fd_sc_hd__mux2_1
X_15366_ _15366_/A vssd1 vssd1 vccd1 vccd1 _15366_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11869__B _11869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12578_ _12574_/X _12577_/Y _12770_/S vssd1 vssd1 vccd1 vccd1 _12578_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ _17105_/A vssd1 vssd1 vccd1 vccd1 _19491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11529_ _11529_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11580_/C sky130_fd_sc_hd__nand2_1
X_14317_ _18671_/Q _18670_/Q _18669_/Q _14317_/D vssd1 vssd1 vccd1 vccd1 _14329_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15297_ _18844_/Q _15278_/X _15296_/X vssd1 vssd1 vccd1 vccd1 _18844_/D sky130_fd_sc_hd__o21a_1
X_18085_ _18084_/X _19897_/Q _18095_/S vssd1 vssd1 vccd1 vccd1 _18086_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17036_ _17036_/A vssd1 vssd1 vccd1 vccd1 _17036_/X sky130_fd_sc_hd__clkbuf_2
X_14248_ _14278_/D _14279_/C _14247_/Y vssd1 vssd1 vccd1 vccd1 _18650_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14179_ _18631_/Q _14180_/C _18632_/Q vssd1 vssd1 vccd1 vccd1 _14181_/B sky130_fd_sc_hd__a21oi_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _18992_/CLK _18987_/D vssd1 vssd1 vccd1 vccd1 _18987_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _17938_/A vssd1 vssd1 vccd1 vccd1 _19839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17869_ _17869_/A vssd1 vssd1 vccd1 vccd1 _19808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19608_ _19864_/CLK _19608_/D vssd1 vssd1 vccd1 vccd1 _19608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19539_ _19989_/CLK _19539_/D vssd1 vssd1 vccd1 vccd1 _19539_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09905__S0 _09903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ _09230_/A _09274_/A vssd1 vssd1 vccd1 vccd1 _09306_/C sky130_fd_sc_hd__and2b_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16127__S _16133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13340__A _13340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_10_0_clock clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_147_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18342__S _18346_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09987_ _09987_/A vssd1 vssd1 vccd1 vccd1 _09988_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16797__S _16797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11856__B1 _13189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10754__S1 _10626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ _10900_/A _10900_/B vssd1 vssd1 vccd1 vccd1 _10900_/X sky130_fd_sc_hd__or2_1
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11880_ _11773_/A _11879_/X _11812_/B vssd1 vssd1 vccd1 vccd1 _11880_/X sky130_fd_sc_hd__a21bo_1
XFILLER_83_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ _19924_/Q _19538_/Q _19988_/Q _19107_/Q _11467_/S _10820_/A vssd1 vssd1 vccd1
+ vccd1 _10832_/B sky130_fd_sc_hd__mux4_1
XFILLER_26_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ _13550_/A vssd1 vssd1 vccd1 vccd1 _18459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10762_ _19667_/Q _19433_/Q _18498_/Q _19763_/Q _10872_/S _10664_/A vssd1 vssd1 vccd1
+ vccd1 _10763_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12281__B1 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12501_ _12501_/A _12501_/B _12501_/C vssd1 vssd1 vccd1 vccd1 _12523_/B sky130_fd_sc_hd__and3_1
XFILLER_158_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13481_ _17732_/A vssd1 vssd1 vccd1 vccd1 _13481_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10693_ _10643_/A _10688_/X _10690_/Y _10692_/Y vssd1 vssd1 vccd1 vccd1 _10693_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12033__A0 _14749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15220_ _15218_/X _15210_/Y _15219_/Y vssd1 vssd1 vccd1 vccd1 _15221_/C sky130_fd_sc_hd__a21oi_1
X_12432_ _11949_/X _12432_/B _12432_/C vssd1 vssd1 vccd1 vccd1 _14966_/A sky130_fd_sc_hd__nand3b_4
XFILLER_173_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15770__A1 _09466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10044__C1 _09807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15151_ _15151_/A vssd1 vssd1 vccd1 vccd1 _15151_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12363_ _12334_/A _12334_/B _12329_/A vssd1 vssd1 vccd1 vccd1 _12364_/B sky130_fd_sc_hd__a21oi_2
XFILLER_153_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18252__S _18252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14102_ _14102_/A vssd1 vssd1 vccd1 vccd1 _14102_/X sky130_fd_sc_hd__buf_2
XFILLER_153_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11314_ _18836_/Q _09841_/A _09881_/A _11313_/X vssd1 vssd1 vccd1 vccd1 _12826_/B
+ sky130_fd_sc_hd__o2bb2a_4
X_15082_ _15082_/A _15082_/B vssd1 vssd1 vccd1 vccd1 _15082_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12294_ _12294_/A _15291_/A vssd1 vssd1 vccd1 vccd1 _12297_/A sky130_fd_sc_hd__xor2_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14033_ _14034_/B _14034_/C _14032_/Y vssd1 vssd1 vccd1 vccd1 _18586_/D sky130_fd_sc_hd__o21a_1
X_18910_ _18911_/CLK _18910_/D vssd1 vssd1 vccd1 vccd1 _18910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11245_ _09774_/A _11240_/X _11242_/X _11244_/X _09817_/A vssd1 vssd1 vccd1 vccd1
+ _11245_/X sky130_fd_sc_hd__a221o_1
X_19890_ _19896_/CLK _19890_/D vssd1 vssd1 vccd1 vccd1 _19890_/Q sky130_fd_sc_hd__dfxtp_1
X_18841_ _19324_/CLK _18841_/D vssd1 vssd1 vccd1 vccd1 _18841_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_121_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11176_ _11164_/A _11175_/X _11095_/A vssd1 vssd1 vccd1 vccd1 _11176_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10127_ _10497_/A vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__buf_2
XFILLER_121_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18772_ _19899_/CLK _18772_/D vssd1 vssd1 vccd1 vccd1 _18772_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16500__S _16508_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15984_ _17098_/A _16846_/B _16846_/C vssd1 vssd1 vccd1 vccd1 _17738_/B sky130_fd_sc_hd__or3_2
XFILLER_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17723_ _17723_/A vssd1 vssd1 vccd1 vccd1 _17723_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09903__A _09903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ _10058_/A vssd1 vssd1 vccd1 vccd1 _10059_/S sky130_fd_sc_hd__clkbuf_4
X_14935_ _14933_/X _14934_/X _14938_/S vssd1 vssd1 vccd1 vccd1 _14935_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17654_ _17652_/X _19724_/Q _17666_/S vssd1 vssd1 vccd1 vccd1 _17655_/A sky130_fd_sc_hd__mux2_1
X_14866_ _15029_/A vssd1 vssd1 vccd1 vccd1 _14916_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_91_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16605_ _19281_/Q _13838_/X _16613_/S vssd1 vssd1 vccd1 vccd1 _16606_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13817_ _18504_/Q _13816_/X _13820_/S vssd1 vssd1 vccd1 vccd1 _13818_/A sky130_fd_sc_hd__mux2_1
X_17585_ _17585_/A vssd1 vssd1 vccd1 vccd1 _19696_/D sky130_fd_sc_hd__clkbuf_1
X_14797_ _14800_/A _14797_/B vssd1 vssd1 vccd1 vccd1 _14798_/A sky130_fd_sc_hd__and2_1
XFILLER_63_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17331__S _17337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19324_ _19324_/CLK _19324_/D vssd1 vssd1 vccd1 vccd1 _19324_/Q sky130_fd_sc_hd__dfxtp_1
X_16536_ _16536_/A vssd1 vssd1 vccd1 vccd1 _19250_/D sky130_fd_sc_hd__clkbuf_1
X_13748_ _19025_/Q _13495_/X _13747_/Y _11730_/A vssd1 vssd1 vccd1 vccd1 _13748_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19255_ _19842_/CLK _19255_/D vssd1 vssd1 vccd1 vccd1 _19255_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14549__C1 _14540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16467_ _16467_/A vssd1 vssd1 vccd1 vccd1 _19220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13679_ _18475_/Q _13517_/X _13674_/Y _13678_/X vssd1 vssd1 vccd1 vccd1 _18475_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13160__A _17033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18206_ _17735_/X _19944_/Q _18206_/S vssd1 vssd1 vccd1 vccd1 _18207_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15418_ _15418_/A vssd1 vssd1 vccd1 vccd1 _18852_/D sky130_fd_sc_hd__clkbuf_1
X_19186_ _20035_/CLK _19186_/D vssd1 vssd1 vccd1 vccd1 _19186_/Q sky130_fd_sc_hd__dfxtp_1
X_16398_ _16398_/A vssd1 vssd1 vccd1 vccd1 _19190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12575__A1 _12554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18137_ _18193_/A vssd1 vssd1 vccd1 vccd1 _18206_/S sky130_fd_sc_hd__buf_6
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15349_ _15247_/X _14922_/X _14986_/X vssd1 vssd1 vccd1 vccd1 _15349_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10681__S0 _09726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18068_ _18067_/X _19892_/Q _18078_/S vssd1 vssd1 vccd1 vccd1 _18069_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09910_ _09910_/A vssd1 vssd1 vccd1 vccd1 _09911_/A sky130_fd_sc_hd__clkbuf_4
X_17019_ _17019_/A vssd1 vssd1 vccd1 vccd1 _19460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20030_ _20030_/CLK _20030_/D vssd1 vssd1 vccd1 vccd1 _20030_/Q sky130_fd_sc_hd__dfxtp_1
X_09841_ _09841_/A vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__buf_4
XANTENNA__10433__S0 _10328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18398__A _18409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15815__A _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _09772_/A vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10024__A _10328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10959__A _11344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13054__B _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13055__A2 _11794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17241__S _17243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09206_ _11664_/A _09272_/A vssd1 vssd1 vccd1 vccd1 _09206_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13070__A _13070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15504__A1 _18859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_135_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11030_ _09791_/A _11025_/X _11027_/Y _11029_/Y _09804_/A vssd1 vssd1 vccd1 vccd1
+ _11030_/X sky130_fd_sc_hd__o221a_1
XFILLER_103_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17416__S _17420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09723__A _10906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12981_ _18682_/Q vssd1 vssd1 vccd1 vccd1 _14355_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10869__A _15936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13294__A2 _13081_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14720_ _14720_/A vssd1 vssd1 vccd1 vccd1 _18810_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13245__A _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09442__B _09442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11932_ _11932_/A _11932_/B vssd1 vssd1 vccd1 vccd1 _11932_/X sky130_fd_sc_hd__and2_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _15715_/B vssd1 vssd1 vccd1 vccd1 _14528_/A sky130_fd_sc_hd__clkbuf_8
X_14651_ _14651_/A vssd1 vssd1 vccd1 vccd1 _18783_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _18845_/Q vssd1 vssd1 vccd1 vccd1 _10814_/Y sky130_fd_sc_hd__inv_2
X_13602_ _13602_/A vssd1 vssd1 vccd1 vccd1 _18465_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _19597_/Q _17014_/X _17376_/S vssd1 vssd1 vccd1 vccd1 _17371_/A sky130_fd_sc_hd__mux2_1
X_14582_ _14595_/A _14582_/B vssd1 vssd1 vccd1 vccd1 _14583_/A sky130_fd_sc_hd__and2_1
X_11794_ _11824_/A vssd1 vssd1 vccd1 vccd1 _11794_/X sky130_fd_sc_hd__buf_2
X_16321_ _16320_/X _19166_/Q _16330_/S vssd1 vssd1 vccd1 vccd1 _16322_/A sky130_fd_sc_hd__mux2_1
X_10745_ _09759_/A _10744_/X _10579_/A vssd1 vssd1 vccd1 vccd1 _10745_/Y sky130_fd_sc_hd__o21ai_1
X_13533_ _13528_/X _13529_/X _13531_/Y _13532_/X hold6/X vssd1 vssd1 vccd1 vccd1 hold7/A
+ sky130_fd_sc_hd__a32o_4
XANTENNA__16990__S _16990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19040_ _19637_/CLK _19040_/D vssd1 vssd1 vccd1 vccd1 _19040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16252_ _13150_/X _19139_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _16253_/A sky130_fd_sc_hd__mux2_1
X_13464_ _13463_/X _18453_/Q _13464_/S vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10676_ _10549_/A _10675_/X _09686_/A vssd1 vssd1 vccd1 vccd1 _10676_/X sky130_fd_sc_hd__o21a_1
XFILLER_139_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ _12790_/A vssd1 vssd1 vccd1 vccd1 _12415_/X sky130_fd_sc_hd__clkbuf_4
X_15203_ _15201_/X _14984_/A _15202_/X _14922_/S vssd1 vssd1 vccd1 vccd1 _15203_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_138_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16183_ _16183_/A vssd1 vssd1 vccd1 vccd1 _19109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13395_ _19907_/Q _13431_/B vssd1 vssd1 vccd1 vccd1 _13395_/X sky130_fd_sc_hd__and2_1
XFILLER_154_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15134_ _15132_/X _15095_/X _15347_/S vssd1 vssd1 vccd1 vccd1 _15134_/X sky130_fd_sc_hd__mux2_1
X_12346_ _12338_/X _12342_/X _12345_/Y vssd1 vssd1 vccd1 vccd1 _12346_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19942_ _19942_/CLK _19942_/D vssd1 vssd1 vccd1 vccd1 _19942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15065_ _14916_/X _14900_/X _15114_/S vssd1 vssd1 vccd1 vccd1 _15065_/X sky130_fd_sc_hd__mux2_1
X_12277_ _18526_/Q _12277_/B _18528_/Q _12277_/D vssd1 vssd1 vccd1 vccd1 _12340_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__12324__A _12459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14242__C _14242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14016_ _18580_/Q _14016_/B vssd1 vssd1 vccd1 vccd1 _14017_/B sky130_fd_sc_hd__and2_1
XFILLER_136_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output73_A _12301_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ _19197_/Q _19788_/Q _19950_/Q _19165_/Q _11156_/S _11108_/X vssd1 vssd1 vccd1
+ vccd1 _11228_/X sky130_fd_sc_hd__mux4_1
X_19873_ _19873_/CLK _19873_/D vssd1 vssd1 vccd1 vccd1 _19873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17326__S _17326_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18824_ _18960_/CLK _18824_/D vssd1 vssd1 vccd1 vccd1 _18824_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15635__A _15703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16230__S _16236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159_ _11237_/A _11158_/X _11227_/A vssd1 vssd1 vccd1 vccd1 _11159_/X sky130_fd_sc_hd__a21o_1
XANTENNA__18011__A _18011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18755_ _19063_/CLK _18755_/D vssd1 vssd1 vccd1 vccd1 _18755_/Q sky130_fd_sc_hd__dfxtp_1
X_15967_ _19017_/Q _15951_/X _15966_/X vssd1 vssd1 vccd1 vccd1 _19017_/D sky130_fd_sc_hd__a21o_1
XFILLER_49_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17706_ _17706_/A vssd1 vssd1 vccd1 vccd1 _19740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14918_ _15016_/A vssd1 vssd1 vccd1 vccd1 _15082_/B sky130_fd_sc_hd__clkbuf_2
X_18686_ _18687_/CLK _18686_/D vssd1 vssd1 vccd1 vccd1 _18686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15898_ _15898_/A vssd1 vssd1 vccd1 vccd1 _18992_/D sky130_fd_sc_hd__clkbuf_1
X_17637_ _17736_/S vssd1 vssd1 vccd1 vccd1 _17650_/S sky130_fd_sc_hd__buf_2
XFILLER_91_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14849_ _14990_/A _14993_/B _14849_/C vssd1 vssd1 vccd1 vccd1 _15353_/A sky130_fd_sc_hd__and3_1
XFILLER_90_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17568_ _17568_/A vssd1 vssd1 vccd1 vccd1 _19688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19307_ _19996_/CLK _19307_/D vssd1 vssd1 vccd1 vccd1 _19307_/Q sky130_fd_sc_hd__dfxtp_1
X_16519_ _19243_/Q _13819_/X _16519_/S vssd1 vssd1 vccd1 vccd1 _16520_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17996__S _17998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17499_ _17499_/A vssd1 vssd1 vccd1 vccd1 _19655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19238_ _20023_/CLK _19238_/D vssd1 vssd1 vccd1 vccd1 _19238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09949__C1 _11574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19169_ _19985_/CLK _19169_/D vssd1 vssd1 vccd1 vccd1 _19169_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10019__A _10859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16405__S _16413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12234__A _12234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20013_ _20013_/CLK _20013_/D vssd1 vssd1 vccd1 vccd1 _20013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09824_ _09824_/A vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__buf_2
XFILLER_86_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16140__S _16144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09755_ _09755_/A vssd1 vssd1 vccd1 vccd1 _11032_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13276__A2 _11815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09686_ _09686_/A vssd1 vssd1 vccd1 vccd1 _09687_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11382__S1 _11077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10530_ _10424_/A _10529_/X _10149_/A vssd1 vssd1 vccd1 vccd1 _10530_/X sky130_fd_sc_hd__a21o_1
XFILLER_167_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10461_ _19211_/Q _19802_/Q _19964_/Q _19179_/Q _10180_/S _09610_/A vssd1 vssd1 vccd1
+ vccd1 _10462_/B sky130_fd_sc_hd__mux4_1
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12200_ _12162_/A _12198_/X _12059_/X vssd1 vssd1 vccd1 vccd1 _12200_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11211__A1 _11003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13180_ _17678_/A vssd1 vssd1 vccd1 vccd1 _13180_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09718__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ _10392_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__or2_1
XFILLER_135_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12131_ _12050_/A _12124_/X _12130_/X _12056_/X vssd1 vssd1 vccd1 vccd1 _12131_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12062_ _12062_/A _12163_/B vssd1 vssd1 vccd1 vccd1 _12062_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14161__B1 _14160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11013_ _15930_/B vssd1 vssd1 vccd1 vccd1 _11459_/A sky130_fd_sc_hd__clkinv_2
X_16870_ _16329_/X _19398_/Q _16870_/S vssd1 vssd1 vccd1 vccd1 _16871_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15821_ hold2/A _15816_/X _15820_/X input64/X vssd1 vssd1 vccd1 vccd1 _15822_/B sky130_fd_sc_hd__a22o_1
XANTENNA__10599__A _10832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18540_ _18878_/CLK _18540_/D vssd1 vssd1 vccd1 vccd1 _18540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _15773_/B vssd1 vssd1 vccd1 vccd1 _15752_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _12963_/X _18426_/Q _13003_/S vssd1 vssd1 vccd1 vccd1 _12965_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _18803_/Q _13612_/X _14705_/S vssd1 vssd1 vccd1 vccd1 _14704_/A sky130_fd_sc_hd__mux2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ input66/X _11915_/B vssd1 vssd1 vccd1 vccd1 _12350_/A sky130_fd_sc_hd__nand2_2
X_18471_ _18547_/CLK _18471_/D vssd1 vssd1 vccd1 vccd1 _18471_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _15683_/A vssd1 vssd1 vccd1 vccd1 _18918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12895_/A _12956_/A vssd1 vssd1 vccd1 vccd1 _12895_/Y sky130_fd_sc_hd__nor2_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _19621_/Q _17090_/X _17424_/S vssd1 vssd1 vccd1 vccd1 _17423_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _14634_/A vssd1 vssd1 vccd1 vccd1 _18778_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _12881_/A vssd1 vssd1 vccd1 vccd1 _11847_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _17353_/A vssd1 vssd1 vccd1 vccd1 _19590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _15760_/A _11777_/B _11777_/C vssd1 vssd1 vccd1 vccd1 _11780_/B sky130_fd_sc_hd__or3_1
X_14565_ _14577_/A _14565_/B vssd1 vssd1 vccd1 vccd1 _14566_/A sky130_fd_sc_hd__and2_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _17640_/A vssd1 vssd1 vccd1 vccd1 _16304_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10728_ _09664_/A _10726_/X _11481_/A vssd1 vssd1 vccd1 vccd1 _10728_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13516_ _13520_/A vssd1 vssd1 vccd1 vccd1 _13517_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17284_ _17352_/S vssd1 vssd1 vccd1 vccd1 _17293_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__15716__B2 _15738_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14496_ _14496_/A vssd1 vssd1 vccd1 vccd1 _14501_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12038__B _15103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13849__S _13852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19023_ _19023_/CLK _19023_/D vssd1 vssd1 vccd1 vccd1 _19023_/Q sky130_fd_sc_hd__dfxtp_1
X_16235_ _16235_/A vssd1 vssd1 vccd1 vccd1 _19131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10659_ _19670_/Q _19436_/Q _18501_/Q _19766_/Q _10586_/S _10050_/A vssd1 vssd1 vccd1
+ vccd1 _10659_/X sky130_fd_sc_hd__mux4_1
X_13447_ _18894_/Q vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11202__A1 _10983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16166_ _16166_/A vssd1 vssd1 vccd1 vccd1 _19101_/D sky130_fd_sc_hd__clkbuf_1
X_13378_ _18739_/Q vssd1 vssd1 vccd1 vccd1 _14518_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13742__A3 _09341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11753__A2 _11683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15117_ _15033_/X _15028_/X _15117_/S vssd1 vssd1 vccd1 vccd1 _15117_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17845__A _17867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12950__B2 _12020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12329_ _12329_/A _12329_/B vssd1 vssd1 vccd1 vccd1 _12330_/A sky130_fd_sc_hd__or2_1
X_16097_ _16097_/A vssd1 vssd1 vccd1 vccd1 _19071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19925_ _19989_/CLK _19925_/D vssd1 vssd1 vccd1 vccd1 _19925_/Q sky130_fd_sc_hd__dfxtp_1
X_15048_ _15048_/A vssd1 vssd1 vccd1 vccd1 _15048_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17056__S _17056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19856_ _19856_/CLK _19856_/D vssd1 vssd1 vccd1 vccd1 _19856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18807_ _19887_/CLK _18807_/D vssd1 vssd1 vccd1 vccd1 _18807_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16895__S _16903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19787_ _19949_/CLK _19787_/D vssd1 vssd1 vccd1 vccd1 _19787_/Q sky130_fd_sc_hd__dfxtp_1
X_16999_ _19454_/Q _16998_/X _17008_/S vssd1 vssd1 vccd1 vccd1 _17000_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12501__B _12501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09540_ _09540_/A vssd1 vssd1 vccd1 vccd1 _09540_/X sky130_fd_sc_hd__clkbuf_4
X_18738_ _19909_/CLK _18738_/D vssd1 vssd1 vccd1 vccd1 _18738_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09331__B1 _18827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09471_ _09467_/X _14749_/B _09471_/C _14750_/B vssd1 vssd1 vccd1 vccd1 _09471_/X
+ sky130_fd_sc_hd__and4b_1
X_18669_ _18688_/CLK _18669_/D vssd1 vssd1 vccd1 vccd1 _18669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10229__C1 _09807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11116__S1 _11022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13430__A2 _18861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11133__A _11133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10972__A _10972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10627__S0 _10691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10183__S _10314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18350__S _18350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14694__A1 _13579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13497__A2 _13495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11052__S0 _10977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09807_ _09807_/A vssd1 vssd1 vccd1 vccd1 _09807_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09738_ _11157_/A vssd1 vssd1 vccd1 vccd1 _10624_/A sky130_fd_sc_hd__buf_2
XFILLER_28_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09669_ _11533_/A _09668_/X _10073_/A vssd1 vssd1 vccd1 vccd1 _09669_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _15758_/A _11700_/B vssd1 vssd1 vccd1 vccd1 _11701_/A sky130_fd_sc_hd__nor2_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12530_/X _12678_/Y _12700_/B _12583_/X vssd1 vssd1 vccd1 vccd1 _12680_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14338__B _18676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11631_ _11631_/A _11631_/B _11631_/C vssd1 vssd1 vccd1 vccd1 _11633_/B sky130_fd_sc_hd__or3_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ _11558_/A _11559_/X _11561_/X _09809_/X vssd1 vssd1 vccd1 vccd1 _11562_/X
+ sky130_fd_sc_hd__o211a_1
X_14350_ _18681_/Q _14350_/B _14350_/C vssd1 vssd1 vccd1 vccd1 _14355_/C sky130_fd_sc_hd__and3_1
XFILLER_128_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13301_ _17058_/A vssd1 vssd1 vccd1 vccd1 _17700_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10513_ _09547_/A _10502_/Y _10511_/X _10078_/X _10512_/Y vssd1 vssd1 vccd1 vccd1
+ _15956_/B sky130_fd_sc_hd__o32a_2
X_14281_ _18660_/Q _18659_/Q _18658_/Q _14281_/D vssd1 vssd1 vccd1 vccd1 _14290_/D
+ sky130_fd_sc_hd__and4_1
X_11493_ _11493_/A _11493_/B vssd1 vssd1 vccd1 vccd1 _11493_/X sky130_fd_sc_hd__or2_1
XANTENNA__16045__S _16053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10882__A _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16020_ _13202_/X _19040_/Q _16020_/S vssd1 vssd1 vccd1 vccd1 _16021_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13232_ _13092_/A _14789_/A _09354_/A input7/X _13093_/B vssd1 vssd1 vccd1 vccd1
+ _13368_/A sky130_fd_sc_hd__a41o_2
XFILLER_155_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10444_ _10444_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _10445_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09448__A _15147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11196__B1 _09911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13163_ _13163_/A vssd1 vssd1 vccd1 vccd1 _18436_/D sky130_fd_sc_hd__clkbuf_1
X_10375_ _10380_/A _10375_/B vssd1 vssd1 vccd1 vccd1 _10375_/X sky130_fd_sc_hd__or2_1
XANTENNA__17320__A0 _17151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12114_ _12114_/A vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13094_ _13094_/A vssd1 vssd1 vccd1 vccd1 _13094_/X sky130_fd_sc_hd__clkbuf_2
X_17971_ _17971_/A vssd1 vssd1 vccd1 vccd1 _19853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13488__A2 _12881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19710_ _20003_/CLK _19710_/D vssd1 vssd1 vccd1 vccd1 _19710_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output159_A _12681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12045_ _11993_/A _11993_/B _12044_/Y vssd1 vssd1 vccd1 vccd1 _12046_/B sky130_fd_sc_hd__o21a_2
X_16922_ _16990_/S vssd1 vssd1 vccd1 vccd1 _16931_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10821__S _10821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13000__A1_N _12967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09375__B_N _18951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19641_ _19641_/CLK _19641_/D vssd1 vssd1 vccd1 vccd1 _19641_/Q sky130_fd_sc_hd__dfxtp_1
X_16853_ _16304_/X _19390_/Q _16859_/S vssd1 vssd1 vccd1 vccd1 _16854_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17604__S _17606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15804_ _15804_/A vssd1 vssd1 vccd1 vccd1 _18964_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12448__A0 _12443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19572_ _19829_/CLK _19572_/D vssd1 vssd1 vccd1 vccd1 _19572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10122__A _11467_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16784_ _16326_/X _19360_/Q _16786_/S vssd1 vssd1 vccd1 vccd1 _16785_/A sky130_fd_sc_hd__mux2_1
X_13996_ _18573_/Q _13999_/C _13995_/Y vssd1 vssd1 vccd1 vccd1 _18573_/D sky130_fd_sc_hd__o21a_1
XFILLER_46_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18523_ _18997_/CLK _18523_/D vssd1 vssd1 vccd1 vccd1 _18523_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09911__A _09911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735_ _15735_/A vssd1 vssd1 vccd1 vccd1 _16691_/A sky130_fd_sc_hd__buf_4
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _13209_/B vssd1 vssd1 vccd1 vccd1 _13373_/B sky130_fd_sc_hd__buf_2
XFILLER_46_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14529__A _14529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11120__B1 _09911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _19975_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15666_ _18911_/Q _12416_/B _15666_/S vssd1 vssd1 vccd1 vccd1 _15667_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15937__A1 _19005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12878_/A vssd1 vssd1 vccd1 vccd1 _12878_/X sky130_fd_sc_hd__buf_2
XFILLER_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17405_ _19613_/Q _17065_/X _17409_/S vssd1 vssd1 vccd1 vccd1 _17406_/A sky130_fd_sc_hd__mux2_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17139__A0 _17138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14617_ _14617_/A vssd1 vssd1 vccd1 vccd1 _18773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18385_ _17681_/X _20023_/Q _18385_/S vssd1 vssd1 vccd1 vccd1 _18386_/A sky130_fd_sc_hd__mux2_1
X_11829_ _14552_/A vssd1 vssd1 vccd1 vccd1 _13726_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13412__A2 _18860_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15597_ _15597_/A vssd1 vssd1 vccd1 vccd1 _18880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _17336_/A vssd1 vssd1 vccd1 vccd1 _19582_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10857__S0 _11488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14548_ _14548_/A _14547_/X vssd1 vssd1 vccd1 vccd1 _14548_/X sky130_fd_sc_hd__or2b_1
XFILLER_174_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11888__A _13081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17267_ _17267_/A vssd1 vssd1 vccd1 vccd1 _17276_/S sky130_fd_sc_hd__buf_4
X_14479_ _14479_/A vssd1 vssd1 vccd1 vccd1 _14514_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19006_ _19025_/CLK _19006_/D vssd1 vssd1 vccd1 vccd1 _19006_/Q sky130_fd_sc_hd__dfxtp_2
X_16218_ _16218_/A vssd1 vssd1 vccd1 vccd1 _19125_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09358__A _13091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10609__S0 _10657_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17198_ _17735_/A vssd1 vssd1 vccd1 vccd1 _17198_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17311__A0 _17138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__S1 _10028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16149_ _16149_/A vssd1 vssd1 vccd1 vccd1 _19095_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17575__A _17632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__S0 _11063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19908_ _19909_/CLK _19908_/D vssd1 vssd1 vccd1 vccd1 _19908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19839_ _19839_/CLK _19839_/D vssd1 vssd1 vccd1 vccd1 _19839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09821__A _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09523_ _09309_/A _09522_/Y _09520_/B vssd1 vssd1 vccd1 vccd1 _11937_/B sky130_fd_sc_hd__a21o_1
XFILLER_25_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13651__A2 _11764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13343__A _17065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09454_ _14749_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _12055_/A sky130_fd_sc_hd__or2_1
XFILLER_101_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11662__A1 _11650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09385_ _09401_/A vssd1 vssd1 vccd1 vccd1 _11869_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11798__A _11831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10906__S _10906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10207__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10925__B1 _10719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10160_ _10438_/A _10158_/X _10159_/X vssd1 vssd1 vccd1 vccd1 _10160_/X sky130_fd_sc_hd__o21a_1
XANTENNA__15717__B _15740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14667__A1 _13750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15864__B1 _15788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _10084_/Y _10086_/Y _10088_/Y _10090_/Y _09823_/A vssd1 vssd1 vccd1 vccd1
+ _10091_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09769__S1 _09768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17424__S _17424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13850_ _13850_/A vssd1 vssd1 vccd1 vccd1 _18514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09731__A _10277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ _18548_/Q _12790_/X _12796_/X _12800_/X vssd1 vssd1 vccd1 vccd1 _12801_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_28_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13781_ _17017_/A vssd1 vssd1 vccd1 vccd1 _13781_/X sky130_fd_sc_hd__buf_2
X_10993_ _11001_/A _10993_/B vssd1 vssd1 vccd1 vccd1 _10993_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15520_ _15520_/A _15520_/B vssd1 vssd1 vccd1 vccd1 _15520_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15919__A1 _15053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12732_ _12645_/B _12670_/A _12729_/X _12731_/X vssd1 vssd1 vccd1 vccd1 _12742_/A
+ sky130_fd_sc_hd__a31o_2
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _15522_/A _15451_/B _15451_/C vssd1 vssd1 vccd1 vccd1 _15451_/X sky130_fd_sc_hd__and3_1
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _15970_/C _18922_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12664_/A sky130_fd_sc_hd__mux2_2
XANTENNA__18255__S _18263_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14402_ _14413_/A _14409_/C vssd1 vssd1 vccd1 vccd1 _14402_/Y sky130_fd_sc_hd__nor2_1
X_18170_ _18170_/A vssd1 vssd1 vccd1 vccd1 _19927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11614_ _11614_/A _11614_/B _11614_/C _11613_/X vssd1 vssd1 vccd1 vccd1 _11614_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12602__A0 _12599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15382_ _15368_/X _15385_/B _15369_/X _15381_/X vssd1 vssd1 vccd1 vccd1 _15382_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12619_/A _12618_/A vssd1 vssd1 vccd1 vccd1 _12595_/A sky130_fd_sc_hd__xor2_1
XFILLER_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ _17121_/A vssd1 vssd1 vccd1 vccd1 _19496_/D sky130_fd_sc_hd__clkbuf_1
X_14333_ _14336_/B _14338_/D _14332_/X vssd1 vssd1 vccd1 vccd1 _14333_/Y sky130_fd_sc_hd__a21oi_1
X_11545_ _11547_/A _11545_/B vssd1 vssd1 vccd1 vccd1 _11545_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13158__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17052_ _17052_/A vssd1 vssd1 vccd1 vccd1 _17052_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11476_ _19926_/Q _19540_/Q _19990_/Q _19109_/Q _10708_/X _10710_/X vssd1 vssd1 vccd1
+ vccd1 _11477_/B sky130_fd_sc_hd__mux4_1
X_14264_ _18656_/Q _18655_/Q _18654_/Q _14264_/D vssd1 vssd1 vccd1 vccd1 _14275_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_143_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11169__B1 _15923_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16003_ _13042_/X _19032_/Q _16009_/S vssd1 vssd1 vccd1 vccd1 _16004_/A sky130_fd_sc_hd__mux2_1
X_10427_ _10172_/A _10422_/X _10424_/Y _10426_/Y vssd1 vssd1 vccd1 vccd1 _10427_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__18097__A1 _13667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ _18848_/Q _13627_/B _13215_/S vssd1 vssd1 vccd1 vccd1 _13215_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ _14407_/A vssd1 vssd1 vccd1 vccd1 _14315_/A sky130_fd_sc_hd__buf_2
XFILLER_125_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10358_ _10200_/A _10353_/X _10355_/X _10357_/X vssd1 vssd1 vccd1 vccd1 _10358_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_151_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09906__A _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13146_ _13142_/Y _13174_/C _13144_/X _13289_/A vssd1 vssd1 vccd1 vccd1 _13146_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17954_ _18352_/C _17954_/B vssd1 vssd1 vccd1 vccd1 _18011_/A sky130_fd_sc_hd__nor2_4
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _18798_/Q _13071_/X _13074_/X _13076_/Y vssd1 vssd1 vccd1 vccd1 _13077_/X
+ sky130_fd_sc_hd__a211o_2
XANTENNA__11016__S0 _11017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10289_ _20032_/Q _19870_/Q _19279_/Q _19049_/Q _10279_/X _10283_/X vssd1 vssd1 vccd1
+ vccd1 _10290_/B sky130_fd_sc_hd__mux4_1
XFILLER_112_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16905_ _16905_/A vssd1 vssd1 vccd1 vccd1 _16914_/S sky130_fd_sc_hd__buf_4
X_12028_ _11997_/X _12024_/Y _12027_/X vssd1 vssd1 vccd1 vccd1 _12028_/X sky130_fd_sc_hd__a21o_4
XANTENNA__15786__D_N input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17885_ _19815_/Q _16992_/X _17893_/S vssd1 vssd1 vccd1 vccd1 _17886_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19624_ _19979_/CLK _19624_/D vssd1 vssd1 vccd1 vccd1 _19624_/Q sky130_fd_sc_hd__dfxtp_1
X_16836_ _16836_/A vssd1 vssd1 vccd1 vccd1 _17201_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _20013_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09641__A _11538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19555_ _20037_/CLK _19555_/D vssd1 vssd1 vccd1 vccd1 _19555_/Q sky130_fd_sc_hd__dfxtp_1
X_16767_ _16297_/X _19352_/Q _16775_/S vssd1 vssd1 vccd1 vccd1 _16768_/A sky130_fd_sc_hd__mux2_1
X_13979_ _18567_/Q _13982_/C _13969_/X vssd1 vssd1 vccd1 vccd1 _13979_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14259__A _14265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18506_ _19771_/CLK _18506_/D vssd1 vssd1 vccd1 vccd1 _18506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15718_ _09436_/B _15705_/X _15717_/X _15713_/X vssd1 vssd1 vccd1 vccd1 _18934_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19486_ _19487_/CLK _19486_/D vssd1 vssd1 vccd1 vccd1 _19486_/Q sky130_fd_sc_hd__dfxtp_1
X_16698_ _16698_/A vssd1 vssd1 vccd1 vccd1 _19321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18437_ _19636_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15649_ _18903_/Q _12191_/A _15655_/S vssd1 vssd1 vccd1 vccd1 _15650_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18165__S _18169_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16474__A _16691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09170_ _18965_/Q vssd1 vssd1 vccd1 vccd1 _09283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18368_ _17656_/X _20015_/Q _18374_/S vssd1 vssd1 vccd1 vccd1 _18369_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17319_ _17319_/A vssd1 vssd1 vccd1 vccd1 _19574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10726__S _10821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18299_ _18299_/A vssd1 vssd1 vccd1 vccd1 _19984_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12507__A _12508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12619__B_N _15449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__B1 _10078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14897__A1 _12738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18088__A1 _11748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16413__S _16413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17835__A1 _17026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10383__A1 _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14649__A1 _13710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11007__S0 _11048_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13338__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13772__S _13772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15553__A _15553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10230__S1 _10223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13085__A0 _18841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09506_ _14765_/A _09506_/B vssd1 vssd1 vccd1 vccd1 _09508_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16023__A0 _13219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09437_ _09437_/A vssd1 vssd1 vccd1 vccd1 _14761_/C sky130_fd_sc_hd__clkbuf_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15782__C1 _13885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09368_ _18956_/Q _18954_/Q _18953_/Q vssd1 vssd1 vccd1 vccd1 _11680_/B sky130_fd_sc_hd__or3_1
XANTENNA__11494__S0 _10906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09299_ _18980_/Q _18979_/Q _18978_/Q _18977_/Q vssd1 vssd1 vccd1 vccd1 _09465_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_165_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11330_ _11421_/A _11330_/B vssd1 vssd1 vccd1 vccd1 _11330_/X sky130_fd_sc_hd__or2_1
XFILLER_126_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15728__A _16150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ _11122_/A _11258_/X _11260_/X vssd1 vssd1 vccd1 vccd1 _11261_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18104__A _18104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ _10748_/A vssd1 vssd1 vccd1 vccd1 _10695_/A sky130_fd_sc_hd__clkbuf_2
X_13000_ _12967_/X _12999_/X _12906_/A input27/X vssd1 vssd1 vccd1 vccd1 _17007_/A
+ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__09726__A _09726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11192_ _11340_/A _11191_/X _09789_/A vssd1 vssd1 vccd1 vccd1 _11192_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11467__S _11467_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15837__B1 _15789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ _19940_/Q _19554_/Q _20004_/Q _19123_/Q _10141_/X _10283_/A vssd1 vssd1 vccd1
+ vccd1 _10144_/B sky130_fd_sc_hd__mux4_1
XFILLER_43_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10074_ _20033_/Q _19871_/Q _19280_/Q _19050_/Q _09597_/A _09646_/A vssd1 vssd1 vccd1
+ vccd1 _10074_/X sky130_fd_sc_hd__mux4_1
XANTENNA_input35_A io_ibus_inst[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14951_ _14946_/X _14949_/X _15121_/S vssd1 vssd1 vccd1 vccd1 _14951_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13902_ _18542_/Q _13900_/X _12651_/X _12655_/X _13897_/X vssd1 vssd1 vccd1 vccd1
+ _18542_/D sky130_fd_sc_hd__o221a_1
X_17670_ _17668_/X _19729_/Q _17682_/S vssd1 vssd1 vccd1 vccd1 _17671_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14882_ _14878_/X _14881_/X _14916_/S vssd1 vssd1 vccd1 vccd1 _14882_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11874__B2 _18669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16621_ _16689_/S vssd1 vssd1 vccd1 vccd1 _16630_/S sky130_fd_sc_hd__buf_2
X_13833_ _18509_/Q _13832_/X _13836_/S vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13076__B1 _09410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19340_ _19997_/CLK _19340_/D vssd1 vssd1 vccd1 vccd1 _19340_/Q sky130_fd_sc_hd__dfxtp_1
X_16552_ _19257_/Q _13762_/X _16558_/S vssd1 vssd1 vccd1 vccd1 _16553_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10400__A _10400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13764_ _13764_/A vssd1 vssd1 vccd1 vccd1 _18487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _11409_/S vssd1 vssd1 vccd1 vccd1 _10977_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_31_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15503_ _12693_/Y _15458_/X _15502_/X _15454_/X vssd1 vssd1 vccd1 vccd1 _15503_/X
+ sky130_fd_sc_hd__a211o_1
X_19271_ _19960_/CLK _19271_/D vssd1 vssd1 vccd1 vccd1 _19271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12715_ _12715_/A vssd1 vssd1 vccd1 vccd1 _15498_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16483_ _16483_/A vssd1 vssd1 vccd1 vccd1 _19226_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16565__A1 _13781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13695_ _13699_/B _13694_/Y _13648_/X vssd1 vssd1 vccd1 vccd1 _13695_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_94_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14576__A0 _12165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18222_ _19950_/Q _17652_/A _18230_/S vssd1 vssd1 vccd1 vccd1 _18223_/A sky130_fd_sc_hd__mux2_1
X_15434_ _15155_/X _15436_/B _15102_/X _15433_/X vssd1 vssd1 vccd1 vccd1 _15434_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12646_ _18542_/Q _12647_/B vssd1 vssd1 vccd1 vccd1 _12648_/A sky130_fd_sc_hd__nor2_1
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09678__S0 _09920_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18153_ _18153_/A vssd1 vssd1 vccd1 vccd1 _19919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15365_ _15365_/A vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12577_ _12577_/A _12623_/C vssd1 vssd1 vccd1 vccd1 _12577_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17104_ _17103_/X _19491_/Q _17113_/S vssd1 vssd1 vccd1 vccd1 _17105_/A sky130_fd_sc_hd__mux2_1
X_14316_ _18670_/Q _14316_/B _14317_/D vssd1 vssd1 vccd1 vccd1 _14316_/X sky130_fd_sc_hd__and3_1
X_11528_ _15980_/B _12864_/C vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__nand2_1
X_18084_ _18849_/Q _11724_/X _18084_/S vssd1 vssd1 vccd1 vccd1 _18084_/X sky130_fd_sc_hd__mux2_1
X_15296_ _12301_/X _15279_/X _15295_/X _15275_/X vssd1 vssd1 vccd1 vccd1 _15296_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17329__S _17337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17035_ _17035_/A vssd1 vssd1 vccd1 vccd1 _19465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14247_ _14265_/A _14247_/B vssd1 vssd1 vccd1 vccd1 _14247_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14542__A input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11459_ _11459_/A _12834_/A vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__or2_1
XANTENNA__12354__A2 _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09636__A _09636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_140_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18724_/CLK sky130_fd_sc_hd__clkbuf_16
X_14178_ _18631_/Q _14180_/C _14177_/Y vssd1 vssd1 vccd1 vccd1 _18631_/D sky130_fd_sc_hd__o21a_1
XFILLER_140_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _18843_/Q _13588_/B _13349_/S vssd1 vssd1 vccd1 vccd1 _13129_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _18992_/CLK _18986_/D vssd1 vssd1 vccd1 vccd1 _18986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17937_ _19839_/Q _17071_/X _17937_/S vssd1 vssd1 vccd1 vccd1 _17938_/A sky130_fd_sc_hd__mux2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11314__B1 _09881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17868_ _19808_/Q _17074_/X _17876_/S vssd1 vssd1 vccd1 vccd1 _17869_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_155_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19887_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09371__A _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19607_ _19976_/CLK _19607_/D vssd1 vssd1 vccd1 vccd1 _19607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16819_ _16377_/X _19376_/Q _16819_/S vssd1 vssd1 vccd1 vccd1 _16820_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17799_ _17799_/A vssd1 vssd1 vccd1 vccd1 _19777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12814__A0 _12812_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19538_ _19990_/CLK _19538_/D vssd1 vssd1 vccd1 vccd1 _19538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19469_ _20025_/CLK _19469_/D vssd1 vssd1 vccd1 vccd1 _19469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09691__C1 _09690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14567__A0 _12020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09222_ _09306_/A _09480_/A vssd1 vssd1 vccd1 vccd1 _11659_/B sky130_fd_sc_hd__or2_1
XFILLER_148_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17239__S _17243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11228__S0 _11156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15548__A _15624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10980__A _10980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_108_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _20002_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09546__A _09546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13068__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09986_ _19249_/Q _19744_/Q _10251_/S vssd1 vssd1 vccd1 vccd1 _09986_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18233__A1 _17668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17702__S _17714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10830_ _09686_/A _10825_/X _10827_/Y _10829_/Y _09874_/A vssd1 vssd1 vccd1 vccd1
+ _10830_/X sky130_fd_sc_hd__o221a_2
XANTENNA_clkbuf_leaf_131_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10220__A _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10761_ _10759_/X _10761_/B vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__and2b_1
XANTENNA__12281__A1 _18464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16318__S _16330_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13531__A _13531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12500_ _12501_/B _12524_/C vssd1 vssd1 vccd1 vccd1 _12502_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10692_ _10522_/A _10691_/X _10630_/A vssd1 vssd1 vccd1 vccd1 _10692_/Y sky130_fd_sc_hd__a21oi_1
X_13480_ _17090_/A vssd1 vssd1 vccd1 vccd1 _17732_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12033__A1 _12032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ _12514_/A vssd1 vssd1 vccd1 vccd1 _15373_/A sky130_fd_sc_hd__buf_2
XFILLER_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15150_ _18837_/Q _15053_/X _15145_/X _15149_/X vssd1 vssd1 vccd1 vccd1 _18837_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_154_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12362_ _12362_/A vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__clkinv_2
XFILLER_165_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11792__B1 _12876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14101_ _18609_/Q _14097_/B _14100_/Y vssd1 vssd1 vccd1 vccd1 _18609_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17149__S _17161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11313_ _09803_/A _11299_/X _11303_/Y _11307_/Y _11312_/X vssd1 vssd1 vccd1 vccd1
+ _11313_/X sky130_fd_sc_hd__a32o_1
XANTENNA__15458__A _15458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10890__A _18843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12293_ _11904_/A _12839_/B _12292_/X vssd1 vssd1 vccd1 vccd1 _15291_/A sky130_fd_sc_hd__a21o_2
XANTENNA__11219__S0 _11063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15081_ _15369_/A vssd1 vssd1 vccd1 vccd1 _15081_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16053__S _16053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14032_ _14034_/B _14034_/C _14019_/X vssd1 vssd1 vccd1 vccd1 _14032_/Y sky130_fd_sc_hd__a21oi_1
X_11244_ _09755_/A _11243_/X _11095_/A vssd1 vssd1 vccd1 vccd1 _11244_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13533__B2 hold6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15177__B _15177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10347__A1 _10162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16988__S _16990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ _20013_/Q _19851_/Q _19260_/Q _19030_/Q _11348_/S _11015_/A vssd1 vssd1 vccd1
+ vccd1 _11175_/X sky130_fd_sc_hd__mux4_1
X_18840_ _19324_/CLK _18840_/D vssd1 vssd1 vccd1 vccd1 _18840_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10126_ _10448_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _10126_/X sky130_fd_sc_hd__and2_1
XFILLER_110_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_72_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19877_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18771_ _19899_/CLK _18771_/D vssd1 vssd1 vccd1 vccd1 _18771_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output141_A _11908_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15983_ _19025_/Q _15936_/A _15928_/A _15982_/Y vssd1 vssd1 vccd1 vccd1 _19025_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17722_ _17722_/A vssd1 vssd1 vccd1 vccd1 _19745_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18224__A1 _17656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ _10057_/A _10057_/B vssd1 vssd1 vccd1 vccd1 _10057_/Y sky130_fd_sc_hd__nand2_1
X_14934_ _12618_/A _15254_/B _14937_/S vssd1 vssd1 vccd1 vccd1 _14934_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17653_ _17736_/S vssd1 vssd1 vccd1 vccd1 _17666_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14865_ _14865_/A vssd1 vssd1 vccd1 vccd1 _15029_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_87_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 _19965_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16604_ _16604_/A vssd1 vssd1 vccd1 vccd1 _16613_/S sky130_fd_sc_hd__buf_4
X_13816_ _17052_/A vssd1 vssd1 vccd1 vccd1 _13816_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15921__A _15982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17584_ _17128_/X _19696_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17585_/A sky130_fd_sc_hd__mux2_1
X_14796_ _12866_/B _14748_/X _14789_/B _18831_/Q vssd1 vssd1 vccd1 vccd1 _14797_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ _19485_/CLK _19323_/D vssd1 vssd1 vccd1 vccd1 _19323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16535_ _19250_/Q _13842_/X _16541_/S vssd1 vssd1 vccd1 vccd1 _16536_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13747_ _13747_/A _19025_/Q vssd1 vssd1 vccd1 vccd1 _13747_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16228__S _16236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10959_ _11344_/A vssd1 vssd1 vccd1 vccd1 _11149_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19254_ _20039_/CLK _19254_/D vssd1 vssd1 vccd1 vccd1 _19254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_10_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19982_/CLK sky130_fd_sc_hd__clkbuf_16
X_16466_ _19220_/Q _13848_/X _16468_/S vssd1 vssd1 vccd1 vccd1 _16467_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13678_ _13650_/X _13677_/X _13517_/A vssd1 vssd1 vccd1 vccd1 _13678_/X sky130_fd_sc_hd__a21bo_1
XANTENNA_clkbuf_opt_3_0_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18205_ _18205_/A vssd1 vssd1 vccd1 vccd1 _19943_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13221__A0 _13219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15417_ _18852_/Q _15416_/X _15480_/S vssd1 vssd1 vccd1 vccd1 _15418_/A sky130_fd_sc_hd__mux2_1
X_19185_ _19873_/CLK _19185_/D vssd1 vssd1 vccd1 vccd1 _19185_/Q sky130_fd_sc_hd__dfxtp_1
X_12629_ _18780_/Q _12606_/X _12170_/X vssd1 vssd1 vccd1 vccd1 _12629_/Y sky130_fd_sc_hd__o21ai_1
X_16397_ _16396_/X _19190_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _16398_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18136_ _18352_/A _18352_/B _18280_/B vssd1 vssd1 vccd1 vccd1 _18193_/A sky130_fd_sc_hd__or3_4
XFILLER_8_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15348_ _15346_/Y _15347_/X _15348_/S vssd1 vssd1 vccd1 vccd1 _15348_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_25_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19569_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18067_ _18844_/Q _11833_/D _18067_/S vssd1 vssd1 vccd1 vccd1 _18067_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15368__A _15368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16710__A1 _13781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15279_ _15458_/A vssd1 vssd1 vccd1 vccd1 _15279_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10681__S1 _10010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13524__A1 _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17018_ _19460_/Q _17017_/X _17024_/S vssd1 vssd1 vccd1 vccd1 _17019_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10338__A1 _09798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _19485_/Q _09909_/B _09909_/C vssd1 vssd1 vccd1 vccd1 _09841_/A sky130_fd_sc_hd__and3_1
XFILLER_140_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15277__A1 _18843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _11181_/A vssd1 vssd1 vccd1 vccd1 _09772_/A sky130_fd_sc_hd__buf_2
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _18998_/CLK _18969_/D vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfxtp_2
XFILLER_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13335__B _13335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16138__S _16144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10274__B1 _09540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09205_ _09283_/A vssd1 vssd1 vccd1 vccd1 _11664_/A sky130_fd_sc_hd__inv_2
XANTENNA__14881__S _14948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13212__B1 _11794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15278__A _15457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10215__A _10521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_clock clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09969_ _10266_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _09969_/X sky130_fd_sc_hd__or2_1
XANTENNA__13279__B1 _13005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ _12980_/A vssd1 vssd1 vccd1 vccd1 _18427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10869__B _12839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11931_ _09289_/A _14819_/A _11931_/C vssd1 vssd1 vccd1 vccd1 _11931_/X sky130_fd_sc_hd__and3b_1
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10501__A1 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14663_/A _14650_/B vssd1 vssd1 vccd1 vccd1 _14651_/A sky130_fd_sc_hd__and2_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _18711_/Q _14792_/B _11860_/X _11861_/X vssd1 vssd1 vccd1 vccd1 _18713_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _18465_/Q _13600_/X _13617_/S vssd1 vssd1 vccd1 vccd1 _13602_/A sky130_fd_sc_hd__mux2_1
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10813_ _09794_/A _10804_/Y _10808_/Y _10812_/Y _09804_/A vssd1 vssd1 vccd1 vccd1
+ _10813_/X sky130_fd_sc_hd__o311a_2
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14581_ _18763_/Q _13553_/X _14581_/S vssd1 vssd1 vccd1 vccd1 _14582_/B sky130_fd_sc_hd__mux2_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _13057_/A vssd1 vssd1 vccd1 vccd1 _11851_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16320_ _17656_/A vssd1 vssd1 vccd1 vccd1 _16320_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13532_ _13660_/A vssd1 vssd1 vccd1 vccd1 _13532_/X sky130_fd_sc_hd__clkbuf_2
X_10744_ _19206_/Q _19797_/Q _19959_/Q _19174_/Q _10750_/S _10626_/A vssd1 vssd1 vccd1
+ vccd1 _10744_/X sky130_fd_sc_hd__mux4_1
XANTENNA__18390__A0 _17688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16251_ _16251_/A vssd1 vssd1 vccd1 vccd1 _19138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17668__A _17668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13463_ _17729_/A vssd1 vssd1 vccd1 vccd1 _13463_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10675_ _20024_/Q _19862_/Q _19271_/Q _19041_/Q _09652_/A _10656_/A vssd1 vssd1 vccd1
+ vccd1 _10675_/X sky130_fd_sc_hd__mux4_1
XANTENNA__18263__S _18263_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15202_ _15121_/X _15118_/X _15202_/S vssd1 vssd1 vccd1 vccd1 _15202_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12414_ _18533_/Q vssd1 vssd1 vccd1 vccd1 _12416_/C sky130_fd_sc_hd__buf_2
X_16182_ _13180_/X _19109_/Q _16184_/S vssd1 vssd1 vccd1 vccd1 _16183_/A sky130_fd_sc_hd__mux2_1
X_13394_ _13188_/A _18859_/Q _12957_/X vssd1 vssd1 vccd1 vccd1 _13394_/Y sky130_fd_sc_hd__a21oi_1
X_15133_ _15169_/A vssd1 vssd1 vccd1 vccd1 _15347_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12345_ _18466_/Q _12343_/X _12344_/X vssd1 vssd1 vccd1 vccd1 _12345_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19941_ _19941_/CLK _19941_/D vssd1 vssd1 vccd1 vccd1 _19941_/Q sky130_fd_sc_hd__dfxtp_1
X_15064_ _15062_/X _15063_/X _15199_/S vssd1 vssd1 vccd1 vccd1 _15064_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12276_ _12234_/A _12277_/B _12277_/D _18528_/Q vssd1 vssd1 vccd1 vccd1 _12278_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_153_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14015_ _18579_/Q _14010_/B _14014_/Y vssd1 vssd1 vccd1 vccd1 _18579_/D sky130_fd_sc_hd__o21a_1
XFILLER_141_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11227_ _11227_/A _11227_/B vssd1 vssd1 vccd1 vccd1 _11227_/X sky130_fd_sc_hd__or2_1
XANTENNA__16511__S _16519_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19872_ _20002_/CLK _19872_/D vssd1 vssd1 vccd1 vccd1 _19872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09914__A _18862_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18823_ _18960_/CLK _18823_/D vssd1 vssd1 vccd1 vccd1 _18823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11158_ _19230_/Q _19725_/Q _11158_/S vssd1 vssd1 vccd1 vccd1 _11158_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15127__S _15127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ _10398_/A vssd1 vssd1 vccd1 vccd1 _10109_/X sky130_fd_sc_hd__buf_2
X_15966_ _15966_/A _15966_/B _15966_/C vssd1 vssd1 vccd1 vccd1 _15966_/X sky130_fd_sc_hd__and3_1
X_11089_ _19386_/Q vssd1 vssd1 vccd1 vccd1 _11440_/A sky130_fd_sc_hd__clkbuf_1
X_18754_ _18956_/CLK _18754_/D vssd1 vssd1 vccd1 vccd1 _18754_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12340__A _12340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17705_ _17704_/X _19740_/Q _17714_/S vssd1 vssd1 vccd1 vccd1 _17706_/A sky130_fd_sc_hd__mux2_1
X_14917_ _14911_/X _14916_/X _15118_/S vssd1 vssd1 vccd1 vccd1 _14917_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18685_ _19882_/CLK _18685_/D vssd1 vssd1 vccd1 vccd1 _18685_/Q sky130_fd_sc_hd__dfxtp_1
X_15897_ _15897_/A _15897_/B vssd1 vssd1 vccd1 vccd1 _15898_/A sky130_fd_sc_hd__and2_1
XFILLER_64_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09894__C1 _11574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17342__S _17348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17636_ _17717_/A vssd1 vssd1 vccd1 vccd1 _17736_/S sky130_fd_sc_hd__buf_6
XFILLER_1_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14848_ _14973_/B vssd1 vssd1 vccd1 vccd1 _14849_/C sky130_fd_sc_hd__clkinv_2
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15431__A1 _18853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17567_ _17103_/X _19688_/Q _17573_/S vssd1 vssd1 vccd1 vccd1 _17568_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10795__A _10858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14779_ _14748_/X _14766_/A _14789_/B _18826_/Q vssd1 vssd1 vccd1 vccd1 _14780_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14267__A _14745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19306_ _19994_/CLK _19306_/D vssd1 vssd1 vccd1 vccd1 _19306_/Q sky130_fd_sc_hd__dfxtp_1
X_16518_ _16518_/A vssd1 vssd1 vccd1 vccd1 _19242_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17498_ _19655_/Q vssd1 vssd1 vccd1 vccd1 _17499_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16449_ _19212_/Q _13822_/X _16457_/S vssd1 vssd1 vccd1 vccd1 _16450_/A sky130_fd_sc_hd__mux2_1
X_19237_ _19732_/CLK _19237_/D vssd1 vssd1 vccd1 vccd1 _19237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19168_ _19985_/CLK _19168_/D vssd1 vssd1 vccd1 vccd1 _19168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10559__A1 _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18133__B1 _16075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__B1 _13451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18119_ _18118_/X _19907_/Q _18128_/S vssd1 vssd1 vccd1 vccd1 _18120_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19099_ _19979_/CLK _19099_/D vssd1 vssd1 vccd1 vccd1 _19099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12234__B _12234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20012_ _20012_/CLK _20012_/D vssd1 vssd1 vccd1 vccd1 _20012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09823_ _09823_/A vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09754_ _11311_/A vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__buf_2
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12484__A1 _12422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ _09685_/A vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__buf_2
XFILLER_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18348__S _18350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17252__S _17254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10590__S0 _10657_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12236__B2 _18990_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13433__B1 _12879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15973__A2 _14803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13081__A _13081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14933__A0 _12641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10460_ _10415_/A _10459_/X _09565_/A vssd1 vssd1 vccd1 vccd1 _10460_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18124__A0 _18861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10391_ _19149_/Q _19410_/Q _19309_/Q _19644_/Q _10469_/S _09745_/A vssd1 vssd1 vccd1
+ vccd1 _10392_/B sky130_fd_sc_hd__mux4_2
XFILLER_164_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14749__C_N _09467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10645__S1 _10638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__A _12583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12130_ _15633_/C _12153_/B _12153_/C _12130_/D vssd1 vssd1 vccd1 vccd1 _12130_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12061_ _12061_/A _12066_/A _12066_/B vssd1 vssd1 vccd1 vccd1 _12163_/B sky130_fd_sc_hd__or3_2
XANTENNA__15736__A _16691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09734__A _19385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11012_ _11291_/A _10999_/X _11010_/X _10078_/A _11011_/Y vssd1 vssd1 vccd1 vccd1
+ _15930_/B sky130_fd_sc_hd__o32a_4
XFILLER_104_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15820_ _15834_/A vssd1 vssd1 vccd1 vccd1 _15820_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12160__A _18763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15751_ _11982_/X _15734_/X _15750_/X _15743_/X vssd1 vssd1 vccd1 vccd1 _18946_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12963_ _17643_/A vssd1 vssd1 vccd1 vccd1 _12963_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14702_ _14702_/A vssd1 vssd1 vccd1 vccd1 _18802_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10486__B1 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11914_ _12275_/A vssd1 vssd1 vccd1 vccd1 _12503_/A sky130_fd_sc_hd__clkbuf_2
X_18470_ _19900_/CLK _18470_/D vssd1 vssd1 vccd1 vccd1 _18470_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _18918_/Q _18539_/Q _15688_/S vssd1 vssd1 vccd1 vccd1 _15683_/A sky130_fd_sc_hd__mux2_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12894_ _13215_/S vssd1 vssd1 vccd1 vccd1 _12956_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17421_/A vssd1 vssd1 vccd1 vccd1 _19620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14633_ _14646_/A _14633_/B vssd1 vssd1 vccd1 vccd1 _14634_/A sky130_fd_sc_hd__and2_1
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _13290_/B vssd1 vssd1 vccd1 vccd1 _11845_/X sky130_fd_sc_hd__buf_2
XANTENNA__10819__S _10821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output104_A _14791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17352_ _17198_/X _19590_/Q _17352_/S vssd1 vssd1 vccd1 vccd1 _17353_/A sky130_fd_sc_hd__mux2_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _18758_/Q _14562_/X _14581_/S vssd1 vssd1 vccd1 vccd1 _14565_/B sky130_fd_sc_hd__mux2_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11776_ _13194_/A vssd1 vssd1 vccd1 vccd1 _11776_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16303_/A vssd1 vssd1 vccd1 vccd1 _19160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13515_ _13515_/A vssd1 vssd1 vccd1 vccd1 _18456_/D sky130_fd_sc_hd__clkbuf_1
X_10727_ _10727_/A vssd1 vssd1 vccd1 vccd1 _11481_/A sky130_fd_sc_hd__clkbuf_2
X_17283_ _17339_/A vssd1 vssd1 vccd1 vccd1 _17352_/S sky130_fd_sc_hd__buf_6
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16506__S _16508_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15716__A2 _14803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11450__A2 _11438_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14495_ _14495_/A _14495_/B _14495_/C vssd1 vssd1 vccd1 vccd1 _18731_/D sky130_fd_sc_hd__nor3_1
XFILLER_146_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19022_ _19023_/CLK _19022_/D vssd1 vssd1 vccd1 vccd1 _19022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14924__A0 _15410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16234_ _12978_/X _19131_/Q _16236_/S vssd1 vssd1 vccd1 vccd1 _16235_/A sky130_fd_sc_hd__mux2_1
X_13446_ input22/X _13340_/A _13368_/A vssd1 vssd1 vccd1 vccd1 _13446_/X sky130_fd_sc_hd__a21o_1
X_10658_ _10822_/A _10657_/X _10836_/A vssd1 vssd1 vccd1 vccd1 _10658_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12935__C1 _12897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16165_ _13023_/X _19101_/Q _16173_/S vssd1 vssd1 vccd1 vccd1 _16166_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13377_ _18607_/Q vssd1 vssd1 vccd1 vccd1 _14095_/A sky130_fd_sc_hd__clkbuf_2
X_10589_ _10822_/A _10588_/X _10674_/A vssd1 vssd1 vccd1 vccd1 _10589_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15116_ _15112_/X _15115_/X _15190_/S vssd1 vssd1 vccd1 vccd1 _15116_/X sky130_fd_sc_hd__mux2_1
X_12328_ _14885_/A _12328_/B vssd1 vssd1 vccd1 vccd1 _12329_/B sky130_fd_sc_hd__and2b_1
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16096_ _13065_/X _19071_/Q _16100_/S vssd1 vssd1 vccd1 vccd1 _16097_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17337__S _17337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19924_ _20020_/CLK _19924_/D vssd1 vssd1 vccd1 vccd1 _19924_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15646__A _15703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15047_ _15419_/A _15047_/B vssd1 vssd1 vccd1 vccd1 _15047_/X sky130_fd_sc_hd__or2_1
X_12259_ _12259_/A vssd1 vssd1 vccd1 vccd1 _12259_/X sky130_fd_sc_hd__buf_4
XFILLER_69_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16241__S _16247_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19855_ _19855_/CLK _19855_/D vssd1 vssd1 vccd1 vccd1 _19855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18806_ _19885_/CLK _18806_/D vssd1 vssd1 vccd1 vccd1 _18806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19786_ _19948_/CLK _19786_/D vssd1 vssd1 vccd1 vccd1 _19786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16998_ _16998_/A vssd1 vssd1 vccd1 vccd1 _16998_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18737_ _19909_/CLK _18737_/D vssd1 vssd1 vccd1 vccd1 _18737_/Q sky130_fd_sc_hd__dfxtp_1
X_15949_ _15964_/A _15949_/B vssd1 vssd1 vccd1 vccd1 _15949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16477__A _16545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17072__S _17072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09470_ _18990_/Q vssd1 vssd1 vccd1 vccd1 _14750_/B sky130_fd_sc_hd__buf_4
XFILLER_92_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18668_ _18734_/CLK _18668_/D vssd1 vssd1 vccd1 vccd1 _18668_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15404__A1 _18851_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17619_ _17619_/A vssd1 vssd1 vccd1 vccd1 _17628_/S sky130_fd_sc_hd__buf_4
XFILLER_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13415__B1 _12879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18599_ _20037_/CLK _18599_/D vssd1 vssd1 vccd1 vccd1 _18599_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_178_clock_A _18998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17800__S _17804_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16416__S _16424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14915__A0 _15138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09819__A _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15839__A2_N _15834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10627__S1 _10626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09554__A _10194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11052__S1 _11045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11901__B1 _15732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15990__S _15998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11295__S _11295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09806_ _09806_/A vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__buf_4
XFILLER_87_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09737_ _09737_/A vssd1 vssd1 vccd1 vccd1 _11157_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09668_ _19254_/Q _19749_/Q _09668_/S vssd1 vssd1 vccd1 vccd1 _09668_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09599_ _19523_/Q vssd1 vssd1 vccd1 vccd1 _10972_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11629_/Y _11519_/X _10445_/A _11591_/A vssd1 vssd1 vccd1 vccd1 _11631_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ _11572_/A _11561_/B vssd1 vssd1 vccd1 vccd1 _11561_/X sky130_fd_sc_hd__or2_1
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ _13289_/X _13298_/Y _13299_/Y vssd1 vssd1 vccd1 vccd1 _17058_/A sky130_fd_sc_hd__a21oi_4
XFILLER_155_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ _18851_/Q vssd1 vssd1 vccd1 vccd1 _10512_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17011__A _17094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14280_ _14280_/A _18656_/Q _14280_/C vssd1 vssd1 vccd1 vccd1 _14281_/D sky130_fd_sc_hd__and3_1
X_11492_ _19333_/Q _19604_/Q _19828_/Q _19572_/Q _10906_/S _10625_/A vssd1 vssd1 vccd1
+ vccd1 _11493_/B sky130_fd_sc_hd__mux4_1
XFILLER_11_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ _13340_/A vssd1 vssd1 vccd1 vccd1 _13231_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10443_ _10444_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__and2_1
XFILLER_170_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16850__A _16918_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input65_A io_ibus_inst[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13162_ _13161_/X _18436_/Q _13203_/S vssd1 vssd1 vccd1 vccd1 _13163_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12932__A2 _12889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _19934_/Q _19548_/Q _19998_/Q _19117_/Q _10279_/A _09745_/A vssd1 vssd1 vccd1
+ vccd1 _10375_/B sky130_fd_sc_hd__mux4_2
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12113_ _12113_/A _12113_/B vssd1 vssd1 vccd1 vccd1 _12114_/A sky130_fd_sc_hd__and2_1
XANTENNA__11994__A _11994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13093_ _13233_/A _13093_/B vssd1 vssd1 vccd1 vccd1 _13094_/A sky130_fd_sc_hd__or2_1
X_17970_ _19853_/Q _17014_/X _17976_/S vssd1 vssd1 vccd1 vccd1 _17971_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16921_ _16977_/A vssd1 vssd1 vccd1 vccd1 _16990_/S sky130_fd_sc_hd__buf_6
X_12044_ _12044_/A _14898_/A vssd1 vssd1 vccd1 vccd1 _12044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16996__S _17008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17681__A _17681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19640_ _20024_/CLK _19640_/D vssd1 vssd1 vccd1 vccd1 _19640_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_5_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_78_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16852_ _16852_/A vssd1 vssd1 vccd1 vccd1 _19389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15803_ _15813_/A _15803_/B vssd1 vssd1 vccd1 vccd1 _15804_/A sky130_fd_sc_hd__and2_1
X_19571_ _19829_/CLK _19571_/D vssd1 vssd1 vccd1 vccd1 _19571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16783_ _16783_/A vssd1 vssd1 vccd1 vccd1 _19359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13995_ _18573_/Q _13999_/C _13969_/X vssd1 vssd1 vccd1 vccd1 _13995_/Y sky130_fd_sc_hd__a21oi_1
X_15734_ _15773_/B vssd1 vssd1 vccd1 vccd1 _15734_/X sky130_fd_sc_hd__clkbuf_2
X_18522_ _18975_/CLK _18522_/D vssd1 vssd1 vccd1 vccd1 _18522_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ _12946_/A vssd1 vssd1 vccd1 vccd1 _13209_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17387__A1 _17039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11120__A1 _09881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10554__S0 _10125_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ _19747_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_1
X_15665_ _15665_/A vssd1 vssd1 vccd1 vccd1 _18910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _13070_/A vssd1 vssd1 vccd1 vccd1 _12877_/X sky130_fd_sc_hd__buf_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17620__S _17628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _17404_/A vssd1 vssd1 vccd1 vccd1 _19612_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _14629_/A _14616_/B vssd1 vssd1 vccd1 vccd1 _14617_/A sky130_fd_sc_hd__and2_1
X_18384_ _18384_/A vssd1 vssd1 vccd1 vccd1 _20022_/D sky130_fd_sc_hd__clkbuf_1
X_11828_ _19005_/Q _11828_/B vssd1 vssd1 vccd1 vccd1 _11828_/X sky130_fd_sc_hd__or2_1
XFILLER_21_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15596_ _13207_/A _18912_/Q _15600_/S vssd1 vssd1 vccd1 vccd1 _15597_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10306__S0 _10354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17173_/X _19582_/Q _17337_/S vssd1 vssd1 vccd1 vccd1 _17336_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14547_/A _15762_/A _14547_/C vssd1 vssd1 vccd1 vccd1 _14547_/X sky130_fd_sc_hd__and3_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11759_ _18696_/Q _11698_/Y _11758_/X _11712_/Y vssd1 vssd1 vccd1 vccd1 _11759_/X
+ sky130_fd_sc_hd__a211o_2
XANTENNA__16236__S _16236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10857__S1 _10856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17266_ _17266_/A vssd1 vssd1 vccd1 vccd1 _19551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09639__A _09642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14478_ _14495_/A _14478_/B _14478_/C vssd1 vssd1 vccd1 vccd1 _18725_/D sky130_fd_sc_hd__nor3_1
XFILLER_128_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16217_ _13463_/X _19125_/Q _16217_/S vssd1 vssd1 vccd1 vccd1 _16218_/A sky130_fd_sc_hd__mux2_1
X_19005_ _19025_/CLK _19005_/D vssd1 vssd1 vccd1 vccd1 _19005_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__17856__A _17867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13429_ _13449_/B _13429_/B vssd1 vssd1 vccd1 vccd1 _13429_/X sky130_fd_sc_hd__or2_1
XANTENNA__10609__S1 _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17197_ _17197_/A vssd1 vssd1 vccd1 vccd1 _19520_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12065__A _15758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16148_ _13501_/X _19095_/Q _16148_/S vssd1 vssd1 vccd1 vccd1 _16149_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11282__S1 _11065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16079_ _16135_/A vssd1 vssd1 vccd1 vccd1 _16148_/S sky130_fd_sc_hd__buf_4
XFILLER_130_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12136__B1 _12165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09374__A _18950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19907_ _19909_/CLK _19907_/D vssd1 vssd1 vccd1 vccd1 _19907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19838_ _20030_/CLK _19838_/D vssd1 vssd1 vccd1 vccd1 _19838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput1 io_dbus_rdata[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_8
X_19769_ _19995_/CLK _19769_/D vssd1 vssd1 vccd1 vccd1 _19769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12206__A2_N _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09522_ _09522_/A _11663_/A vssd1 vssd1 vccd1 vccd1 _09522_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16000__A _16057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10545__S0 _10493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09453_ _18983_/Q vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__buf_4
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09384_ _18950_/Q _11699_/A _11783_/C vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__or3b_4
XANTENNA__12611__A1 _14749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16146__S _16148_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15050__S _15127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15561__A0 _18864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18361__S _18363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15864__B2 input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10090_ _09765_/A _10089_/X _09799_/A vssd1 vssd1 vccd1 vccd1 _10090_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17705__S _17714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10223__A _10223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12800_ _12170_/X _12798_/X _12799_/Y _12234_/B vssd1 vssd1 vccd1 vccd1 _12800_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__15092__A2 _15053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13780_ _13780_/A vssd1 vssd1 vccd1 vccd1 _18492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10992_ _19136_/Q _19397_/Q _19296_/Q _19631_/Q _11048_/S _10978_/A vssd1 vssd1 vccd1
+ vccd1 _10993_/B sky130_fd_sc_hd__mux4_1
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12731_ _12729_/B _12690_/Y _12729_/C _12730_/X _12714_/B vssd1 vssd1 vccd1 vccd1
+ _12731_/X sky130_fd_sc_hd__a311o_1
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15919__A2 _15928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12976__A1_N _12967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _15384_/X _15445_/Y _15449_/Y vssd1 vssd1 vccd1 vccd1 _15451_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__18318__A0 _17688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _15487_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _12667_/A sky130_fd_sc_hd__xor2_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14411_/D vssd1 vssd1 vccd1 vccd1 _14409_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11613_ _11604_/A _11462_/A _11462_/B _11462_/C vssd1 vssd1 vccd1 vccd1 _11613_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15381_/A _15385_/A vssd1 vssd1 vccd1 vccd1 _15381_/X sky130_fd_sc_hd__or2_1
XANTENNA__10893__A _10893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ _10351_/A _18919_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _12618_/A sky130_fd_sc_hd__mux2_2
X_17120_ _17119_/X _19496_/Q _17129_/S vssd1 vssd1 vccd1 vccd1 _17121_/A sky130_fd_sc_hd__mux2_1
X_14332_ _14427_/A vssd1 vssd1 vccd1 vccd1 _14332_/X sky130_fd_sc_hd__clkbuf_2
X_11544_ _20040_/Q _19878_/Q _19287_/Q _19057_/Q _11534_/S _09660_/A vssd1 vssd1 vccd1
+ vccd1 _11545_/B sky130_fd_sc_hd__mux4_2
XANTENNA__09459__A _18971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ _17051_/A vssd1 vssd1 vccd1 vccd1 _19470_/D sky130_fd_sc_hd__clkbuf_1
X_14263_ _18655_/Q _14259_/B _14262_/Y vssd1 vssd1 vccd1 vccd1 _18655_/D sky130_fd_sc_hd__o21a_1
X_11475_ _10712_/X _11466_/X _11470_/X _11474_/X _09551_/A vssd1 vssd1 vccd1 vccd1
+ _11475_/X sky130_fd_sc_hd__a311o_2
XFILLER_109_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11169__A1 _15925_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11169__B2 _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16002_ _16002_/A vssd1 vssd1 vccd1 vccd1 _19031_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13214_ _18597_/Q _11732_/X _13211_/X _13212_/X _13213_/X vssd1 vssd1 vccd1 vccd1
+ _13627_/B sky130_fd_sc_hd__a2111o_4
X_10426_ _10027_/A _10425_/X _10376_/A vssd1 vssd1 vccd1 vccd1 _10426_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14194_ _18637_/Q _14197_/C _14193_/Y vssd1 vssd1 vccd1 vccd1 _18637_/D sky130_fd_sc_hd__o21a_1
XFILLER_152_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_126_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _13145_/A vssd1 vssd1 vccd1 vccd1 _13289_/A sky130_fd_sc_hd__buf_2
X_10357_ _10054_/A _10356_/X _10305_/A vssd1 vssd1 vccd1 vccd1 _10357_/X sky130_fd_sc_hd__a21o_1
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _17953_/A vssd1 vssd1 vccd1 vccd1 _19846_/D sky130_fd_sc_hd__clkbuf_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _13075_/Y _11845_/X _09410_/A vssd1 vssd1 vccd1 vccd1 _13076_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11016__S1 _11015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10288_ _09780_/A _10285_/Y _10287_/Y _09807_/A vssd1 vssd1 vccd1 vccd1 _10288_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17615__S _17617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16904_ _16904_/A vssd1 vssd1 vccd1 vccd1 _19413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12027_ _18520_/Q _12234_/B vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__and2_1
XFILLER_120_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17884_ _17952_/S vssd1 vssd1 vccd1 vccd1 _17893_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_78_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19623_ _19979_/CLK _19623_/D vssd1 vssd1 vccd1 vccd1 _19623_/Q sky130_fd_sc_hd__dfxtp_1
X_16835_ _16835_/A vssd1 vssd1 vccd1 vccd1 _19383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15083__A2 _15078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19554_ _19942_/CLK _19554_/D vssd1 vssd1 vccd1 vccd1 _19554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13978_ _18566_/Q _13976_/B _13977_/Y vssd1 vssd1 vccd1 vccd1 _18566_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16766_ _16834_/S vssd1 vssd1 vccd1 vccd1 _16775_/S sky130_fd_sc_hd__buf_2
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14291__B1 _14792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18505_ _19996_/CLK _18505_/D vssd1 vssd1 vccd1 vccd1 _18505_/Q sky130_fd_sc_hd__dfxtp_1
X_15717_ _18934_/Q _15740_/B vssd1 vssd1 vccd1 vccd1 _15717_/X sky130_fd_sc_hd__or2_1
X_12929_ _18583_/Q vssd1 vssd1 vccd1 vccd1 _14026_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16697_ _19321_/Q _13762_/X _16703_/S vssd1 vssd1 vccd1 vccd1 _16698_/A sky130_fd_sc_hd__mux2_1
X_19485_ _19485_/CLK _19485_/D vssd1 vssd1 vccd1 vccd1 _19485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17350__S _17352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18436_ _19633_/CLK _18436_/D vssd1 vssd1 vccd1 vccd1 _18436_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15648_ _15648_/A vssd1 vssd1 vccd1 vccd1 _18902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16474__B _16474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14594__A1 _13591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13397__A2 _13269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15579_ _15579_/A vssd1 vssd1 vccd1 vccd1 _18872_/D sky130_fd_sc_hd__clkbuf_1
X_18367_ _18367_/A vssd1 vssd1 vccd1 vccd1 _20014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10604__B1 _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17318_ _17147_/X _19574_/Q _17326_/S vssd1 vssd1 vccd1 vccd1 _17319_/A sky130_fd_sc_hd__mux2_1
X_18298_ _17659_/X _19984_/Q _18302_/S vssd1 vssd1 vccd1 vccd1 _18299_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10080__A1 _09547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17586__A _17632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17249_ _17249_/A vssd1 vssd1 vccd1 vccd1 _19543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17296__A0 _17115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12523__A _18537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13338__B _18855_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18210__A _18278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09832__A _10424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15553__B _15553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13085__A1 _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14282__B1 _14792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09505_ _09516_/A _09248_/X _09206_/Y _09272_/C vssd1 vssd1 vccd1 vccd1 _09506_/B
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11096__B1 _11095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11191__S0 _10618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _11925_/B _09436_/B _09436_/C _09436_/D vssd1 vssd1 vccd1 vccd1 _09437_/A
+ sky130_fd_sc_hd__nand4_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14585__A1 _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ _11697_/A vssd1 vssd1 vccd1 vccd1 _15773_/A sky130_fd_sc_hd__inv_2
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09298_ _18936_/Q vssd1 vssd1 vccd1 vccd1 _16846_/B sky130_fd_sc_hd__inv_4
XANTENNA__11494__S1 _10625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ _11050_/A _11259_/X _11425_/A vssd1 vssd1 vccd1 vccd1 _11260_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17287__A0 _17103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ _10211_/A vssd1 vssd1 vccd1 vccd1 _10748_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13529__A hold6/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ _19324_/Q _19595_/Q _19819_/Q _19563_/Q _10618_/A _11086_/A vssd1 vssd1 vccd1
+ vccd1 _11191_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10142_ _10473_/A vssd1 vssd1 vccd1 vccd1 _10283_/A sky130_fd_sc_hd__buf_2
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10073_ _10073_/A _10073_/B vssd1 vssd1 vccd1 vccd1 _10073_/Y sky130_fd_sc_hd__nor2_1
X_14950_ _15020_/A vssd1 vssd1 vccd1 vccd1 _15121_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__13312__A2 _13071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09742__A _10638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13901_ _18541_/Q _13900_/X _12627_/X _12630_/Y _13897_/X vssd1 vssd1 vccd1 vccd1
+ _18541_/D sky130_fd_sc_hd__o221a_1
X_14881_ _15338_/B _15385_/B _14948_/S vssd1 vssd1 vccd1 vccd1 _14881_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input28_A io_dbus_rdata[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__A2 _09405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13832_ _17068_/A vssd1 vssd1 vccd1 vccd1 _13832_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16620_ _16676_/A vssd1 vssd1 vccd1 vccd1 _16689_/S sky130_fd_sc_hd__buf_6
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16551_ _16551_/A vssd1 vssd1 vccd1 vccd1 _19256_/D sky130_fd_sc_hd__clkbuf_1
X_13763_ _18487_/Q _13762_/X _13772_/S vssd1 vssd1 vccd1 vccd1 _13764_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18266__S _18274_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10975_ _11328_/A vssd1 vssd1 vccd1 vccd1 _11409_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_44_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15502_ _15419_/X _15153_/X _15501_/X _15428_/X vssd1 vssd1 vccd1 vccd1 _15502_/X
+ sky130_fd_sc_hd__o211a_2
X_12714_ _12714_/A _12714_/B vssd1 vssd1 vccd1 vccd1 _12729_/C sky130_fd_sc_hd__nor2_2
X_19270_ _19861_/CLK _19270_/D vssd1 vssd1 vccd1 vccd1 _19270_/Q sky130_fd_sc_hd__dfxtp_1
X_16482_ _19226_/Q _13765_/X _16486_/S vssd1 vssd1 vccd1 vccd1 _16483_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_52_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ _13688_/A _13693_/C _18889_/Q vssd1 vssd1 vccd1 vccd1 _13694_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15433_ _15539_/A _15436_/A vssd1 vssd1 vccd1 vccd1 _15433_/X sky130_fd_sc_hd__or2_1
X_18221_ _18278_/S vssd1 vssd1 vccd1 vccd1 _18230_/S sky130_fd_sc_hd__buf_4
XANTENNA__13379__A2 _13120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14576__A1 _13546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12645_ _12729_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _12645_/X sky130_fd_sc_hd__xor2_4
XFILLER_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13203__S _13203_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__S1 _10057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15364_ _15458_/A vssd1 vssd1 vccd1 vccd1 _15364_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18152_ _17656_/X _19919_/Q _18158_/S vssd1 vssd1 vccd1 vccd1 _18153_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12576_ _18538_/Q _18539_/Q _12576_/C vssd1 vssd1 vccd1 vccd1 _12623_/C sky130_fd_sc_hd__and3_1
XFILLER_12_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17103_ _17640_/A vssd1 vssd1 vccd1 vccd1 _17103_/X sky130_fd_sc_hd__buf_2
X_14315_ _14315_/A _14315_/B _14325_/D vssd1 vssd1 vccd1 vccd1 _18670_/D sky130_fd_sc_hd__nor3_1
XFILLER_156_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11527_ _11644_/A _10247_/Y _11524_/Y _11643_/A _11526_/Y vssd1 vssd1 vccd1 vccd1
+ _11582_/B sky130_fd_sc_hd__a311o_1
X_18083_ _18083_/A vssd1 vssd1 vccd1 vccd1 _19896_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15525__B1 _15524_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15295_ _15243_/X _15281_/X _15294_/X _15258_/X vssd1 vssd1 vccd1 vccd1 _15295_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10128__A _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17034_ _19465_/Q _17033_/X _17040_/S vssd1 vssd1 vccd1 vccd1 _17035_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output96_A _12046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14246_ _14278_/D _14279_/C vssd1 vssd1 vccd1 vccd1 _14247_/B sky130_fd_sc_hd__and2_1
X_11458_ _11269_/X _11455_/X _11607_/B _11611_/C _11609_/A vssd1 vssd1 vccd1 vccd1
+ _11606_/B sky130_fd_sc_hd__a2111o_1
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13000__B2 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ _10502_/A _10409_/B _10409_/C vssd1 vssd1 vccd1 vccd1 _10409_/Y sky130_fd_sc_hd__nor3_1
XFILLER_125_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13439__A _13439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14177_ _18631_/Q _14180_/C _14160_/X vssd1 vssd1 vccd1 vccd1 _14177_/Y sky130_fd_sc_hd__a21oi_1
X_11389_ _19225_/Q _19720_/Q _11442_/S vssd1 vssd1 vccd1 vccd1 _11389_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12343__A _12722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14261__C _14264_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _14051_/B _13120_/X _13124_/X _13125_/X _13127_/X vssd1 vssd1 vccd1 vccd1
+ _13588_/B sky130_fd_sc_hd__a2111o_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _19526_/CLK _18985_/D vssd1 vssd1 vccd1 vccd1 _18985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _17936_/A vssd1 vssd1 vccd1 vccd1 _19838_/D sky130_fd_sc_hd__clkbuf_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _14042_/A _13120_/A _13194_/A _14468_/A vssd1 vssd1 vccd1 vccd1 _13059_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18030__A _18115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15795__A1_N _15793_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17867_ _17867_/A vssd1 vssd1 vccd1 vccd1 _17876_/S sky130_fd_sc_hd__buf_4
Xclkbuf_2_2_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_39_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19606_ _19976_/CLK _19606_/D vssd1 vssd1 vccd1 vccd1 _19606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16818_ _16818_/A vssd1 vssd1 vccd1 vccd1 _19375_/D sky130_fd_sc_hd__clkbuf_1
X_17798_ _17720_/X _19777_/Q _17804_/S vssd1 vssd1 vccd1 vccd1 _17799_/A sky130_fd_sc_hd__mux2_1
X_19537_ _20021_/CLK _19537_/D vssd1 vssd1 vccd1 vccd1 _19537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16749_ _16749_/A vssd1 vssd1 vccd1 vccd1 _16758_/S sky130_fd_sc_hd__buf_4
XANTENNA__18176__S _18180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11173__S0 _11171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19468_ _20025_/CLK _19468_/D vssd1 vssd1 vccd1 vccd1 _19468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09221_ _09435_/A _09436_/B _09434_/A vssd1 vssd1 vccd1 vccd1 _09480_/A sky130_fd_sc_hd__nand3b_2
X_18419_ _18419_/A vssd1 vssd1 vccd1 vccd1 _20038_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14567__A1 _13508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19399_ _19633_/CLK _19399_/D vssd1 vssd1 vccd1 vccd1 _19399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12578__A0 _12574_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11779__D _15760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16424__S _16424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput70 reset vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_4
XANTENNA__11228__S1 _11108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10987__S0 _11121_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09985_ _19377_/Q _19712_/Q _10254_/A vssd1 vssd1 vccd1 vccd1 _09985_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11856__A2 _11815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10760_ _10760_/A _12843_/A vssd1 vssd1 vccd1 vccd1 _10761_/B sky130_fd_sc_hd__or2_1
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12281__A2 _12556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09419_ _18825_/Q _09417_/X _11722_/A vssd1 vssd1 vccd1 vccd1 _11772_/B sky130_fd_sc_hd__a21o_1
XFILLER_73_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_clock clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__13531__B hold6/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ _19367_/Q _19702_/Q _10691_/S vssd1 vssd1 vccd1 vccd1 _10691_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12569__A0 _15962_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12430_ _15847_/A _14763_/C _12429_/Y vssd1 vssd1 vccd1 vccd1 _12514_/A sky130_fd_sc_hd__a21o_2
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12361_ _12361_/A _12361_/B vssd1 vssd1 vccd1 vccd1 _12362_/A sky130_fd_sc_hd__or2_1
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16334__S _16346_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18115__A _18115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14100_ _14146_/A _14105_/C vssd1 vssd1 vccd1 vccd1 _14100_/Y sky130_fd_sc_hd__nor2_2
XFILLER_154_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _11181_/X _11309_/Y _11311_/Y _09816_/A vssd1 vssd1 vccd1 vccd1 _11312_/X
+ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_6_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19755_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09737__A _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15080_ _15102_/A vssd1 vssd1 vccd1 vccd1 _15369_/A sky130_fd_sc_hd__clkbuf_2
X_12292_ _09467_/X _12317_/A _12260_/C _12291_/X vssd1 vssd1 vccd1 vccd1 _12292_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14031_ _18585_/Q _14028_/B _14030_/Y vssd1 vssd1 vccd1 vccd1 _18585_/D sky130_fd_sc_hd__o21a_1
X_11243_ _19325_/Q _19596_/Q _19820_/Q _19564_/Q _11158_/S _11022_/A vssd1 vssd1 vccd1
+ vccd1 _11243_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11174_ _11227_/A _11174_/B vssd1 vssd1 vccd1 vccd1 _11174_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17165__S _17177_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ _19251_/Q _19746_/Q _10125_/S vssd1 vssd1 vccd1 vccd1 _10126_/B sky130_fd_sc_hd__mux2_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15474__A _15474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18770_ _19899_/CLK _18770_/D vssd1 vssd1 vccd1 vccd1 _18770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15982_ _15982_/A _15982_/B vssd1 vssd1 vccd1 vccd1 _15982_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17721_ _17720_/X _19745_/Q _17730_/S vssd1 vssd1 vccd1 vccd1 _17722_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10056_ _19376_/Q _19711_/Q _10254_/A vssd1 vssd1 vccd1 vccd1 _10057_/B sky130_fd_sc_hd__mux2_1
X_14933_ _12641_/A _15234_/B _14933_/S vssd1 vssd1 vccd1 vccd1 _14933_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12610__B _12855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output134_A _12826_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17652_ _17652_/A vssd1 vssd1 vccd1 vccd1 _17652_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10411__A _10411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14864_ _15270_/B _15436_/B _14948_/S vssd1 vssd1 vccd1 vccd1 _14864_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17983__A1 _17033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16603_ _16603_/A vssd1 vssd1 vccd1 vccd1 _19280_/D sky130_fd_sc_hd__clkbuf_1
X_13815_ _13815_/A vssd1 vssd1 vccd1 vccd1 _18503_/D sky130_fd_sc_hd__clkbuf_1
X_14795_ _14795_/A _14795_/B vssd1 vssd1 vccd1 vccd1 _18830_/D sky130_fd_sc_hd__nor2_1
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17583_ _17583_/A vssd1 vssd1 vccd1 vccd1 _19695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19322_ _19947_/CLK _19322_/D vssd1 vssd1 vccd1 vccd1 _19322_/Q sky130_fd_sc_hd__dfxtp_1
X_16534_ _16534_/A vssd1 vssd1 vccd1 vccd1 _19249_/D sky130_fd_sc_hd__clkbuf_1
X_13746_ _18896_/Q _13746_/B vssd1 vssd1 vccd1 vccd1 _13746_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10958_ _11435_/A vssd1 vssd1 vccd1 vccd1 _11344_/A sky130_fd_sc_hd__buf_2
XFILLER_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19253_ _20006_/CLK _19253_/D vssd1 vssd1 vccd1 vccd1 _19253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16465_ _16465_/A vssd1 vssd1 vccd1 vccd1 _19219_/D sky130_fd_sc_hd__clkbuf_1
X_13677_ _13656_/X _13675_/X _13676_/Y _13660_/X _19015_/Q vssd1 vssd1 vccd1 vccd1
+ _13677_/X sky130_fd_sc_hd__a32o_2
X_10889_ _10882_/Y _10884_/Y _10886_/Y _10888_/Y _09550_/A vssd1 vssd1 vccd1 vccd1
+ _10889_/X sky130_fd_sc_hd__o221a_1
XFILLER_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12338__A _12338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18204_ _17732_/X _19943_/Q _18206_/S vssd1 vssd1 vccd1 vccd1 _18205_/A sky130_fd_sc_hd__mux2_1
X_12628_ _18780_/Q _18779_/Q _12628_/C vssd1 vssd1 vccd1 vccd1 _12679_/C sky130_fd_sc_hd__and3_1
X_15416_ _15405_/X _15414_/X _15415_/X _15048_/X _12521_/Y vssd1 vssd1 vccd1 vccd1
+ _15416_/X sky130_fd_sc_hd__a32o_1
X_19184_ _20034_/CLK _19184_/D vssd1 vssd1 vccd1 vccd1 _19184_/Q sky130_fd_sc_hd__dfxtp_1
X_16396_ _17732_/A vssd1 vssd1 vccd1 vccd1 _16396_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15347_ _15199_/X _15202_/X _15347_/S vssd1 vssd1 vccd1 vccd1 _15347_/X sky130_fd_sc_hd__mux2_1
X_18135_ _18135_/A vssd1 vssd1 vccd1 vccd1 _19912_/D sky130_fd_sc_hd__clkbuf_1
X_12559_ _12338_/X _12555_/X _12558_/Y vssd1 vssd1 vccd1 vccd1 _12559_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_117_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_opt_7_0_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15278_ _15457_/A vssd1 vssd1 vccd1 vccd1 _15278_/X sky130_fd_sc_hd__clkbuf_2
X_18066_ _18066_/A vssd1 vssd1 vccd1 vccd1 _19891_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11896__B _11896_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14229_ _18646_/Q _14242_/C vssd1 vssd1 vccd1 vccd1 _14231_/B sky130_fd_sc_hd__or2_1
XANTENNA__14721__A1 _13677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17017_ _17017_/A vssd1 vssd1 vccd1 vccd1 _17017_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11535__A1 _09639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15277__A2 _09433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ _19387_/Q vssd1 vssd1 vccd1 vccd1 _11181_/A sky130_fd_sc_hd__inv_2
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ _18997_/CLK _18968_/D vssd1 vssd1 vccd1 vccd1 _18968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _17919_/A vssd1 vssd1 vccd1 vccd1 _19830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18899_ _18997_/CLK _18899_/D vssd1 vssd1 vccd1 vccd1 _18899_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10197__S1 _10182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__S0 _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11146__S0 _11023_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14447__B _14447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10274__B2 _18856_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09204_ _11956_/A vssd1 vssd1 vccd1 vccd1 _14811_/A sky130_fd_sc_hd__inv_2
XFILLER_50_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13748__C1 _11730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16154__S _16162_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14463__A _14472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10991__A _11049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12971__B1 _11796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14712__A1 _11748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10734__C1 _09874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09968_ _19938_/Q _19552_/Q _20002_/Q _19121_/Q _09967_/X _09612_/A vssd1 vssd1 vccd1
+ vccd1 _09969_/B sky130_fd_sc_hd__mux4_1
XFILLER_103_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13279__A1 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__A _12713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09899_ _09833_/X _09898_/X _09942_/A vssd1 vssd1 vccd1 vccd1 _09899_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _12078_/A vssd1 vssd1 vccd1 vccd1 _14931_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _13879_/A _18713_/Q _14534_/S vssd1 vssd1 vccd1 vccd1 _11861_/X sky130_fd_sc_hd__or3_1
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _11833_/D _13599_/Y _13623_/S vssd1 vssd1 vccd1 vccd1 _13600_/X sky130_fd_sc_hd__mux2_1
X_10812_ _10211_/A _10809_/X _10811_/X vssd1 vssd1 vccd1 vccd1 _10812_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13542__A _18999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17014__A _17014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14580_ _14648_/A vssd1 vssd1 vccd1 vccd1 _14595_/A sky130_fd_sc_hd__buf_2
X_11792_ _18649_/Q _11815_/A _12876_/A _18553_/Q vssd1 vssd1 vccd1 vccd1 _11796_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13531_ _13531_/A hold6/A vssd1 vssd1 vccd1 vccd1 _13531_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10743_ _10748_/A _10743_/B vssd1 vssd1 vccd1 vccd1 _10743_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12158__A _18104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16250_ _13137_/X _19138_/Q _16258_/S vssd1 vssd1 vccd1 vccd1 _16251_/A sky130_fd_sc_hd__mux2_1
X_13462_ _17087_/A vssd1 vssd1 vccd1 vccd1 _17729_/A sky130_fd_sc_hd__clkbuf_2
X_10674_ _10674_/A _10674_/B vssd1 vssd1 vccd1 vccd1 _10674_/X sky130_fd_sc_hd__or2_1
XFILLER_139_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15201_ _12031_/B _15201_/B vssd1 vssd1 vccd1 vccd1 _15201_/X sky130_fd_sc_hd__and2b_1
X_12413_ _12438_/A _12413_/B vssd1 vssd1 vccd1 vccd1 _12413_/Y sky130_fd_sc_hd__xnor2_4
X_16181_ _16181_/A vssd1 vssd1 vccd1 vccd1 _19108_/D sky130_fd_sc_hd__clkbuf_1
X_13393_ _13427_/C _13393_/B vssd1 vssd1 vccd1 vccd1 _13393_/X sky130_fd_sc_hd__or2_1
XFILLER_154_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_154_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _18789_/CLK sky130_fd_sc_hd__clkbuf_16
X_15132_ _14917_/X _14876_/X _15132_/S vssd1 vssd1 vccd1 vccd1 _15132_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12344_ _12344_/A vssd1 vssd1 vccd1 vccd1 _12344_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16999__S _17008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19940_ _19940_/CLK _19940_/D vssd1 vssd1 vccd1 vccd1 _19940_/Q sky130_fd_sc_hd__dfxtp_1
X_15063_ _14874_/X _14911_/X _15117_/S vssd1 vssd1 vccd1 vccd1 _15063_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14703__A1 _13612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12275_ _12275_/A vssd1 vssd1 vccd1 vccd1 _12814_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14014_ _14046_/A _14016_/B vssd1 vssd1 vccd1 vccd1 _14014_/Y sky130_fd_sc_hd__nor2_1
XFILLER_136_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13911__C1 _14792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11226_ _18429_/Q _19458_/Q _19495_/Q _19069_/Q _11293_/A _09737_/A vssd1 vssd1 vccd1
+ vccd1 _11227_/B sky130_fd_sc_hd__mux4_1
X_19871_ _20033_/CLK _19871_/D vssd1 vssd1 vccd1 vccd1 _19871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_169_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _18526_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold6_A hold6/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18822_ _18960_/CLK _18822_/D vssd1 vssd1 vccd1 vccd1 _18822_/Q sky130_fd_sc_hd__dfxtp_1
X_11157_ _11157_/A _11157_/B vssd1 vssd1 vccd1 vccd1 _11157_/X sky130_fd_sc_hd__and2_1
XFILLER_96_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10108_ _10129_/S vssd1 vssd1 vccd1 vccd1 _10314_/S sky130_fd_sc_hd__buf_4
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18753_ _18956_/CLK _18753_/D vssd1 vssd1 vccd1 vccd1 _18753_/Q sky130_fd_sc_hd__dfxtp_2
X_15965_ _19016_/Q _15954_/X _15955_/X _15964_/Y vssd1 vssd1 vccd1 vccd1 _19016_/D
+ sky130_fd_sc_hd__a22o_1
X_11088_ _11088_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11088_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11376__S0 _11328_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17704_ _17704_/A vssd1 vssd1 vccd1 vccd1 _17704_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__15932__A _19003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11237__A _11237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ _10294_/A _10034_/X _10036_/Y _10038_/Y vssd1 vssd1 vccd1 vccd1 _10039_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_14916_ _14913_/X _14915_/X _14916_/S vssd1 vssd1 vccd1 vccd1 _14916_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18684_ _19882_/CLK _18684_/D vssd1 vssd1 vccd1 vccd1 _18684_/Q sky130_fd_sc_hd__dfxtp_1
X_15896_ _12316_/A _15842_/X _15843_/X input58/X vssd1 vssd1 vccd1 vccd1 _15897_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17635_ _17635_/A _17635_/B vssd1 vssd1 vccd1 vccd1 _17717_/A sky130_fd_sc_hd__or2_4
X_14847_ _11971_/B _15142_/A _15151_/A _12871_/B vssd1 vssd1 vccd1 vccd1 _14847_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14548__A _14548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16239__S _16247_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17566_ _17566_/A vssd1 vssd1 vccd1 vccd1 _19687_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_107_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19971_/CLK sky130_fd_sc_hd__clkbuf_16
X_14778_ _14778_/A vssd1 vssd1 vccd1 vccd1 _14789_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19305_ _19993_/CLK _19305_/D vssd1 vssd1 vccd1 vccd1 _19305_/Q sky130_fd_sc_hd__dfxtp_1
X_16517_ _19242_/Q _13816_/X _16519_/S vssd1 vssd1 vccd1 vccd1 _16518_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13729_ _18482_/Q _13526_/A _13724_/Y _13728_/X vssd1 vssd1 vccd1 vccd1 _18482_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17497_ _17497_/A vssd1 vssd1 vccd1 vccd1 _19654_/D sky130_fd_sc_hd__clkbuf_1
X_19236_ _19827_/CLK _19236_/D vssd1 vssd1 vccd1 vccd1 _19236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16448_ _16459_/A vssd1 vssd1 vccd1 vccd1 _16457_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__15195__B2 _12150_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19167_ _20016_/CLK _19167_/D vssd1 vssd1 vccd1 vccd1 _19167_/Q sky130_fd_sc_hd__dfxtp_1
X_16379_ _16379_/A vssd1 vssd1 vccd1 vccd1 _19184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18133__A1 _18864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11756__A1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__A _15758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__S0 _11171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18118_ _18859_/Q _13710_/X _18118_/S vssd1 vssd1 vccd1 vccd1 _18118_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19098_ _19979_/CLK _19098_/D vssd1 vssd1 vccd1 vccd1 _19098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18049_ _18049_/A vssd1 vssd1 vccd1 vccd1 _19886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_174_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _09822_/A vssd1 vssd1 vccd1 vccd1 _09823_/A sky130_fd_sc_hd__clkbuf_4
X_20011_ _20012_/CLK _20011_/D vssd1 vssd1 vccd1 vccd1 _20011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10750__S _10750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13627__A _19009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09753_ _11111_/A vssd1 vssd1 vccd1 vccd1 _11311_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15842__A _15875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10051__A _10587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ _10719_/A vssd1 vssd1 vccd1 vccd1 _09685_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10986__A _11212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14458__A _15715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10590__S1 _09607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12236__A2 _12835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_99_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09986__S _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_71_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19975_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14933__A1 _15234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18124__A1 _13727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10390_ _10380_/A _10385_/X _10387_/X _10389_/X vssd1 vssd1 vccd1 vccd1 _10390_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_163_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_86_clock clkbuf_opt_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19996_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17708__S _17714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10226__A _10388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ _12060_/A _12060_/B vssd1 vssd1 vccd1 vccd1 _12060_/X sky130_fd_sc_hd__or2_1
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11011_ _18841_/Q vssd1 vssd1 vccd1 vccd1 _11011_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_89_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11358__S0 _11356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _18946_/Q _15760_/B vssd1 vssd1 vccd1 vccd1 _15750_/X sky130_fd_sc_hd__or2_1
X_12962_ _17001_/A vssd1 vssd1 vccd1 vccd1 _17643_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11132__C1 _11058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input10_A io_dbus_rdata[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18060__A0 _18842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10486__A1 _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _15633_/C _12153_/B _12153_/C vssd1 vssd1 vccd1 vccd1 _12275_/A sky130_fd_sc_hd__and3_1
X_14701_ _18802_/Q _11860_/D _14705_/S vssd1 vssd1 vccd1 vccd1 _14702_/A sky130_fd_sc_hd__mux2_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19957_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15471__B _15474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _15681_/A vssd1 vssd1 vccd1 vccd1 _18917_/D sky130_fd_sc_hd__clkbuf_1
X_12893_ _19488_/Q vssd1 vssd1 vccd1 vccd1 _13215_/S sky130_fd_sc_hd__buf_2
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _19620_/Q _17087_/X _17420_/S vssd1 vssd1 vccd1 vccd1 _17421_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _18769_/Q vssd1 vssd1 vccd1 vccd1 _12349_/A sky130_fd_sc_hd__clkbuf_2
X_14632_ _18778_/Q _13677_/X _14632_/S vssd1 vssd1 vccd1 vccd1 _14633_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _17351_/A vssd1 vssd1 vccd1 vccd1 _19589_/D sky130_fd_sc_hd__clkbuf_1
X_14563_ _14601_/A vssd1 vssd1 vccd1 vccd1 _14581_/S sky130_fd_sc_hd__buf_2
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _13082_/A vssd1 vssd1 vccd1 vccd1 _13194_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18274__S _18274_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09896__S _09903_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16302_ _16297_/X _19160_/Q _16314_/S vssd1 vssd1 vccd1 vccd1 _16303_/A sky130_fd_sc_hd__mux2_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _19238_/Q _19733_/Q _10821_/S vssd1 vssd1 vccd1 vccd1 _10726_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19796_/CLK sky130_fd_sc_hd__clkbuf_16
X_13514_ _18456_/Q _13509_/Y _13514_/S vssd1 vssd1 vccd1 vccd1 _13515_/A sky130_fd_sc_hd__mux2_1
X_17282_ _17426_/A _17882_/B vssd1 vssd1 vccd1 vccd1 _17339_/A sky130_fd_sc_hd__or2_4
X_14494_ _14493_/B _14493_/C _18731_/Q vssd1 vssd1 vccd1 vccd1 _14495_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__11450__A3 _11449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_110_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19021_ _19973_/CLK _19021_/D vssd1 vssd1 vccd1 vccd1 _19021_/Q sky130_fd_sc_hd__dfxtp_1
X_13445_ _13445_/A vssd1 vssd1 vccd1 vccd1 _18452_/D sky130_fd_sc_hd__clkbuf_1
X_16233_ _16233_/A vssd1 vssd1 vccd1 vccd1 _19130_/D sky130_fd_sc_hd__clkbuf_1
X_10657_ _19239_/Q _19734_/Q _10657_/S vssd1 vssd1 vccd1 vccd1 _10657_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16164_ _16221_/S vssd1 vssd1 vccd1 vccd1 _16173_/S sky130_fd_sc_hd__clkbuf_4
X_13376_ _18671_/Q _12889_/X _11852_/X _18639_/Q vssd1 vssd1 vccd1 vccd1 _13376_/X
+ sky130_fd_sc_hd__a22o_2
X_10588_ _19240_/Q _19735_/Q _10657_/S vssd1 vssd1 vccd1 vccd1 _10588_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09800__B1 _09809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15115_ _15113_/X _15114_/X _15189_/S vssd1 vssd1 vccd1 vccd1 _15115_/X sky130_fd_sc_hd__mux2_1
X_12327_ _12328_/B _14885_/A vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__and2b_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15927__A _15954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16095_ _16095_/A vssd1 vssd1 vccd1 vccd1 _19070_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16522__S _16530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19923_ _20021_/CLK _19923_/D vssd1 vssd1 vccd1 vccd1 _19923_/Q sky130_fd_sc_hd__dfxtp_1
X_15046_ _15027_/X _15044_/X _15247_/A vssd1 vssd1 vccd1 vccd1 _15047_/B sky130_fd_sc_hd__mux2_1
XFILLER_170_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12258_ _12258_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12259_/A sky130_fd_sc_hd__and2_1
XANTENNA__17626__A0 _17189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11209_ _19324_/Q _19595_/Q _19819_/Q _19563_/Q _11273_/A _11208_/X vssd1 vssd1 vccd1
+ vccd1 _11209_/X sky130_fd_sc_hd__mux4_1
X_19854_ _19949_/CLK _19854_/D vssd1 vssd1 vccd1 vccd1 _19854_/Q sky130_fd_sc_hd__dfxtp_1
X_12189_ _12275_/A vssd1 vssd1 vccd1 vccd1 _12479_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18805_ _19896_/CLK _18805_/D vssd1 vssd1 vccd1 vccd1 _18805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19785_ _19947_/CLK _19785_/D vssd1 vssd1 vccd1 vccd1 _19785_/Q sky130_fd_sc_hd__dfxtp_1
X_16997_ _16997_/A vssd1 vssd1 vccd1 vccd1 _19453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18736_ _19909_/CLK _18736_/D vssd1 vssd1 vccd1 vccd1 _18736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15948_ _19009_/Q _15921_/X _15947_/X vssd1 vssd1 vccd1 vccd1 _19009_/D sky130_fd_sc_hd__a21o_1
XANTENNA__13663__A1 _18473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__A1 _10380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__A _09660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__A2 _18939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18667_ _18734_/CLK _18667_/D vssd1 vssd1 vccd1 vccd1 _18667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15879_ _15879_/A vssd1 vssd1 vccd1 vccd1 _15879_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14278__A _18653_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17618_ _17618_/A vssd1 vssd1 vccd1 vccd1 _19711_/D sky130_fd_sc_hd__clkbuf_1
X_18598_ _20037_/CLK _18598_/D vssd1 vssd1 vccd1 vccd1 _18598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10229__A1 _09798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17549_ _17549_/A vssd1 vssd1 vccd1 vccd1 _19680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13910__A _13910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19219_ _20036_/CLK _19219_/D vssd1 vssd1 vccd1 vccd1 _19219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14915__A1 _12713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11901__A1 _18711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input2_A io_dbus_rdata[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _09805_/A vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__buf_2
XFILLER_140_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18359__S _18363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17263__S _17265_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09736_ _11172_/A vssd1 vssd1 vccd1 vccd1 _09737_/A sky130_fd_sc_hd__buf_2
XFILLER_83_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09667_ _10355_/A vssd1 vssd1 vccd1 vccd1 _11533_/A sky130_fd_sc_hd__buf_4
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09598_ _09668_/S vssd1 vssd1 vccd1 vccd1 _09598_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16607__S _16613_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11560_ _20040_/Q _19878_/Q _19287_/Q _19057_/Q _11566_/S _11554_/A vssd1 vssd1 vccd1
+ vccd1 _11561_/B sky130_fd_sc_hd__mux4_1
XFILLER_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10511_ _10504_/Y _10506_/Y _10508_/Y _10510_/Y _10668_/A vssd1 vssd1 vccd1 vccd1
+ _10511_/X sky130_fd_sc_hd__o221a_1
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10655__S _10655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ _11487_/X _11489_/X _11490_/X _10211_/A _09776_/A vssd1 vssd1 vccd1 vccd1
+ _11491_/X sky130_fd_sc_hd__o221a_1
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11340__A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ _13268_/A _13256_/C _13225_/Y _13229_/X vssd1 vssd1 vccd1 vccd1 _13230_/X
+ sky130_fd_sc_hd__o31a_1
X_10442_ _09884_/A _10432_/X _10441_/X _09913_/A _10419_/Y vssd1 vssd1 vccd1 vccd1
+ _12851_/B sky130_fd_sc_hd__o32a_4
XFILLER_136_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _17675_/A vssd1 vssd1 vccd1 vccd1 _13161_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10373_ _09849_/X _10363_/X _10372_/X _09540_/A _18854_/Q vssd1 vssd1 vccd1 vccd1
+ _15962_/C sky130_fd_sc_hd__a32o_4
XFILLER_152_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12112_ _13508_/A _12098_/X _12099_/X _12111_/Y _12402_/B vssd1 vssd1 vccd1 vccd1
+ _12113_/B sky130_fd_sc_hd__a311o_1
XFILLER_151_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input58_A io_ibus_inst[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _13092_/A _14789_/A _18828_/Q input30/X vssd1 vssd1 vccd1 vccd1 _13093_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11486__S _11486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16920_ _17738_/A _17635_/B vssd1 vssd1 vccd1 vccd1 _16977_/A sky130_fd_sc_hd__or2_4
X_12043_ _12043_/A _12043_/B vssd1 vssd1 vccd1 vccd1 _12046_/A sky130_fd_sc_hd__nor2_2
XFILLER_132_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16851_ _16297_/X _19389_/Q _16859_/S vssd1 vssd1 vccd1 vccd1 _16852_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15802_ _09481_/A _11860_/A _15798_/X input59/X vssd1 vssd1 vccd1 vccd1 _15803_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15482__A _15482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19570_ _19732_/CLK _19570_/D vssd1 vssd1 vccd1 vccd1 _19570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16782_ _16323_/X _19359_/Q _16786_/S vssd1 vssd1 vccd1 vccd1 _16783_/A sky130_fd_sc_hd__mux2_1
X_13994_ _18572_/Q _13992_/B _13993_/Y vssd1 vssd1 vccd1 vccd1 _18572_/D sky130_fd_sc_hd__o21a_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18521_ _18975_/CLK _18521_/D vssd1 vssd1 vccd1 vccd1 _18521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _18971_/Q _15720_/X _15732_/Y _15730_/X vssd1 vssd1 vccd1 vccd1 _18939_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _18680_/Q vssd1 vssd1 vccd1 vccd1 _14350_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14098__A _14245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11515__A _15952_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _19587_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_122_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15664_ _18910_/Q _12368_/A _15666_/S vssd1 vssd1 vccd1 vccd1 _15665_/A sky130_fd_sc_hd__mux2_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _12876_/A vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__buf_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _19612_/Q _17062_/X _17409_/S vssd1 vssd1 vccd1 vccd1 _17404_/A sky130_fd_sc_hd__mux2_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _12452_/A _11724_/X _14615_/S vssd1 vssd1 vccd1 vccd1 _14616_/B sky130_fd_sc_hd__mux2_1
XFILLER_92_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18383_ _17678_/X _20022_/Q _18385_/S vssd1 vssd1 vccd1 vccd1 _18384_/A sky130_fd_sc_hd__mux2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _14280_/A _11815_/X _11823_/X _11825_/X _11826_/X vssd1 vssd1 vccd1 vccd1
+ _11828_/B sky130_fd_sc_hd__a2111o_2
XANTENNA__16517__S _16519_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _15595_/A vssd1 vssd1 vccd1 vccd1 _18879_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10306__S1 _10182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11503__S0 _11488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17334_/A vssd1 vssd1 vccd1 vccd1 _19581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _18747_/Q _11677_/B _14555_/B _12508_/A _11757_/X vssd1 vssd1 vccd1 vccd1
+ _11758_/X sky130_fd_sc_hd__a221o_1
X_14546_ _14546_/A vssd1 vssd1 vccd1 vccd1 _14547_/C sky130_fd_sc_hd__inv_2
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ _10709_/A vssd1 vssd1 vccd1 vccd1 _10710_/A sky130_fd_sc_hd__buf_2
X_17265_ _17176_/X _19551_/Q _17265_/S vssd1 vssd1 vccd1 vccd1 _17266_/A sky130_fd_sc_hd__mux2_1
X_11689_ _11734_/A vssd1 vssd1 vccd1 vccd1 _13081_/A sky130_fd_sc_hd__buf_2
X_14477_ _14476_/B _14476_/C _18725_/Q vssd1 vssd1 vccd1 vccd1 _14478_/C sky130_fd_sc_hd__a21oi_1
X_19004_ _19025_/CLK _19004_/D vssd1 vssd1 vccd1 vccd1 _19004_/Q sky130_fd_sc_hd__dfxtp_1
X_16216_ _16216_/A vssd1 vssd1 vccd1 vccd1 _19124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15570__A1 _18900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13428_ _13714_/B _13427_/C _18893_/Q vssd1 vssd1 vccd1 vccd1 _13429_/B sky130_fd_sc_hd__a21oi_1
XFILLER_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17196_ _17195_/X _19520_/Q _17199_/S vssd1 vssd1 vccd1 vccd1 _17197_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17348__S _17348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16147_ _16147_/A vssd1 vssd1 vccd1 vccd1 _19094_/D sky130_fd_sc_hd__clkbuf_1
X_13359_ _13390_/C _13359_/B _13359_/C vssd1 vssd1 vccd1 vccd1 _13359_/X sky130_fd_sc_hd__and3b_1
XANTENNA__15657__A _15703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16252__S _16258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09655__A _09655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16078_ _16993_/A _17738_/B vssd1 vssd1 vccd1 vccd1 _16135_/A sky130_fd_sc_hd__or2_4
XFILLER_130_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15029_ _15029_/A vssd1 vssd1 vccd1 vccd1 _15039_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_69_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19906_ _19910_/CLK _19906_/D vssd1 vssd1 vccd1 vccd1 _19906_/Q sky130_fd_sc_hd__dfxtp_1
X_19837_ _19997_/CLK _19837_/D vssd1 vssd1 vccd1 vccd1 _19837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16488__A _16545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15392__A _15397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 io_dbus_rdata[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_6
X_19768_ _19993_/CLK _19768_/D vssd1 vssd1 vccd1 vccd1 _19768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09521_ _09521_/A vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__clkbuf_4
X_18719_ _18719_/CLK _18719_/D vssd1 vssd1 vccd1 vccd1 _18719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19699_ _19796_/CLK _19699_/D vssd1 vssd1 vccd1 vccd1 _19699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10545__S1 _10587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13116__S _13116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11425__A _11425_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ _18984_/Q vssd1 vssd1 vccd1 vccd1 _14749_/A sky130_fd_sc_hd__buf_4
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09383_ _18952_/Q _18951_/Q vssd1 vssd1 vccd1 vccd1 _11783_/C sky130_fd_sc_hd__nor2_1
XANTENNA__16427__S _16435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15561__A1 _15560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12406__D _15338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16162__S _16162_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10481__S0 _10388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15864__A2 _15856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10504__A _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09719_ _10960_/A vssd1 vssd1 vccd1 vccd1 _11348_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_16_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10991_ _11049_/S vssd1 vssd1 vccd1 vccd1 _11048_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_16_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17721__S _17730_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15870__A2_N _15834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _12713_/A _15509_/B _12689_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _12730_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15919__A3 _12118_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10861__A1 _09830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12613_/A _12612_/A _15474_/A _12632_/A vssd1 vssd1 vccd1 vccd1 _12662_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16337__S _16346_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14400_ _18696_/Q _18695_/Q _18694_/Q _14400_/D vssd1 vssd1 vccd1 vccd1 _14411_/D
+ sky130_fd_sc_hd__and4_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11462_/C _11606_/Y _11608_/Y _11611_/X vssd1 vssd1 vccd1 vccd1 _11614_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_169_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12687_/A vssd1 vssd1 vccd1 vccd1 _12805_/S sky130_fd_sc_hd__clkbuf_4
X_15380_ _15385_/A _15385_/B vssd1 vssd1 vccd1 vccd1 _15380_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11543_ _11543_/A _11543_/B vssd1 vssd1 vccd1 vccd1 _11543_/Y sky130_fd_sc_hd__nor2_1
X_14331_ _18674_/Q _14327_/X _14330_/Y vssd1 vssd1 vccd1 vccd1 _18674_/D sky130_fd_sc_hd__o21a_1
XFILLER_129_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09459__B hold2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16861__A _16918_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17050_ _19470_/Q _17049_/X _17056_/S vssd1 vssd1 vccd1 vccd1 _17051_/A sky130_fd_sc_hd__mux2_1
X_14262_ _14265_/A _14262_/B vssd1 vssd1 vccd1 vccd1 _14262_/Y sky130_fd_sc_hd__nor2_1
X_11474_ _11481_/A _11471_/X _11473_/X _10719_/X vssd1 vssd1 vccd1 vccd1 _11474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16001_ _13023_/X _19031_/Q _16009_/S vssd1 vssd1 vccd1 vccd1 _16002_/A sky130_fd_sc_hd__mux2_1
X_13213_ _18565_/Q _12876_/A _11855_/B _18729_/Q vssd1 vssd1 vccd1 vccd1 _13213_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17168__S _17177_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10425_ _19372_/Q _19707_/Q _10470_/S vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14193_ _18637_/Q _14197_/C _14160_/X vssd1 vssd1 vccd1 vccd1 _14193_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14381__A _18690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13144_ _18844_/Q _11828_/B _13349_/S vssd1 vssd1 vccd1 vccd1 _13144_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10356_ _19373_/Q _19708_/Q _10356_/S vssd1 vssd1 vccd1 vccd1 _10356_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output164_A _12028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13315__B1 _13312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17952_ _19846_/Q _17093_/X _17952_/S vssd1 vssd1 vccd1 vccd1 _17953_/A sky130_fd_sc_hd__mux2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _19889_/Q vssd1 vssd1 vccd1 vccd1 _13075_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16800__S _16808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10287_ _10290_/A _10287_/B vssd1 vssd1 vccd1 vccd1 _10287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16903_ _16377_/X _19413_/Q _16903_/S vssd1 vssd1 vccd1 vccd1 _16904_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12026_ _12402_/B vssd1 vssd1 vccd1 vccd1 _12234_/B sky130_fd_sc_hd__buf_2
XANTENNA__10224__S0 _10166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17883_ _17939_/A vssd1 vssd1 vccd1 vccd1 _17952_/S sky130_fd_sc_hd__buf_6
XFILLER_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19622_ _19622_/CLK _19622_/D vssd1 vssd1 vccd1 vccd1 _19622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16834_ _16399_/X _19383_/Q _16834_/S vssd1 vssd1 vccd1 vccd1 _16835_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19553_ _19971_/CLK _19553_/D vssd1 vssd1 vccd1 vccd1 _19553_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09917__S0 _09920_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16765_ _16821_/A vssd1 vssd1 vccd1 vccd1 _16834_/S sky130_fd_sc_hd__buf_6
XFILLER_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13977_ _14010_/A _13982_/C vssd1 vssd1 vccd1 vccd1 _13977_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18504_ _19995_/CLK _18504_/D vssd1 vssd1 vccd1 vccd1 _18504_/Q sky130_fd_sc_hd__dfxtp_1
X_15716_ _09436_/C _14803_/X _15715_/X _15738_/B vssd1 vssd1 vccd1 vccd1 _18933_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15940__A _15940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19484_ _19846_/CLK _19484_/D vssd1 vssd1 vccd1 vccd1 _19484_/Q sky130_fd_sc_hd__dfxtp_1
X_12928_ _19060_/Q _12878_/X _12879_/X _18758_/Q _12927_/X vssd1 vssd1 vccd1 vccd1
+ _12928_/X sky130_fd_sc_hd__a221o_2
X_16696_ _16696_/A vssd1 vssd1 vccd1 vccd1 _19320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18435_ _19636_/CLK _18435_/D vssd1 vssd1 vccd1 vccd1 _18435_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15647_ _18902_/Q _18523_/Q _15655_/S vssd1 vssd1 vccd1 vccd1 _15648_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16247__S _16247_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12859_ _12859_/A vssd1 vssd1 vccd1 vccd1 _12866_/A sky130_fd_sc_hd__buf_2
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18366_ _17652_/X _20014_/Q _18374_/S vssd1 vssd1 vccd1 vccd1 _18367_/A sky130_fd_sc_hd__mux2_1
X_15578_ _18872_/Q _18904_/Q _15578_/S vssd1 vssd1 vccd1 vccd1 _15579_/A sky130_fd_sc_hd__mux2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17317_ _17339_/A vssd1 vssd1 vccd1 vccd1 _17326_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__17867__A _17867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14529_ _14529_/A _14529_/B vssd1 vssd1 vccd1 vccd1 _14529_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18297_ _18297_/A vssd1 vssd1 vccd1 vccd1 _19983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17248_ _17151_/X _19543_/Q _17254_/S vssd1 vssd1 vccd1 vccd1 _17249_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10080__A2 _10067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17179_ _17716_/A vssd1 vssd1 vccd1 vccd1 _17179_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12804__A _15982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10463__S0 _10314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13619__B _13619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17806__S _17808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16710__S _16714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16011__A _16057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09504_ _11948_/A _11956_/B _09504_/C vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__and3b_1
XFILLER_37_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09435_ _09435_/A vssd1 vssd1 vccd1 vccd1 _09436_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__11191__S1 _11086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ _18955_/Q vssd1 vssd1 vccd1 vccd1 _11697_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15782__A1 _12260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15996__S _15998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18372__S _18374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ _18977_/Q _09322_/A _09294_/X _09295_/X _09296_/X vssd1 vssd1 vccd1 vccd1
+ _09542_/B sky130_fd_sc_hd__a2111o_1
XFILLER_166_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10210_ _10210_/A _10210_/B vssd1 vssd1 vccd1 vccd1 _10210_/Y sky130_fd_sc_hd__nand2_1
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10454__S0 _09995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__B _13529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ _19132_/Q _19393_/Q _19292_/Q _19627_/Q _11156_/S _11108_/X vssd1 vssd1 vccd1
+ vccd1 _11190_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ _10573_/S vssd1 vssd1 vccd1 vccd1 _10141_/X sky130_fd_sc_hd__buf_4
XFILLER_161_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_clock clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_153_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10072_ _19216_/Q _19807_/Q _19969_/Q _19184_/Q _09918_/S _10057_/A vssd1 vssd1 vccd1
+ vccd1 _10073_/B sky130_fd_sc_hd__mux4_1
XFILLER_43_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13900_ _13900_/A vssd1 vssd1 vccd1 vccd1 _13900_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17017__A _17017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14880_ _14880_/A vssd1 vssd1 vccd1 vccd1 _15385_/B sky130_fd_sc_hd__clkbuf_2
X_13831_ _13831_/A vssd1 vssd1 vccd1 vccd1 _18508_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13076__A2 _11845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10509__S1 _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17451__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15760__A _15760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11065__A _11073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16550_ _19256_/Q _13754_/X _16558_/S vssd1 vssd1 vccd1 vccd1 _16551_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10974_ _19522_/Q vssd1 vssd1 vccd1 vccd1 _11328_/A sky130_fd_sc_hd__clkbuf_2
X_13762_ _16998_/A vssd1 vssd1 vccd1 vccd1 _13762_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15501_ _14977_/X _15172_/B _15500_/X _15400_/X vssd1 vssd1 vccd1 vccd1 _15501_/X
+ sky130_fd_sc_hd__a211o_1
X_12713_ _12713_/A _12713_/B vssd1 vssd1 vccd1 vccd1 _12714_/B sky130_fd_sc_hd__and2_1
X_16481_ _16481_/A vssd1 vssd1 vccd1 vccd1 _19225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13693_ _18888_/Q _18889_/Q _13693_/C vssd1 vssd1 vccd1 vccd1 _13699_/B sky130_fd_sc_hd__or3_2
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18220_ _18220_/A vssd1 vssd1 vccd1 vccd1 _19949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15432_ _15436_/A _15436_/B vssd1 vssd1 vccd1 vccd1 _15432_/Y sky130_fd_sc_hd__nand2_1
X_12644_ _12598_/A _12598_/B _12621_/A _12643_/Y vssd1 vssd1 vccd1 vccd1 _12645_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18151_ _18151_/A vssd1 vssd1 vccd1 vccd1 _19918_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12575_ _12554_/A _12576_/C _18539_/Q vssd1 vssd1 vccd1 vccd1 _12577_/A sky130_fd_sc_hd__a21oi_1
X_15363_ _15457_/A vssd1 vssd1 vccd1 vccd1 _15363_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10409__A _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17102_ _17102_/A vssd1 vssd1 vccd1 vccd1 _19490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14314_ _18670_/Q _14316_/B _14314_/C vssd1 vssd1 vccd1 vccd1 _14325_/D sky130_fd_sc_hd__and3_1
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11526_ _15978_/C _12863_/B vssd1 vssd1 vccd1 vccd1 _11526_/Y sky130_fd_sc_hd__nor2_1
X_18082_ _18080_/X _19896_/Q _18095_/S vssd1 vssd1 vccd1 vccd1 _18083_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15525__A1 _12743_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15294_ _15282_/X _15283_/X _15293_/X _15238_/X vssd1 vssd1 vccd1 vccd1 _15294_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12339__A1 _12340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14823__B _15004_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17033_ _17033_/A vssd1 vssd1 vccd1 vccd1 _17033_/X sky130_fd_sc_hd__clkbuf_2
X_11457_ _15923_/C _12830_/B vssd1 vssd1 vccd1 vccd1 _11611_/C sky130_fd_sc_hd__nor2_1
X_14245_ _14245_/A vssd1 vssd1 vccd1 vccd1 _14265_/A sky130_fd_sc_hd__buf_2
XFILLER_171_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10408_ _10415_/A _10405_/X _10407_/X _10192_/X vssd1 vssd1 vccd1 vccd1 _10409_/C
+ sky130_fd_sc_hd__o211a_1
X_14176_ _18630_/Q _14174_/B _14175_/Y vssd1 vssd1 vccd1 vccd1 _18630_/D sky130_fd_sc_hd__o21a_1
XANTENNA_output89_A _12693_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11388_ _11388_/A _11388_/B vssd1 vssd1 vccd1 vccd1 _11388_/X sky130_fd_sc_hd__and2_1
XANTENNA__13439__B _13725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17626__S _17628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _20031_/Q _19869_/Q _19278_/Q _19048_/Q _10330_/S _10223_/X vssd1 vssd1 vccd1
+ vccd1 _10340_/B sky130_fd_sc_hd__mux4_1
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13127_ _18560_/Q _13070_/A _13082_/X _14476_/B vssd1 vssd1 vccd1 vccd1 _13127_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16530__S _16530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18984_ _19523_/CLK _18984_/D vssd1 vssd1 vccd1 vccd1 _18984_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _19838_/Q _17068_/X _17937_/S vssd1 vssd1 vccd1 vccd1 _17936_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09933__A _09933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _18721_/Q vssd1 vssd1 vccd1 vccd1 _14468_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12511__A1 _12082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12009_ _15633_/B vssd1 vssd1 vccd1 vccd1 _12722_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17866_ _17866_/A vssd1 vssd1 vccd1 vccd1 _19807_/D sky130_fd_sc_hd__clkbuf_1
X_19605_ _19828_/CLK _19605_/D vssd1 vssd1 vccd1 vccd1 _19605_/Q sky130_fd_sc_hd__dfxtp_1
X_16817_ _16374_/X _19375_/Q _16819_/S vssd1 vssd1 vccd1 vccd1 _16818_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17797_ _17797_/A vssd1 vssd1 vccd1 vccd1 _19776_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16766__A _16834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17361__S _17365_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19536_ _19986_/CLK _19536_/D vssd1 vssd1 vccd1 vccd1 _19536_/Q sky130_fd_sc_hd__dfxtp_1
X_16748_ _16748_/A vssd1 vssd1 vccd1 vccd1 _19344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11173__S1 _11172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19467_ _20022_/CLK _19467_/D vssd1 vssd1 vccd1 vccd1 _19467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16679_ _16384_/X _19314_/Q _16685_/S vssd1 vssd1 vccd1 vccd1 _16680_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09220_ _09283_/B vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18418_ _17729_/X _20038_/Q _18418_/S vssd1 vssd1 vccd1 vccd1 _18419_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15764__A1 _09454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19398_ _19985_/CLK _19398_/D vssd1 vssd1 vccd1 vccd1 _19398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17597__A _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18349_ _18349_/A vssd1 vssd1 vccd1 vccd1 _20007_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10589__B1 _10674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput60 io_ibus_inst[4] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10987__S1 _10973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10054__A _10054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16440__S _16446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09984_ _10266_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _09984_/X sky130_fd_sc_hd__or2_1
XFILLER_104_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18221__A _18278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09843__A _09843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10513__B1 _10078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15580__A _15602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12709__A _15974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_169_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13304__S _13366_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10911__S1 _10893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09418_ _18824_/Q _09418_/B vssd1 vssd1 vccd1 vccd1 _11722_/A sky130_fd_sc_hd__and2_1
XFILLER_41_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10690_ _10690_/A _10690_/B vssd1 vssd1 vccd1 vccd1 _10690_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09349_ _18831_/Q _12895_/A _18832_/Q vssd1 vssd1 vccd1 vccd1 _09349_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16615__S _16617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12360_ _12360_/A _14883_/A vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ _11311_/A _11311_/B vssd1 vssd1 vccd1 vccd1 _11311_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11792__A2 _11815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12291_ _18968_/Q _14805_/A _14812_/B _12290_/X vssd1 vssd1 vccd1 vccd1 _12291_/X
+ sky130_fd_sc_hd__a211o_1
X_14030_ _14046_/A _14034_/C vssd1 vssd1 vccd1 vccd1 _14030_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11242_ _11242_/A _11242_/B vssd1 vssd1 vccd1 vccd1 _11242_/X sky130_fd_sc_hd__or2_1
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11173_ _19196_/Q _19787_/Q _19949_/Q _19164_/Q _11171_/X _11172_/X vssd1 vssd1 vccd1
+ vccd1 _11174_/B sky130_fd_sc_hd__mux4_1
XFILLER_161_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16350__S _16362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10124_ _10543_/S vssd1 vssd1 vccd1 vccd1 _10125_/S sky130_fd_sc_hd__buf_4
XANTENNA_input40_A io_ibus_inst[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15474__B _15474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15981_ _19024_/Q _15936_/A _15928_/A _15980_/Y vssd1 vssd1 vccd1 vccd1 _19024_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17720_ _17720_/A vssd1 vssd1 vccd1 vccd1 _17720_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10055_ _19679_/Q _19445_/Q _18510_/Q _19775_/Q _10254_/A _10054_/X vssd1 vssd1 vccd1
+ vccd1 _10055_/X sky130_fd_sc_hd__mux4_1
X_14932_ _14926_/X _14930_/X _15041_/S vssd1 vssd1 vccd1 vccd1 _14932_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17651_ _17651_/A vssd1 vssd1 vccd1 vccd1 _19723_/D sky130_fd_sc_hd__clkbuf_1
X_14863_ _14863_/A vssd1 vssd1 vccd1 vccd1 _15436_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_91_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output127_A _12858_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16602_ _19280_/Q _13835_/X _16602_/S vssd1 vssd1 vccd1 vccd1 _16603_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17181__S _17193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13814_ _18503_/Q _13813_/X _13820_/S vssd1 vssd1 vccd1 vccd1 _13815_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17582_ _17125_/X _19695_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17583_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14794_ _18830_/Q _14789_/B _15765_/A _11956_/A vssd1 vssd1 vccd1 vccd1 _14795_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_16_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19321_ _19526_/CLK _19321_/D vssd1 vssd1 vccd1 vccd1 _19321_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10807__A1 _09830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16533_ _19249_/Q _13838_/X _16541_/S vssd1 vssd1 vccd1 vccd1 _16534_/A sky130_fd_sc_hd__mux2_1
X_13745_ _13745_/A vssd1 vssd1 vccd1 vccd1 _18484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10957_ _19329_/Q _19600_/Q _19824_/Q _19568_/Q _10892_/X _10893_/X vssd1 vssd1 vccd1
+ vccd1 _10957_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11507__A1_N _18846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19252_ _19747_/CLK _19252_/D vssd1 vssd1 vccd1 vccd1 _19252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16464_ _19219_/Q _13845_/X _16468_/S vssd1 vssd1 vccd1 vccd1 _16465_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15746__A1 _09458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13676_ _13732_/A _19015_/Q vssd1 vssd1 vccd1 vccd1 _13676_/Y sky130_fd_sc_hd__nand2_1
X_10888_ _11473_/A _10887_/X _10719_/A vssd1 vssd1 vccd1 vccd1 _10888_/Y sky130_fd_sc_hd__o21ai_1
X_18203_ _18203_/A vssd1 vssd1 vccd1 vccd1 _19942_/D sky130_fd_sc_hd__clkbuf_1
X_15415_ _15478_/A _15415_/B vssd1 vssd1 vccd1 vccd1 _15415_/X sky130_fd_sc_hd__or2_1
X_19183_ _20030_/CLK _19183_/D vssd1 vssd1 vccd1 vccd1 _19183_/Q sky130_fd_sc_hd__dfxtp_1
X_12627_ _12522_/X _12625_/X _12626_/X _12480_/X vssd1 vssd1 vccd1 vccd1 _12627_/X
+ sky130_fd_sc_hd__o211a_1
X_16395_ _16395_/A vssd1 vssd1 vccd1 vccd1 _19189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14834__A _15183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12835__A_N _12833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18134_ _18133_/X _19912_/Q _18134_/S vssd1 vssd1 vccd1 vccd1 _18135_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15346_ _15346_/A vssd1 vssd1 vccd1 vccd1 _15346_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _18474_/Q _12556_/X _12557_/X vssd1 vssd1 vccd1 vccd1 _12558_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_156_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13509__B1 _16069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11509_ _15940_/C _12842_/A vssd1 vssd1 vccd1 vccd1 _11510_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18065_ _18063_/X _19891_/Q _18078_/S vssd1 vssd1 vccd1 vccd1 _18066_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15277_ _18843_/Q _09433_/X _15276_/X vssd1 vssd1 vccd1 vccd1 _18843_/D sky130_fd_sc_hd__o21a_1
X_12489_ _15373_/A _12458_/Y _15385_/A _12632_/A vssd1 vssd1 vccd1 vccd1 _12490_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_7_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17016_ _17016_/A vssd1 vssd1 vccd1 vccd1 _19459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14228_ _12065_/B _12918_/B _14227_/X _09345_/A vssd1 vssd1 vccd1 vccd1 _14242_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_160_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14159_ _14159_/A vssd1 vssd1 vccd1 vccd1 _14427_/A sky130_fd_sc_hd__clkbuf_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09663__A _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ _18967_/CLK _18967_/D vssd1 vssd1 vccd1 vccd1 _18967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11299__A1 _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17918_ _19830_/Q _17042_/X _17926_/S vssd1 vssd1 vccd1 vccd1 _17919_/A sky130_fd_sc_hd__mux2_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18898_ _18997_/CLK _18898_/D vssd1 vssd1 vccd1 vccd1 _18898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17849_ _17849_/A vssd1 vssd1 vccd1 vccd1 _19799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18187__S _18191_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17091__S _17094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11146__S1 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19519_ _20038_/CLK _19519_/D vssd1 vssd1 vccd1 vccd1 _19519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_170_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10274__A2 _10264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15737__A1 hold4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09203_ _11961_/A _12003_/B _14761_/B vssd1 vssd1 vccd1 vccd1 _11956_/A sky130_fd_sc_hd__or3_4
XFILLER_50_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16435__S _16435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10049__A _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13212__A2 _11815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11223__A1 _18837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12971__A1 _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12723__A1 _12522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_95_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09967_ _10313_/S vssd1 vssd1 vccd1 vccd1 _09967_/X sky130_fd_sc_hd__buf_4
XFILLER_131_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10512__A _18851_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09898_ _19253_/Q _19748_/Q _09898_/S vssd1 vssd1 vccd1 vccd1 _09898_/X sky130_fd_sc_hd__mux2_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14779__A2 _14766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ _11860_/A _11860_/B _11860_/C _11860_/D vssd1 vssd1 vccd1 vccd1 _11860_/X
+ sky130_fd_sc_hd__or4_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _11502_/A _10810_/X _09793_/A vssd1 vssd1 vccd1 vccd1 _10811_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13542__B _13542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11791_ _11791_/A vssd1 vssd1 vccd1 vccd1 _12876_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13530_ _13747_/A vssd1 vssd1 vccd1 vccd1 _13531_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10742_ _20023_/Q _19861_/Q _19270_/Q _19040_/Q _09725_/A _10009_/A vssd1 vssd1 vccd1
+ vccd1 _10743_/B sky130_fd_sc_hd__mux4_1
XFILLER_43_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10673_ _19207_/Q _19798_/Q _19960_/Q _19175_/Q _09652_/A _10656_/A vssd1 vssd1 vccd1
+ vccd1 _10674_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13461_ _12967_/X _13446_/X _13450_/Y _13460_/Y vssd1 vssd1 vccd1 vccd1 _17087_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15200_ _15198_/X _15199_/X _15298_/S vssd1 vssd1 vccd1 vccd1 _15200_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17030__A _17030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ _12389_/A _12389_/B _12386_/A vssd1 vssd1 vccd1 vccd1 _12413_/B sky130_fd_sc_hd__a21bo_1
XFILLER_139_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16180_ _13161_/X _19108_/Q _16184_/S vssd1 vssd1 vccd1 vccd1 _16181_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09748__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13392_ _13699_/A _13390_/C _13714_/A vssd1 vssd1 vccd1 vccd1 _13393_/B sky130_fd_sc_hd__a21oi_1
X_15131_ _15129_/X _15130_/X _15280_/S vssd1 vssd1 vccd1 vccd1 _15131_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12343_ _12722_/B vssd1 vssd1 vccd1 vccd1 _12343_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15062_ _14888_/X _14867_/X _15118_/S vssd1 vssd1 vccd1 vccd1 _15062_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12274_ _18528_/Q _12303_/B vssd1 vssd1 vccd1 vccd1 _12287_/A sky130_fd_sc_hd__or2_1
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14013_ _18579_/Q _18578_/Q _14013_/C vssd1 vssd1 vccd1 vccd1 _14016_/B sky130_fd_sc_hd__and3_1
X_11225_ _11225_/A _11225_/B vssd1 vssd1 vccd1 vccd1 _11225_/X sky130_fd_sc_hd__or2_1
X_19870_ _20030_/CLK _19870_/D vssd1 vssd1 vccd1 vccd1 _19870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18821_ _19887_/CLK _18821_/D vssd1 vssd1 vccd1 vccd1 _18821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11156_ _19358_/Q _19693_/Q _11156_/S vssd1 vssd1 vccd1 vccd1 _11157_/B sky130_fd_sc_hd__mux2_1
XFILLER_150_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10107_ _10107_/A vssd1 vssd1 vccd1 vccd1 _10107_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17904__S _17904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18752_ _18762_/CLK _18752_/D vssd1 vssd1 vccd1 vccd1 _18752_/Q sky130_fd_sc_hd__dfxtp_1
X_15964_ _15964_/A _15964_/B vssd1 vssd1 vccd1 vccd1 _15964_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11087_ _19199_/Q _19790_/Q _19952_/Q _19167_/Q _11023_/S _11296_/A vssd1 vssd1 vccd1
+ vccd1 _11088_/B sky130_fd_sc_hd__mux4_1
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17703_ _17703_/A vssd1 vssd1 vccd1 vccd1 _19739_/D sky130_fd_sc_hd__clkbuf_1
X_10038_ _10028_/X _10037_/X _10342_/A vssd1 vssd1 vccd1 vccd1 _10038_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11376__S1 _11322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14915_ _15138_/B _12713_/B _14915_/S vssd1 vssd1 vccd1 vccd1 _14915_/X sky130_fd_sc_hd__mux2_1
X_18683_ _18687_/CLK _18683_/D vssd1 vssd1 vccd1 vccd1 _18683_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15932__B _15942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15895_ _15895_/A vssd1 vssd1 vccd1 vccd1 _18991_/D sky130_fd_sc_hd__clkbuf_1
X_17634_ _17634_/A vssd1 vssd1 vccd1 vccd1 _17634_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14846_ _14990_/C _14846_/B vssd1 vssd1 vccd1 vccd1 _15151_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17565_ _17097_/X _19687_/Q _17573_/S vssd1 vssd1 vccd1 vccd1 _17566_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14777_ _14777_/A vssd1 vssd1 vccd1 vccd1 _18825_/D sky130_fd_sc_hd__clkbuf_1
X_11989_ _11452_/A _18899_/Q _12039_/A vssd1 vssd1 vccd1 vccd1 _14898_/A sky130_fd_sc_hd__mux2_2
X_19304_ _19828_/CLK _19304_/D vssd1 vssd1 vccd1 vccd1 _19304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16516_ _16516_/A vssd1 vssd1 vccd1 vccd1 _19241_/D sky130_fd_sc_hd__clkbuf_1
X_13728_ _12422_/X _13727_/X _13514_/S vssd1 vssd1 vccd1 vccd1 _13728_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__10887__S0 _10776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17496_ _17198_/X _19654_/Q _17496_/S vssd1 vssd1 vccd1 vccd1 _17497_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19235_ _19861_/CLK _19235_/D vssd1 vssd1 vccd1 vccd1 _19235_/Q sky130_fd_sc_hd__dfxtp_1
X_16447_ _16447_/A vssd1 vssd1 vccd1 vccd1 _19211_/D sky130_fd_sc_hd__clkbuf_1
X_13659_ _13732_/A _19013_/Q vssd1 vssd1 vccd1 vccd1 _13659_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09658__A _09918_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19166_ _20015_/CLK _19166_/D vssd1 vssd1 vccd1 vccd1 _19166_/Q sky130_fd_sc_hd__dfxtp_1
X_16378_ _16377_/X _19184_/Q _16378_/S vssd1 vssd1 vccd1 vccd1 _16379_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12106__B_N _12134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11300__S1 _11172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18117_ _18117_/A vssd1 vssd1 vccd1 vccd1 _19906_/D sky130_fd_sc_hd__clkbuf_1
X_15329_ _15419_/A vssd1 vssd1 vccd1 vccd1 _15329_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19097_ _19978_/CLK _19097_/D vssd1 vssd1 vccd1 vccd1 _19097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18048_ _18046_/X _19886_/Q _18061_/S vssd1 vssd1 vccd1 vccd1 _18049_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_117_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20010_ _20010_/CLK _20010_/D vssd1 vssd1 vccd1 vccd1 _20010_/Q sky130_fd_sc_hd__dfxtp_1
X_09821_ _09821_/A vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__buf_2
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13627__B _13627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15655__A0 _18906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19999_ _19999_/CLK _19999_/D vssd1 vssd1 vccd1 vccd1 _19999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09752_ _11404_/A vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09683_ _09683_/A vssd1 vssd1 vccd1 vccd1 _10719_/A sky130_fd_sc_hd__buf_2
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19948_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13418__C1 _13416_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13433__A2 _13269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11444__A1 _11086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16165__S _16173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09568__A _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14697__A1 _13591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11055__S0 _11367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12722__A _18481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11010_ _11001_/Y _11004_/Y _11006_/Y _11008_/Y _11133_/A vssd1 vssd1 vccd1 vccd1
+ _11010_/X sky130_fd_sc_hd__o221a_1
XFILLER_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17724__S _17730_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10242__A _15972_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11358__S1 _11357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12961_ _13223_/A _12958_/X _12960_/Y input23/X _12906_/X vssd1 vssd1 vccd1 vccd1
+ _17001_/A sky130_fd_sc_hd__a32o_4
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _14700_/A vssd1 vssd1 vccd1 vccd1 _18801_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _11912_/A vssd1 vssd1 vccd1 vccd1 _15633_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18060__A1 _13579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _18917_/Q _12554_/A _15688_/S vssd1 vssd1 vccd1 vccd1 _15681_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _18550_/Q _12877_/X _12886_/X _12888_/X _12891_/X vssd1 vssd1 vccd1 vccd1
+ _12892_/X sky130_fd_sc_hd__a2111o_2
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _14648_/A vssd1 vssd1 vccd1 vccd1 _14646_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10388__S _10388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _12879_/A vssd1 vssd1 vccd1 vccd1 _11843_/X sky130_fd_sc_hd__buf_2
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11073__A _11073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _17195_/X _19589_/Q _17352_/S vssd1 vssd1 vccd1 vccd1 _17351_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _13531_/A _18995_/Q _09341_/X _14561_/X vssd1 vssd1 vccd1 vccd1 _14562_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11774_ _11774_/A _11860_/B vssd1 vssd1 vccd1 vccd1 _11774_/X sky130_fd_sc_hd__and2_1
XFILLER_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16400_/S vssd1 vssd1 vccd1 vccd1 _16314_/S sky130_fd_sc_hd__buf_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13520_/A vssd1 vssd1 vccd1 vccd1 _13514_/S sky130_fd_sc_hd__clkbuf_2
X_10725_ _10919_/S vssd1 vssd1 vccd1 vccd1 _10821_/S sky130_fd_sc_hd__clkbuf_4
X_17281_ _17281_/A vssd1 vssd1 vccd1 vccd1 _19558_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14493_ _18731_/Q _14493_/B _14493_/C vssd1 vssd1 vccd1 vccd1 _14495_/B sky130_fd_sc_hd__and3_1
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19020_ _19023_/CLK _19020_/D vssd1 vssd1 vccd1 vccd1 _19020_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11801__A _11801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16232_ _12963_/X _19130_/Q _16236_/S vssd1 vssd1 vccd1 vccd1 _16233_/A sky130_fd_sc_hd__mux2_1
X_13444_ _13443_/X _18452_/Q _13464_/S vssd1 vssd1 vccd1 vccd1 _13445_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10656_ _10656_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10656_/X sky130_fd_sc_hd__and2_1
XFILLER_139_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12935__A1 _12875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16163_ _16163_/A vssd1 vssd1 vccd1 vccd1 _19100_/D sky130_fd_sc_hd__clkbuf_1
X_10587_ _10587_/A _10587_/B vssd1 vssd1 vccd1 vccd1 _10587_/Y sky130_fd_sc_hd__nand2_1
X_13375_ _18815_/Q _13269_/X _11843_/X _18782_/Q _13374_/X vssd1 vssd1 vccd1 vccd1
+ _13375_/X sky130_fd_sc_hd__a221o_1
XFILLER_126_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15114_ _15019_/X _15032_/X _15114_/S vssd1 vssd1 vccd1 vccd1 _15114_/X sky130_fd_sc_hd__mux2_1
X_12326_ _15938_/C _18909_/Q _12409_/A vssd1 vssd1 vccd1 vccd1 _14885_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16094_ _13042_/X _19070_/Q _16100_/S vssd1 vssd1 vccd1 vccd1 _16095_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14688__A1 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19922_ _20018_/CLK _19922_/D vssd1 vssd1 vccd1 vccd1 _19922_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11046__S0 _10977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15045_ _15068_/A vssd1 vssd1 vccd1 vccd1 _15247_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12257_ _12188_/X _12251_/X _12252_/X _12256_/Y vssd1 vssd1 vccd1 vccd1 _12258_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output71_A _12871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _11208_/A vssd1 vssd1 vccd1 vccd1 _11208_/X sky130_fd_sc_hd__clkbuf_4
X_12188_ _12188_/A vssd1 vssd1 vccd1 vccd1 _12188_/X sky130_fd_sc_hd__buf_2
X_19853_ _19853_/CLK _19853_/D vssd1 vssd1 vccd1 vccd1 _19853_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10174__A1 _10162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15943__A _15964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18804_ _19912_/CLK _18804_/D vssd1 vssd1 vccd1 vccd1 _18804_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10152__A _10208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ _19198_/Q _19789_/Q _19951_/Q _19166_/Q _11049_/S _10973_/A vssd1 vssd1 vccd1
+ vccd1 _11140_/B sky130_fd_sc_hd__mux4_1
X_19784_ _19946_/CLK _19784_/D vssd1 vssd1 vccd1 vccd1 _19784_/Q sky130_fd_sc_hd__dfxtp_1
X_16996_ _19453_/Q _16992_/X _17008_/S vssd1 vssd1 vccd1 vccd1 _16997_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13112__A1 _13350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18735_ _20005_/CLK _18735_/D vssd1 vssd1 vccd1 vccd1 _18735_/Q sky130_fd_sc_hd__dfxtp_1
X_15947_ _15966_/A _15966_/B _15947_/C vssd1 vssd1 vccd1 vccd1 _15947_/X sky130_fd_sc_hd__and3_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13663__A2 _13517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18666_ _19683_/CLK _18666_/D vssd1 vssd1 vccd1 vccd1 _18666_/Q sky130_fd_sc_hd__dfxtp_1
X_15878_ _15878_/A vssd1 vssd1 vccd1 vccd1 _18986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17617_ _17176_/X _19711_/Q _17617_/S vssd1 vssd1 vccd1 vccd1 _17618_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14829_ _15546_/A vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__clkbuf_2
X_18597_ _19941_/CLK _18597_/D vssd1 vssd1 vccd1 vccd1 _18597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13415__A2 _13269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17548_ _19680_/Q vssd1 vssd1 vccd1 vccd1 _17549_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_43_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17479_ _17173_/X _19646_/Q _17481_/S vssd1 vssd1 vccd1 vccd1 _17480_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12807__A _15553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19218_ _19971_/CLK _19218_/D vssd1 vssd1 vccd1 vccd1 _19218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11729__A2 _11724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19149_ _19966_/CLK _19149_/D vssd1 vssd1 vccd1 vccd1 _19149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14679__A1 _13508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13351__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ _09804_/A vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11901__A2 _11884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09851__A _09851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09735_ _11019_/A vssd1 vssd1 vccd1 vccd1 _11172_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_153_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19062_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09666_ _10448_/A vssd1 vssd1 vccd1 vccd1 _10355_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09597_ _09597_/A vssd1 vssd1 vccd1 vccd1 _09668_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12614__A0 _15966_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__A1 _11206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_168_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _18868_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10510_ _09988_/A _10509_/X _09687_/A vssd1 vssd1 vccd1 vccd1 _10510_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__14367__B1 _14366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11490_ _19668_/Q _19434_/Q _18499_/Q _19764_/Q _10797_/X _11487_/A vssd1 vssd1 vccd1
+ vccd1 _11490_/X sky130_fd_sc_hd__mux4_1
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ _10434_/Y _10436_/Y _10438_/Y _10440_/Y _09821_/A vssd1 vssd1 vccd1 vccd1
+ _10441_/X sky130_fd_sc_hd__o221a_1
X_10372_ _10365_/X _10367_/X _10369_/X _10371_/X _09876_/A vssd1 vssd1 vccd1 vccd1
+ _10372_/X sky130_fd_sc_hd__a221o_2
XFILLER_137_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13160_ _17033_/A vssd1 vssd1 vccd1 vccd1 _17675_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15867__B1 _15788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12111_ _12108_/Y _12109_/X _12110_/Y vssd1 vssd1 vccd1 vccd1 _12111_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_124_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13091_ _13091_/A vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12452__A _12452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13342__A1 _13005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ _12042_/A _14895_/A vssd1 vssd1 vccd1 vccd1 _12043_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_106_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _20035_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13267__B _18884_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__B1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15763__A _18951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16850_ _16918_/S vssd1 vssd1 vccd1 vccd1 _16859_/S sky130_fd_sc_hd__buf_2
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15801_ _15801_/A vssd1 vssd1 vccd1 vccd1 _18963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15482__B _15482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16781_ _16781_/A vssd1 vssd1 vccd1 vccd1 _19358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13993_ _14010_/A _13999_/C vssd1 vssd1 vccd1 vccd1 _13993_/Y sky130_fd_sc_hd__nor2_1
X_18520_ _18526_/CLK _18520_/D vssd1 vssd1 vccd1 vccd1 _18520_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _16691_/B _15732_/B vssd1 vssd1 vccd1 vccd1 _15732_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12944_ _12944_/A vssd1 vssd1 vccd1 vccd1 _12944_/X sky130_fd_sc_hd__buf_2
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _19942_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11120__A3 _11118_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11515__B _12848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15663_ _15663_/A vssd1 vssd1 vccd1 vccd1 _18909_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18285__S _18291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12875_ _13473_/A vssd1 vssd1 vccd1 vccd1 _12875_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _17402_/A vssd1 vssd1 vccd1 vccd1 _19611_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _14648_/A vssd1 vssd1 vccd1 vccd1 _14629_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18382_ _18382_/A vssd1 vssd1 vccd1 vccd1 _20021_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _18561_/Q _12876_/A _13194_/A _18725_/Q vssd1 vssd1 vccd1 vccd1 _11826_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _13630_/A _18911_/Q _15600_/S vssd1 vssd1 vccd1 vccd1 _15595_/A sky130_fd_sc_hd__mux2_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17333_ _17170_/X _19581_/Q _17337_/S vssd1 vssd1 vccd1 vccd1 _17334_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11503__S1 _10856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _18754_/Q _11865_/X _14544_/X _14540_/X vssd1 vssd1 vccd1 vccd1 _18754_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _18472_/Q _11755_/X _14672_/A _18808_/Q _11756_/X vssd1 vssd1 vccd1 vccd1
+ _11757_/X sky130_fd_sc_hd__a221o_1
XFILLER_42_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17264_ _17264_/A vssd1 vssd1 vccd1 vccd1 _19550_/D sky130_fd_sc_hd__clkbuf_1
X_10708_ _10919_/S vssd1 vssd1 vccd1 vccd1 _10708_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14476_ _18725_/Q _14476_/B _14476_/C vssd1 vssd1 vccd1 vccd1 _14478_/B sky130_fd_sc_hd__and3_1
X_11688_ _11688_/A _11785_/A vssd1 vssd1 vccd1 vccd1 _11734_/A sky130_fd_sc_hd__nor2_2
X_19003_ _19488_/CLK _19003_/D vssd1 vssd1 vccd1 vccd1 _19003_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_174_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16215_ _13443_/X _19124_/Q _16217_/S vssd1 vssd1 vccd1 vccd1 _16216_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14264__D _14264_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15938__A _15940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13427_ _18892_/Q _18893_/Q _13427_/C vssd1 vssd1 vccd1 vccd1 _13449_/B sky130_fd_sc_hd__and3_1
XFILLER_174_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10639_ _19368_/Q _19703_/Q _10749_/S vssd1 vssd1 vccd1 vccd1 _10639_/X sky130_fd_sc_hd__mux2_1
X_17195_ _17732_/A vssd1 vssd1 vccd1 vccd1 _17195_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__10147__A _10843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16533__S _16541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16146_ _13481_/X _19094_/Q _16148_/S vssd1 vssd1 vccd1 vccd1 _16147_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13358_ _13688_/A _13357_/C _18889_/Q vssd1 vssd1 vccd1 vccd1 _13359_/C sky130_fd_sc_hd__a21o_1
XFILLER_6_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10395__A1 _10162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12309_ _18768_/Q _18767_/Q _12309_/C vssd1 vssd1 vccd1 vccd1 _12374_/C sky130_fd_sc_hd__and3_1
XFILLER_115_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16077_ _16077_/A vssd1 vssd1 vccd1 vccd1 _19063_/D sky130_fd_sc_hd__clkbuf_1
X_13289_ _13289_/A _13289_/B _13326_/C vssd1 vssd1 vccd1 vccd1 _13289_/X sky130_fd_sc_hd__or3_2
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15028_ _14864_/X _14870_/X _15032_/S vssd1 vssd1 vccd1 vccd1 _15028_/X sky130_fd_sc_hd__mux2_1
X_19905_ _19910_/CLK _19905_/D vssd1 vssd1 vccd1 vccd1 _19905_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13333__B2 _13332_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19836_ _19836_/CLK _19836_/D vssd1 vssd1 vccd1 vccd1 _19836_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11895__A1 _18670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16283__A0 _13385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _20007_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09671__A _10254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19767_ _19767_/CLK _19767_/D vssd1 vssd1 vccd1 vccd1 _19767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16979_ _16979_/A vssd1 vssd1 vccd1 vccd1 _19446_/D sky130_fd_sc_hd__clkbuf_1
Xinput3 io_dbus_rdata[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
X_09520_ _14756_/B _09520_/B vssd1 vssd1 vccd1 vccd1 _14819_/B sky130_fd_sc_hd__or2_1
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09390__B _11869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18718_ _18719_/CLK _18718_/D vssd1 vssd1 vccd1 vccd1 _18718_/Q sky130_fd_sc_hd__dfxtp_1
X_19698_ _19732_/CLK _19698_/D vssd1 vssd1 vccd1 vccd1 _19698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09451_ _12033_/S vssd1 vssd1 vccd1 vccd1 _15899_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18649_ _18688_/CLK _18649_/D vssd1 vssd1 vccd1 vccd1 _18649_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16708__S _16714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19706_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09382_ _18949_/Q vssd1 vssd1 vccd1 vccd1 _11699_/A sky130_fd_sc_hd__inv_2
XFILLER_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10057__A _10057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13572__B2 _19002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19856_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13368__A _13368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10491__S _10493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10481__S1 _10223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10138__A1 _10194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17274__S _17276_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11430__S0 _11356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19827_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14199__A _14245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09718_ _11153_/A vssd1 vssd1 vccd1 vccd1 _10960_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ _11212_/A vssd1 vssd1 vccd1 vccd1 _11049_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09649_ _10872_/S vssd1 vssd1 vccd1 vccd1 _09650_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14927__A _14927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12660_ _09261_/B _12657_/X _12682_/A _12659_/Y vssd1 vssd1 vccd1 vccd1 _15487_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11611_/A _11611_/B _11611_/C _11610_/X vssd1 vssd1 vccd1 vccd1 _11611_/X
+ sky130_fd_sc_hd__or4b_1
XANTENNA__11497__S0 _11486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12591_ _12591_/A _15449_/A vssd1 vssd1 vccd1 vccd1 _12619_/A sky130_fd_sc_hd__xnor2_2
X_14330_ _14413_/A _14338_/D vssd1 vssd1 vccd1 vccd1 _14330_/Y sky130_fd_sc_hd__nor2_1
X_11542_ _19223_/Q _19814_/Q _19976_/Q _19191_/Q _11534_/S _09660_/A vssd1 vssd1 vccd1
+ vccd1 _11543_/B sky130_fd_sc_hd__mux4_2
XFILLER_168_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15758__A _15758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11249__S0 _11212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14261_ _18655_/Q _14279_/B _14264_/D vssd1 vssd1 vccd1 vccd1 _14262_/B sky130_fd_sc_hd__and3_1
X_11473_ _11473_/A _11473_/B vssd1 vssd1 vccd1 vccd1 _11473_/X sky130_fd_sc_hd__or2_1
XANTENNA__16353__S _16362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13012__B1 _11855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16000_ _16057_/S vssd1 vssd1 vccd1 vccd1 _16009_/S sky130_fd_sc_hd__clkbuf_4
X_13212_ _18661_/Q _11815_/A _11794_/X _18629_/Q vssd1 vssd1 vccd1 vccd1 _13212_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input70_A reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ _10424_/A _10424_/B vssd1 vssd1 vccd1 vccd1 _10424_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14192_ _18636_/Q _14190_/B _14191_/Y vssd1 vssd1 vccd1 vccd1 _18636_/D sky130_fd_sc_hd__o21a_1
XFILLER_100_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13143_ _18876_/Q _13143_/B vssd1 vssd1 vccd1 vccd1 _13174_/C sky130_fd_sc_hd__and2_1
X_10355_ _10355_/A _10355_/B vssd1 vssd1 vccd1 vccd1 _10355_/X sky130_fd_sc_hd__and2_1
XFILLER_140_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10286_ _19151_/Q _19412_/Q _19311_/Q _19646_/Q _10279_/X _10283_/X vssd1 vssd1 vccd1
+ vccd1 _10287_/B sky130_fd_sc_hd__mux4_1
X_17951_ _17951_/A vssd1 vssd1 vccd1 vccd1 _19845_/D sky130_fd_sc_hd__clkbuf_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _12231_/A _12984_/A _13073_/X vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output157_A _12631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17184__S _17193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16902_ _16902_/A vssd1 vssd1 vccd1 vccd1 _19412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12025_ _12350_/A vssd1 vssd1 vccd1 vccd1 _12402_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10224__S1 _10223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17882_ _18208_/A _17882_/B vssd1 vssd1 vccd1 vccd1 _17939_/A sky130_fd_sc_hd__nor2_2
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12910__A _18937_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19621_ _19975_/CLK _19621_/D vssd1 vssd1 vccd1 vccd1 _19621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16833_ _16833_/A vssd1 vssd1 vccd1 vccd1 _19382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13079__B1 _11687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13725__B _13725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__A _15978_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764_ _18280_/A _17635_/A vssd1 vssd1 vccd1 vccd1 _16821_/A sky130_fd_sc_hd__or2_2
X_19552_ _20002_/CLK _19552_/D vssd1 vssd1 vccd1 vccd1 _19552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13976_ _18566_/Q _13976_/B vssd1 vssd1 vccd1 vccd1 _13982_/C sky130_fd_sc_hd__and2_1
XFILLER_19_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14838__B_N _15004_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18503_ _20024_/CLK _18503_/D vssd1 vssd1 vccd1 vccd1 _18503_/Q sky130_fd_sc_hd__dfxtp_1
X_15715_ _18933_/Q _15715_/B vssd1 vssd1 vccd1 vccd1 _15715_/X sky130_fd_sc_hd__or2_1
XFILLER_74_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12927_ _18791_/Q _12880_/X _12881_/X _18679_/Q _12926_/X vssd1 vssd1 vccd1 vccd1
+ _12927_/X sky130_fd_sc_hd__a221o_1
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15940__B _15955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19483_ _20007_/CLK _19483_/D vssd1 vssd1 vccd1 vccd1 _19483_/Q sky130_fd_sc_hd__dfxtp_1
X_16695_ _19320_/Q _13754_/X _16703_/S vssd1 vssd1 vccd1 vccd1 _16696_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16528__S _16530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18434_ _19664_/CLK _18434_/D vssd1 vssd1 vccd1 vccd1 _18434_/Q sky130_fd_sc_hd__dfxtp_1
X_15646_ _15703_/S vssd1 vssd1 vccd1 vccd1 _15655_/S sky130_fd_sc_hd__clkbuf_2
X_12858_ _12863_/A _12858_/B vssd1 vssd1 vccd1 vccd1 _12858_/Y sky130_fd_sc_hd__nor2_2
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11809_ _15633_/A _15786_/B vssd1 vssd1 vccd1 vccd1 _14792_/B sky130_fd_sc_hd__nand2_2
X_18365_ _18422_/S vssd1 vssd1 vccd1 vccd1 _18374_/S sky130_fd_sc_hd__clkbuf_4
X_15577_ _15577_/A vssd1 vssd1 vccd1 vccd1 _18871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12789_/A _12789_/B vssd1 vssd1 vccd1 vccd1 _12791_/B sky130_fd_sc_hd__xnor2_4
XFILLER_42_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17316_/A vssd1 vssd1 vccd1 vccd1 _19573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14528_ _14528_/A _14528_/B _14528_/C vssd1 vssd1 vccd1 vccd1 _18743_/D sky130_fd_sc_hd__nor3_1
XFILLER_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18296_ _17656_/X _19983_/Q _18302_/S vssd1 vssd1 vccd1 vccd1 _18297_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17247_ _17247_/A vssd1 vssd1 vccd1 vccd1 _19542_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17359__S _17365_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15668__A _15690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16263__S _16269_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__A3 _10076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14459_ _18719_/Q _14459_/B _14459_/C vssd1 vssd1 vccd1 vccd1 _14461_/B sky130_fd_sc_hd__and3_1
XFILLER_116_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09666__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17178_ _17178_/A vssd1 vssd1 vccd1 vccd1 _19514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14751__B1 _12833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16129_ _13344_/X _19086_/Q _16133_/S vssd1 vssd1 vccd1 vccd1 _16130_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10463__S1 _10400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11200__S _11270_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16499__A _16545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17094__S _17094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15607__S _15611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11868__A1 _12060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19819_ _19948_/CLK _19819_/D vssd1 vssd1 vccd1 vccd1 _19819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09503_ _14804_/B _14804_/C vssd1 vssd1 vccd1 vccd1 _09504_/C sky130_fd_sc_hd__nor2_1
XFILLER_71_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16438__S _16446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09434_ _09434_/A vssd1 vssd1 vccd1 vccd1 _11925_/B sky130_fd_sc_hd__buf_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _18825_/Q _18824_/Q vssd1 vssd1 vccd1 vccd1 _09423_/B sky130_fd_sc_hd__or2_1
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09296_ _18979_/Q _18939_/Q vssd1 vssd1 vccd1 vccd1 _09296_/X sky130_fd_sc_hd__xor2_1
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16173__S _16173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13098__A _17662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09295__B _18940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16901__S _16903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10454__S1 _10400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11110__S _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _10172_/A vssd1 vssd1 vccd1 vccd1 _10392_/A sky130_fd_sc_hd__buf_2
XFILLER_133_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_165_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput170 _12173_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[6] sky130_fd_sc_hd__buf_2
XFILLER_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13826__A _17062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ _10064_/X _10070_/X _09567_/A vssd1 vssd1 vccd1 vccd1 _10071_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11859__B2 _19006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09921__B1 _10073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13545__B _18999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ _18508_/Q _13829_/X _13836_/S vssd1 vssd1 vccd1 vccd1 _13831_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ _13761_/A vssd1 vssd1 vccd1 vccd1 _18486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10973_ _10973_/A vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__buf_2
XFILLER_16_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15500_ _15522_/A _15500_/B _15500_/C vssd1 vssd1 vccd1 vccd1 _15500_/X sky130_fd_sc_hd__and3_1
XANTENNA__17033__A _17033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ _12713_/A _15509_/B vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__nor2_1
X_16480_ _19225_/Q _13762_/X _16486_/S vssd1 vssd1 vccd1 vccd1 _16481_/A sky130_fd_sc_hd__mux2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13692_ _13692_/A vssd1 vssd1 vccd1 vccd1 _18477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15431_ _18853_/Q _15363_/X _15430_/X vssd1 vssd1 vccd1 vccd1 _18853_/D sky130_fd_sc_hd__o21a_1
X_12643_ _12619_/X _12642_/X _12617_/B vssd1 vssd1 vccd1 vccd1 _12643_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16872__A _16918_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18150_ _17652_/X _19918_/Q _18158_/S vssd1 vssd1 vccd1 vccd1 _18151_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15362_ _18848_/Q _15278_/X _15361_/X vssd1 vssd1 vccd1 vccd1 _18848_/D sky130_fd_sc_hd__o21a_1
XFILLER_156_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12574_ _12574_/A _12574_/B vssd1 vssd1 vccd1 vccd1 _12574_/X sky130_fd_sc_hd__xor2_4
XFILLER_8_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17101_ _17097_/X _19490_/Q _17113_/S vssd1 vssd1 vccd1 vccd1 _17102_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11795__B1 _11794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14313_ _14316_/B _14314_/C _18670_/Q vssd1 vssd1 vccd1 vccd1 _14315_/B sky130_fd_sc_hd__a21oi_1
XFILLER_168_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11525_ _15976_/C _12862_/B vssd1 vssd1 vccd1 vccd1 _11643_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18081_ _18115_/A vssd1 vssd1 vccd1 vccd1 _18095_/S sky130_fd_sc_hd__buf_2
XANTENNA__16083__S _16089_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15293_ _15323_/A _15293_/B _15293_/C vssd1 vssd1 vccd1 vccd1 _15293_/X sky130_fd_sc_hd__and3_1
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17032_ _17032_/A vssd1 vssd1 vccd1 vccd1 _19464_/D sky130_fd_sc_hd__clkbuf_1
X_14244_ _14315_/A _14244_/B _14279_/C vssd1 vssd1 vccd1 vccd1 _18649_/D sky130_fd_sc_hd__nor3_1
XANTENNA__09486__A _15624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11456_ _15925_/C _12831_/B _12118_/A _12828_/B vssd1 vssd1 vccd1 vccd1 _11607_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10407_ _10508_/A _10407_/B vssd1 vssd1 vccd1 vccd1 _10407_/X sky130_fd_sc_hd__or2_1
XANTENNA__17907__S _17915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14175_ _14191_/A _14180_/C vssd1 vssd1 vccd1 vccd1 _14175_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16811__S _16819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ _19353_/Q _19688_/Q _11442_/S vssd1 vssd1 vccd1 vccd1 _11388_/B sky130_fd_sc_hd__mux2_1
XFILLER_125_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13126_ _18724_/Q vssd1 vssd1 vccd1 vccd1 _14476_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10338_ _09798_/A _10335_/X _10337_/X _09822_/A vssd1 vssd1 vccd1 vccd1 _10338_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_113_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _19523_/CLK _18983_/D vssd1 vssd1 vccd1 vccd1 _18983_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _17934_/A vssd1 vssd1 vccd1 vccd1 _19837_/D sky130_fd_sc_hd__clkbuf_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13057_/A vssd1 vssd1 vccd1 vccd1 _13120_/A sky130_fd_sc_hd__clkbuf_2
X_10269_ _20032_/Q _19870_/Q _19279_/Q _19049_/Q _10059_/S _10261_/X vssd1 vssd1 vccd1
+ vccd1 _10270_/B sky130_fd_sc_hd__mux4_1
XFILLER_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12008_ _12393_/A _12393_/B _12393_/C _12008_/D vssd1 vssd1 vccd1 vccd1 _12008_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17865_ _19807_/Q _17071_/X _17865_/S vssd1 vssd1 vccd1 vccd1 _17866_/A sky130_fd_sc_hd__mux2_1
X_19604_ _19828_/CLK _19604_/D vssd1 vssd1 vccd1 vccd1 _19604_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15951__A _15951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16816_ _16816_/A vssd1 vssd1 vccd1 vccd1 _19374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17796_ _17716_/X _19776_/Q _17804_/S vssd1 vssd1 vccd1 vccd1 _17797_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19535_ _19986_/CLK _19535_/D vssd1 vssd1 vccd1 vccd1 _19535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16747_ _19344_/Q _13835_/X _16747_/S vssd1 vssd1 vccd1 vccd1 _16748_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13959_ _13967_/A _13964_/C vssd1 vssd1 vccd1 vccd1 _13959_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16258__S _16258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19466_ _19990_/CLK _19466_/D vssd1 vssd1 vccd1 vccd1 _19466_/Q sky130_fd_sc_hd__dfxtp_1
X_16678_ _16678_/A vssd1 vssd1 vccd1 vccd1 _19313_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10381__S0 _10469_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18417_ _18417_/A vssd1 vssd1 vccd1 vccd1 _20037_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13190__B _13373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15629_ _18895_/Q _18927_/Q _15901_/S vssd1 vssd1 vccd1 vccd1 _15630_/A sky130_fd_sc_hd__mux2_1
X_19397_ _19985_/CLK _19397_/D vssd1 vssd1 vccd1 vccd1 _19397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10038__B1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18348_ _17732_/X _20007_/Q _18350_/S vssd1 vssd1 vccd1 vccd1 _18349_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10589__A1 _10822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10133__S0 _10449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18279_ _18279_/A vssd1 vssd1 vccd1 vccd1 _19976_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13527__A1 _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09396__A _18952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput50 io_ibus_inst[24] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_2
Xinput61 io_ibus_inst[5] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_8
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17817__S _17821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10335__A _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16721__S _16725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09983_ _19680_/Q _19446_/Q _18511_/Q _19776_/Q _09967_/X _09612_/A vssd1 vssd1 vccd1
+ vccd1 _09984_/B sky130_fd_sc_hd__mux4_1
XFILLER_103_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16022__A _16044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10513__A1 _09547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11710__B1 _14672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11166__A _11166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13381__A _13439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09417_ _18946_/Q _18945_/Q _18944_/Q _14225_/C vssd1 vssd1 vccd1 vccd1 _09417_/X
+ sky130_fd_sc_hd__or4_2
XANTENNA__13215__A0 _18848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18383__S _18385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_91_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09348_ _18833_/Q vssd1 vssd1 vccd1 vccd1 _12895_/A sky130_fd_sc_hd__clkinv_4
XFILLER_138_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09279_ _09434_/A _09285_/C _09435_/A _09436_/D vssd1 vssd1 vccd1 vccd1 _09279_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_154_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11310_ _19195_/Q _19786_/Q _19948_/Q _19163_/Q _11230_/X _11021_/A vssd1 vssd1 vccd1
+ vccd1 _11311_/B sky130_fd_sc_hd__mux4_1
XANTENNA__15101__A _15368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12290_ _18992_/Q _12290_/B _12315_/A vssd1 vssd1 vccd1 vccd1 _12290_/X sky130_fd_sc_hd__and3_1
XFILLER_147_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17727__S _17730_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11241_ _19133_/Q _19394_/Q _19293_/Q _19628_/Q _11156_/S _11108_/X vssd1 vssd1 vccd1
+ vccd1 _11242_/B sky130_fd_sc_hd__mux4_1
XANTENNA__15837__A2_N _15834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11172_ _11172_/A vssd1 vssd1 vccd1 vccd1 _11172_/X sky130_fd_sc_hd__buf_2
XFILLER_79_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ _10657_/S vssd1 vssd1 vccd1 vccd1 _10543_/S sky130_fd_sc_hd__clkbuf_2
X_15980_ _15982_/A _15980_/B vssd1 vssd1 vccd1 vccd1 _15980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A io_dbus_valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ _10054_/A vssd1 vssd1 vccd1 vccd1 _10054_/X sky130_fd_sc_hd__buf_2
XFILLER_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14931_ _14931_/A vssd1 vssd1 vccd1 vccd1 _15041_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_76_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17462__S _17470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17650_ _17649_/X _19723_/Q _17650_/S vssd1 vssd1 vccd1 vccd1 _17651_/A sky130_fd_sc_hd__mux2_1
X_14862_ _15291_/B _15424_/B _14915_/S vssd1 vssd1 vccd1 vccd1 _14862_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16601_ _16601_/A vssd1 vssd1 vccd1 vccd1 _19279_/D sky130_fd_sc_hd__clkbuf_1
X_13813_ _17049_/A vssd1 vssd1 vccd1 vccd1 _13813_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12257__A1 _12188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17581_ _17581_/A vssd1 vssd1 vccd1 vccd1 _19694_/D sky130_fd_sc_hd__clkbuf_1
X_14793_ _14789_/Y _14791_/Y _14795_/A vssd1 vssd1 vccd1 vccd1 _18829_/D sky130_fd_sc_hd__a21oi_1
X_16532_ _16532_/A vssd1 vssd1 vccd1 vccd1 _16541_/S sky130_fd_sc_hd__buf_4
X_19320_ _19816_/CLK _19320_/D vssd1 vssd1 vccd1 vccd1 _19320_/Q sky130_fd_sc_hd__dfxtp_1
X_13744_ _18484_/Q _13743_/X _13752_/S vssd1 vssd1 vccd1 vccd1 _13745_/A sky130_fd_sc_hd__mux2_1
X_10956_ _10856_/X _10953_/X _10955_/X vssd1 vssd1 vccd1 vccd1 _10956_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19251_ _20036_/CLK _19251_/D vssd1 vssd1 vccd1 vccd1 _19251_/Q sky130_fd_sc_hd__dfxtp_1
X_16463_ _16463_/A vssd1 vssd1 vccd1 vccd1 _19218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13675_ _19015_/Q _13675_/B vssd1 vssd1 vccd1 vccd1 _13675_/X sky130_fd_sc_hd__or2_1
XANTENNA__16806__S _16808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887_ _20019_/Q _19857_/Q _19266_/Q _19036_/Q _10776_/X _10596_/A vssd1 vssd1 vccd1
+ vccd1 _10887_/X sky130_fd_sc_hd__mux4_1
X_18202_ _17729_/X _19942_/Q _18202_/S vssd1 vssd1 vccd1 vccd1 _18203_/A sky130_fd_sc_hd__mux2_1
X_15414_ _15151_/X _15299_/X _15412_/X _15413_/X vssd1 vssd1 vccd1 vccd1 _15414_/X
+ sky130_fd_sc_hd__a211o_1
X_19182_ _19999_/CLK _19182_/D vssd1 vssd1 vccd1 vccd1 _19182_/Q sky130_fd_sc_hd__dfxtp_1
X_12626_ _18477_/Q _12722_/B vssd1 vssd1 vccd1 vccd1 _12626_/X sky130_fd_sc_hd__or2_1
X_16394_ _16393_/X _19189_/Q _16394_/S vssd1 vssd1 vccd1 vccd1 _16395_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18133_ _18864_/Q _12347_/A _16075_/B vssd1 vssd1 vccd1 vccd1 _18133_/X sky130_fd_sc_hd__a21o_1
XFILLER_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15345_ _18847_/Q _15278_/X _15344_/X vssd1 vssd1 vccd1 vccd1 _18847_/D sky130_fd_sc_hd__o21a_1
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _12557_/A vssd1 vssd1 vccd1 vccd1 _12557_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11661__A1_N _11667_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13509__A1 _13648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11508_ _15940_/C _12842_/A vssd1 vssd1 vccd1 vccd1 _11508_/Y sky130_fd_sc_hd__nor2_1
X_18064_ _18134_/S vssd1 vssd1 vccd1 vccd1 _18078_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_157_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15276_ _12273_/Y _15146_/X _15274_/X _15275_/X vssd1 vssd1 vccd1 vccd1 _15276_/X
+ sky130_fd_sc_hd__a211o_1
X_12488_ _12515_/A vssd1 vssd1 vccd1 vccd1 _12632_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17015_ _19459_/Q _17014_/X _17024_/S vssd1 vssd1 vccd1 vccd1 _17016_/A sky130_fd_sc_hd__mux2_1
X_14227_ _14227_/A _14227_/B _14227_/C _14227_/D vssd1 vssd1 vccd1 vccd1 _14227_/X
+ sky130_fd_sc_hd__or4_1
X_11439_ _19655_/Q _19421_/Q _18486_/Q _19751_/Q _11356_/X _11357_/X vssd1 vssd1 vccd1
+ vccd1 _11440_/B sky130_fd_sc_hd__mux4_1
XANTENNA__15946__A _15946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16541__S _16541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14158_ _18624_/Q _14154_/C _14157_/Y vssd1 vssd1 vccd1 vccd1 _18624_/D sky130_fd_sc_hd__o21a_1
XFILLER_113_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _18874_/Q vssd1 vssd1 vccd1 vccd1 _13110_/A sky130_fd_sc_hd__clkbuf_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14089_ _14089_/A vssd1 vssd1 vccd1 vccd1 _14095_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ _18992_/CLK _18966_/D vssd1 vssd1 vccd1 vccd1 _18966_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15682__A1 _18539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17917_ _17939_/A vssd1 vssd1 vccd1 vccd1 _17926_/S sky130_fd_sc_hd__clkbuf_4
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18897_ _18997_/CLK _18897_/D vssd1 vssd1 vccd1 vccd1 _18897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16777__A _16834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09361__A1 _18753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17372__S _17376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09361__B2 _18754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17848_ _19799_/Q _17046_/X _17854_/S vssd1 vssd1 vccd1 vccd1 _17849_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17779_ _17779_/A vssd1 vssd1 vccd1 vccd1 _19768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19518_ _19587_/CLK _19518_/D vssd1 vssd1 vccd1 vccd1 _19518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_113_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19449_ _19973_/CLK _19449_/D vssd1 vssd1 vccd1 vccd1 _19449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10274__A3 _10273_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09202_ _09256_/A vssd1 vssd1 vccd1 vccd1 _14761_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13748__A1 _19025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10764__S _10764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12420__A1 _18469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11223__A2 _09537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10431__B1 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12971__A2 _18836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16451__S _16457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18232__A _18278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10734__A1 _09686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_38_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _10180_/S vssd1 vssd1 vccd1 vccd1 _10313_/S sky130_fd_sc_hd__buf_2
XFILLER_104_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15673__A1 _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12487__A1 _12032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ _11554_/A _09897_/B vssd1 vssd1 vccd1 vccd1 _09897_/X sky130_fd_sc_hd__and2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15591__A _15602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14228__A2 _12918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _19332_/Q _19603_/Q _19827_/Q _19571_/Q _11486_/S _10625_/A vssd1 vssd1 vccd1
+ vccd1 _10810_/X sky130_fd_sc_hd__mux4_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11869_/A _11790_/B vssd1 vssd1 vccd1 vccd1 _11791_/A sky130_fd_sc_hd__nor2_2
XANTENNA__14000__A _14044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__S0 _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10741_ _09759_/A _10740_/X _09776_/A vssd1 vssd1 vccd1 vccd1 _10741_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16626__S _16630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13460_ _13460_/A _13460_/B vssd1 vssd1 vccd1 vccd1 _13460_/Y sky130_fd_sc_hd__nor2_1
X_10672_ _09987_/A _10671_/X _09563_/A vssd1 vssd1 vccd1 vccd1 _10672_/X sky130_fd_sc_hd__o21a_1
XANTENNA__18127__A0 _18862_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12411_ _12411_/A _14877_/A vssd1 vssd1 vccd1 vccd1 _12438_/A sky130_fd_sc_hd__xnor2_4
XFILLER_139_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13391_ _18891_/Q vssd1 vssd1 vccd1 vccd1 _13714_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15130_ _14932_/X _14891_/X _15199_/S vssd1 vssd1 vccd1 vccd1 _15130_/X sky130_fd_sc_hd__mux2_1
X_12342_ _12335_/A _12341_/X _12448_/S vssd1 vssd1 vccd1 vccd1 _12342_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17457__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15766__A _18952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15061_ _15056_/X _15059_/X _15280_/S vssd1 vssd1 vccd1 vccd1 _15061_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12273_ _12273_/A vssd1 vssd1 vccd1 vccd1 _12273_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14012_ _14507_/A vssd1 vssd1 vccd1 vccd1 _14046_/A sky130_fd_sc_hd__buf_2
X_11224_ _19918_/Q _19532_/Q _19982_/Q _19101_/Q _11171_/X _09737_/A vssd1 vssd1 vccd1
+ vccd1 _11225_/B sky130_fd_sc_hd__mux4_1
XFILLER_122_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18820_ _19912_/CLK _18820_/D vssd1 vssd1 vccd1 vccd1 _18820_/Q sky130_fd_sc_hd__dfxtp_1
X_11155_ _11155_/A vssd1 vssd1 vccd1 vccd1 _11156_/S sky130_fd_sc_hd__buf_4
XANTENNA__10703__A _10703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15664__A1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ _10047_/Y _10104_/Y _10248_/A vssd1 vssd1 vccd1 vccd1 _10106_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18751_ _19062_/CLK _18751_/D vssd1 vssd1 vccd1 vccd1 _18751_/Q sky130_fd_sc_hd__dfxtp_1
X_15963_ _19015_/Q _15951_/X _15962_/X vssd1 vssd1 vccd1 vccd1 _19015_/D sky130_fd_sc_hd__a21o_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11086_ _11086_/A vssd1 vssd1 vccd1 vccd1 _11296_/A sky130_fd_sc_hd__buf_2
XFILLER_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17702_ _17700_/X _19739_/Q _17714_/S vssd1 vssd1 vccd1 vccd1 _17703_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10489__B1 _09913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ _19377_/Q _19712_/Q _10037_/S vssd1 vssd1 vccd1 vccd1 _10037_/X sky130_fd_sc_hd__mux2_1
X_14914_ _14914_/A vssd1 vssd1 vccd1 vccd1 _15138_/B sky130_fd_sc_hd__buf_2
X_15894_ _15897_/A _15894_/B vssd1 vssd1 vccd1 vccd1 _15895_/A sky130_fd_sc_hd__and2_1
X_18682_ _19882_/CLK _18682_/D vssd1 vssd1 vccd1 vccd1 _18682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15416__B2 _12521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17633_ _17633_/A vssd1 vssd1 vccd1 vccd1 _19718_/D sky130_fd_sc_hd__clkbuf_1
X_14845_ _15384_/A vssd1 vssd1 vccd1 vccd1 _15142_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15967__A2 _15951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17920__S _17926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14776_ _14780_/A _14776_/B vssd1 vssd1 vccd1 vccd1 _14777_/A sky130_fd_sc_hd__and2_1
X_17564_ _17632_/S vssd1 vssd1 vccd1 vccd1 _17573_/S sky130_fd_sc_hd__buf_2
XANTENNA__10336__S0 _10152_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11989__A0 _11452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11988_ _11988_/A _15094_/A vssd1 vssd1 vccd1 vccd1 _12044_/A sky130_fd_sc_hd__xnor2_2
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19303_ _19767_/CLK _19303_/D vssd1 vssd1 vccd1 vccd1 _19303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16515_ _19241_/Q _13813_/X _16519_/S vssd1 vssd1 vccd1 vccd1 _16516_/A sky130_fd_sc_hd__mux2_1
X_13727_ _11813_/X _13725_/X _13726_/Y _11831_/X _19022_/Q vssd1 vssd1 vccd1 vccd1
+ _13727_/X sky130_fd_sc_hd__a32o_2
X_10939_ _10712_/A _10932_/Y _10934_/Y _10936_/Y _10938_/Y vssd1 vssd1 vccd1 vccd1
+ _10939_/X sky130_fd_sc_hd__o32a_1
XANTENNA__10887__S1 _10596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17495_ _17495_/A vssd1 vssd1 vccd1 vccd1 _19653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19234_ _19827_/CLK _19234_/D vssd1 vssd1 vccd1 vccd1 _19234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16446_ _19211_/Q _13819_/X _16446_/S vssd1 vssd1 vccd1 vccd1 _16447_/A sky130_fd_sc_hd__mux2_1
X_13658_ _14552_/A vssd1 vssd1 vccd1 vccd1 _13732_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18118__A0 _18859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12609_ _12515_/A _15449_/A _12591_/A vssd1 vssd1 vccd1 vccd1 _12613_/A sky130_fd_sc_hd__a21o_1
X_16377_ _17713_/A vssd1 vssd1 vccd1 vccd1 _16377_/X sky130_fd_sc_hd__clkbuf_2
X_19165_ _19758_/CLK _19165_/D vssd1 vssd1 vccd1 vccd1 _19165_/Q sky130_fd_sc_hd__dfxtp_1
X_13589_ _13589_/A _19004_/Q vssd1 vssd1 vccd1 vccd1 _13589_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15328_ _18846_/Q _15278_/X _15327_/X vssd1 vssd1 vccd1 vccd1 _18846_/D sky130_fd_sc_hd__o21a_1
X_18116_ _18114_/X _19906_/Q _18128_/S vssd1 vssd1 vccd1 vccd1 _18117_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12953__A2 _11732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19096_ _19978_/CLK _19096_/D vssd1 vssd1 vccd1 vccd1 _19096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18047_ _18134_/S vssd1 vssd1 vccd1 vccd1 _18061_/S sky130_fd_sc_hd__clkbuf_2
X_15259_ _15243_/X _15246_/X _15257_/X _15258_/X vssd1 vssd1 vccd1 vccd1 _15259_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14580__A _14648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09674__A _10069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13902__A1 _18542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ _09820_/A vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__buf_2
XFILLER_101_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19998_ _19998_/CLK _19998_/D vssd1 vssd1 vccd1 vccd1 _19998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09751_ _19386_/Q vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__inv_2
X_18949_ _18956_/CLK _18949_/D vssd1 vssd1 vccd1 vccd1 _18949_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18198__S _18202_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09682_ _09682_/A vssd1 vssd1 vccd1 vccd1 _09683_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17830__S _17832_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16446__S _16446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17131__A _17668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09849__A _09849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10955__A1 _11237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11055__S1 _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12722__B _12722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09949_ _09942_/Y _09944_/Y _09946_/Y _09948_/Y _11574_/A vssd1 vssd1 vccd1 vccd1
+ _09949_/X sky130_fd_sc_hd__o221a_1
XFILLER_131_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10242__B _12858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17306__A _17352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12960_ _12960_/A _13504_/A vssd1 vssd1 vccd1 vccd1 _12960_/Y sky130_fd_sc_hd__nand2_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11911_ _12196_/A vssd1 vssd1 vccd1 vccd1 _12472_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13409__B1 _13368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ _18646_/Q _12889_/X _12890_/X _18714_/Q vssd1 vssd1 vccd1 vccd1 _12891_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14630_/A vssd1 vssd1 vccd1 vccd1 _18777_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10891__B1 _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11842_ _12984_/A vssd1 vssd1 vccd1 vccd1 _12879_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _18995_/Q _12933_/X _14560_/Y _11717_/X vssd1 vssd1 vccd1 vccd1 _14561_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11773_ _11773_/A vssd1 vssd1 vccd1 vccd1 _11860_/B sky130_fd_sc_hd__inv_2
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16356__S _16362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14665__A _14665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18137__A _18193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16300_ _16381_/A vssd1 vssd1 vccd1 vccd1 _16400_/S sky130_fd_sc_hd__buf_6
X_13512_ _19489_/Q _14792_/B _13511_/X _11915_/B vssd1 vssd1 vccd1 vccd1 _13520_/A
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _19366_/Q _19701_/Q _10724_/S vssd1 vssd1 vccd1 vccd1 _10724_/X sky130_fd_sc_hd__mux2_1
X_17280_ _17198_/X _19558_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17281_/A sky130_fd_sc_hd__mux2_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14492_ _14493_/B _14493_/C _14491_/Y vssd1 vssd1 vccd1 vccd1 _18730_/D sky130_fd_sc_hd__o21a_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14384__B _18690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16231_ _16231_/A vssd1 vssd1 vccd1 vccd1 _19129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13443_ _17726_/A vssd1 vssd1 vccd1 vccd1 _13443_/X sky130_fd_sc_hd__clkbuf_2
X_10655_ _19367_/Q _19702_/Q _10655_/S vssd1 vssd1 vccd1 vccd1 _10656_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12935__A2 _12933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16162_ _13002_/X _19100_/Q _16162_/S vssd1 vssd1 vccd1 vccd1 _16163_/A sky130_fd_sc_hd__mux2_1
X_13374_ _18479_/Q _12943_/X _12944_/X _18703_/Q _13373_/X vssd1 vssd1 vccd1 vccd1
+ _13374_/X sky130_fd_sc_hd__a221o_1
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10586_ _19368_/Q _19703_/Q _10586_/S vssd1 vssd1 vccd1 vccd1 _10587_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15113_ _15023_/X _15018_/X _15113_/S vssd1 vssd1 vccd1 vccd1 _15113_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17187__S _17193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12325_ _15306_/A _12325_/B vssd1 vssd1 vccd1 vccd1 _12328_/B sky130_fd_sc_hd__xor2_1
X_16093_ _16093_/A vssd1 vssd1 vccd1 vccd1 _19069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19921_ _19985_/CLK _19921_/D vssd1 vssd1 vccd1 vccd1 _19921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15044_ _15035_/X _15043_/X _15100_/A vssd1 vssd1 vccd1 vccd1 _15044_/X sky130_fd_sc_hd__mux2_1
X_12256_ _12344_/A _12254_/Y _12309_/C _12366_/B vssd1 vssd1 vccd1 vccd1 _12256_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_135_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12699__A1 _12338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11046__S1 _11045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17915__S _17915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ _11322_/A vssd1 vssd1 vccd1 vccd1 _11208_/A sky130_fd_sc_hd__clkbuf_4
X_19852_ _19949_/CLK _19852_/D vssd1 vssd1 vccd1 vccd1 _19852_/Q sky130_fd_sc_hd__dfxtp_1
X_12187_ _18525_/Q _12303_/B vssd1 vssd1 vccd1 vccd1 _12204_/A sky130_fd_sc_hd__or2_1
XFILLER_69_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18803_ _19883_/CLK _18803_/D vssd1 vssd1 vccd1 vccd1 _18803_/Q sky130_fd_sc_hd__dfxtp_1
X_11138_ _20015_/Q _19853_/Q _19262_/Q _19032_/Q _10995_/X _10996_/X vssd1 vssd1 vccd1
+ vccd1 _11138_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15943__B _15943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19783_ _19947_/CLK _19783_/D vssd1 vssd1 vccd1 vccd1 _19783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16995_ _17094_/S vssd1 vssd1 vccd1 vccd1 _17008_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18734_ _18734_/CLK _18734_/D vssd1 vssd1 vccd1 vccd1 _18734_/Q sky130_fd_sc_hd__dfxtp_1
X_11069_ _11335_/A vssd1 vssd1 vccd1 vccd1 _11332_/A sky130_fd_sc_hd__clkbuf_2
X_15946_ _15946_/A vssd1 vssd1 vccd1 vccd1 _15966_/B sky130_fd_sc_hd__buf_2
XFILLER_95_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18665_ _19683_/CLK _18665_/D vssd1 vssd1 vccd1 vccd1 _18665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15877_ _15881_/A _15877_/B vssd1 vssd1 vccd1 vccd1 _15878_/A sky130_fd_sc_hd__and2_1
XFILLER_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17650__S _17650_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17616_ _17616_/A vssd1 vssd1 vccd1 vccd1 _19710_/D sky130_fd_sc_hd__clkbuf_1
X_14828_ _14973_/A _15004_/B _14955_/S vssd1 vssd1 vccd1 vccd1 _15546_/A sky130_fd_sc_hd__or3b_1
X_18596_ _19683_/CLK _18596_/D vssd1 vssd1 vccd1 vccd1 _18596_/Q sky130_fd_sc_hd__dfxtp_1
X_17547_ _17547_/A vssd1 vssd1 vccd1 vccd1 _19679_/D sky130_fd_sc_hd__clkbuf_1
X_14759_ _15393_/A vssd1 vssd1 vccd1 vccd1 _15539_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17478_ _17478_/A vssd1 vssd1 vccd1 vccd1 _19645_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12807__B _12807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19217_ _20002_/CLK _19217_/D vssd1 vssd1 vccd1 vccd1 _19217_/Q sky130_fd_sc_hd__dfxtp_1
X_16429_ _19203_/Q _13794_/X _16435_/S vssd1 vssd1 vccd1 vccd1 _16430_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10608__A _10836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19148_ _19965_/CLK _19148_/D vssd1 vssd1 vccd1 vccd1 _19148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19079_ _20026_/CLK _19079_/D vssd1 vssd1 vccd1 vccd1 _19079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12823__A _15899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15876__A1 _09261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15876__B2 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13887__B1 _14447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09803_ _09803_/A vssd1 vssd1 vccd1 vccd1 _09804_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__13639__A0 _11724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10570__C1 _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _19385_/Q vssd1 vssd1 vccd1 vccd1 _11019_/A sky130_fd_sc_hd__buf_2
XANTENNA__13654__A _18884_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09665_ _10822_/A vssd1 vssd1 vccd1 vccd1 _10448_/A sky130_fd_sc_hd__buf_2
XANTENNA__13373__B _13373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11174__A _11227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09596_ _10251_/S vssd1 vssd1 vccd1 vccd1 _09597_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16176__S _16184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11902__A _12831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09579__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _10392_/A _10439_/X _10159_/X vssd1 vssd1 vccd1 vccd1 _10440_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13829__A _17065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _10365_/A _10370_/X _09980_/A vssd1 vssd1 vccd1 vccd1 _10371_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12733__A _12753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15867__A1 _09454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12110_ _12134_/B _12168_/S _13595_/A vssd1 vssd1 vccd1 vccd1 _12110_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__15867__B2 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13090_ _13068_/X _13085_/X _13089_/X vssd1 vssd1 vccd1 vccd1 _13090_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__11028__S1 _11157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12041_ _12042_/A _14895_/A vssd1 vssd1 vccd1 vccd1 _12043_/A sky130_fd_sc_hd__and2_1
XFILLER_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11353__A1 _11344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15800_ _15813_/A _15800_/B vssd1 vssd1 vccd1 vccd1 _15801_/A sky130_fd_sc_hd__and2_1
XANTENNA__17036__A _17036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16780_ _16320_/X _19358_/Q _16786_/S vssd1 vssd1 vccd1 vccd1 _16781_/A sky130_fd_sc_hd__mux2_1
X_13992_ _18572_/Q _13992_/B vssd1 vssd1 vccd1 vccd1 _13999_/C sky130_fd_sc_hd__and2_1
XFILLER_19_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15731_ _18970_/Q _15720_/X _15729_/X _15730_/X vssd1 vssd1 vccd1 vccd1 _18938_/D
+ sky130_fd_sc_hd__o211a_1
X_12943_ _12943_/A vssd1 vssd1 vccd1 vccd1 _12943_/X sky130_fd_sc_hd__buf_2
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17241__A0 _17141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17470__S _17470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11084__A _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _19942_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _13223_/A vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__buf_4
X_15662_ _18909_/Q _12340_/B _15666_/S vssd1 vssd1 vccd1 vccd1 _15663_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _19611_/Q _17058_/X _17409_/S vssd1 vssd1 vccd1 vccd1 _17402_/A sky130_fd_sc_hd__mux2_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _14613_/A vssd1 vssd1 vccd1 vccd1 _18772_/D sky130_fd_sc_hd__clkbuf_1
X_11825_ _18593_/Q _11851_/A _12887_/A _18625_/Q vssd1 vssd1 vccd1 vccd1 _11825_/X
+ sky130_fd_sc_hd__a22o_1
X_18381_ _17675_/X _20021_/Q _18385_/S vssd1 vssd1 vccd1 vccd1 _18382_/A sky130_fd_sc_hd__mux2_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output102_A _12246_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15593_ _15593_/A vssd1 vssd1 vccd1 vccd1 _18878_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12908__A _16992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _17332_/A vssd1 vssd1 vccd1 vccd1 _19580_/D sky130_fd_sc_hd__clkbuf_1
X_14544_ input69/X _14544_/B vssd1 vssd1 vccd1 vccd1 _14544_/X sky130_fd_sc_hd__or2_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _18752_/Q _14547_/A _13451_/B _19899_/Q vssd1 vssd1 vccd1 vccd1 _11756_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _10775_/A vssd1 vssd1 vccd1 vccd1 _10919_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_159_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17263_ _17173_/X _19550_/Q _17265_/S vssd1 vssd1 vccd1 vccd1 _17264_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14475_ _14476_/B _14476_/C _14474_/Y vssd1 vssd1 vccd1 vccd1 _18724_/D sky130_fd_sc_hd__o21a_1
XFILLER_174_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11687_ _11824_/A vssd1 vssd1 vccd1 vccd1 _11687_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11023__S _11023_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19002_ _19025_/CLK _19002_/D vssd1 vssd1 vccd1 vccd1 _19002_/Q sky130_fd_sc_hd__dfxtp_2
X_16214_ _16214_/A vssd1 vssd1 vccd1 vccd1 _19123_/D sky130_fd_sc_hd__clkbuf_1
X_13426_ input21/X _13318_/X _13368_/X vssd1 vssd1 vccd1 vccd1 _13426_/Y sky130_fd_sc_hd__a21oi_1
X_10638_ _10638_/A vssd1 vssd1 vccd1 vccd1 _10638_/X sky130_fd_sc_hd__buf_2
X_17194_ _17194_/A vssd1 vssd1 vccd1 vccd1 _19519_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13030__A1 _18460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15938__B _15955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16145_ _16145_/A vssd1 vssd1 vccd1 vccd1 _19093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13357_ _18888_/Q _18889_/Q _13357_/C vssd1 vssd1 vccd1 vccd1 _13390_/C sky130_fd_sc_hd__and3_1
X_10569_ _10572_/A _10568_/X _09796_/A vssd1 vssd1 vccd1 vccd1 _10569_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19562_/CLK sky130_fd_sc_hd__clkbuf_16
X_12308_ _12283_/A _12309_/C _18768_/Q vssd1 vssd1 vccd1 vccd1 _12308_/Y sky130_fd_sc_hd__a21oi_1
X_16076_ _19063_/Q _16075_/X _16076_/S vssd1 vssd1 vccd1 vccd1 _16077_/A sky130_fd_sc_hd__mux2_1
X_13288_ _18885_/Q _13288_/B vssd1 vssd1 vccd1 vccd1 _13326_/C sky130_fd_sc_hd__and2_1
XANTENNA__13458__B _13731_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15027_ _15017_/X _15025_/X _15190_/S vssd1 vssd1 vccd1 vccd1 _15027_/X sky130_fd_sc_hd__mux2_1
X_19904_ _19910_/CLK _19904_/D vssd1 vssd1 vccd1 vccd1 _19904_/Q sky130_fd_sc_hd__dfxtp_1
X_12239_ _12239_/A vssd1 vssd1 vccd1 vccd1 _12239_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15954__A _15954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13333__A2 _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10163__A _10473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19835_ _19965_/CLK _19835_/D vssd1 vssd1 vccd1 vccd1 _19835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15086__A2 _15078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19766_ _19767_/CLK _19766_/D vssd1 vssd1 vccd1 vccd1 _19766_/Q sky130_fd_sc_hd__dfxtp_1
X_16978_ _16380_/X _19446_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16979_/A sky130_fd_sc_hd__mux2_1
Xinput4 io_dbus_rdata[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
XFILLER_77_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18717_ _18744_/CLK _18717_/D vssd1 vssd1 vccd1 vccd1 _18717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15929_ _15942_/A vssd1 vssd1 vccd1 vccd1 _15936_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19697_ _19827_/CLK _19697_/D vssd1 vssd1 vccd1 vccd1 _19697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09450_ _11983_/S vssd1 vssd1 vccd1 vccd1 _12033_/S sky130_fd_sc_hd__clkbuf_2
X_18648_ _18688_/CLK _18648_/D vssd1 vssd1 vccd1 vccd1 _18648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09381_ _13510_/A vssd1 vssd1 vccd1 vccd1 _09381_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18579_ _18819_/CLK _18579_/D vssd1 vssd1 vccd1 vccd1 _18579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14349__A1 _14350_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__B1 _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13021__B2 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10073__A _10073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10769__S0 _10921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09862__A _09862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11430__S1 _11357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13384__A _17074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09717_ _19384_/Q vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__buf_2
XFILLER_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09648_ _10921_/S vssd1 vssd1 vccd1 vccd1 _10872_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14588__A1 _13572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _10458_/A vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__buf_2
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_161_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11610_ _11967_/A _11450_/X _11408_/X vssd1 vssd1 vccd1 vccd1 _11610_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _09454_/B _12657_/A _12682_/A _12589_/Y vssd1 vssd1 vccd1 vccd1 _15449_/A
+ sky130_fd_sc_hd__a211o_4
XANTENNA__13260__A1 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11497__S1 _10856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11541_ _09690_/X _11536_/X _11538_/Y _11540_/Y _09876_/X vssd1 vssd1 vccd1 vccd1
+ _11541_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11271__B1 _11425_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14260_ _14279_/B _14264_/D _14259_/Y vssd1 vssd1 vccd1 vccd1 _18654_/D sky130_fd_sc_hd__o21a_1
XFILLER_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11472_ _19141_/Q _19402_/Q _19301_/Q _19636_/Q _10776_/X _10596_/A vssd1 vssd1 vccd1
+ vccd1 _11473_/B sky130_fd_sc_hd__mux4_1
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11249__S1 _11208_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ _18805_/Q _12880_/X _11817_/X _18772_/Q _13210_/X vssd1 vssd1 vccd1 vccd1
+ _13211_/X sky130_fd_sc_hd__a221o_4
X_10423_ _19244_/Q _19739_/Q _10470_/S vssd1 vssd1 vccd1 vccd1 _10424_/B sky130_fd_sc_hd__mux2_1
X_14191_ _14191_/A _14197_/C vssd1 vssd1 vccd1 vccd1 _14191_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12771__B1 _13648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13142_ _13603_/A _13143_/B _13359_/B vssd1 vssd1 vccd1 vccd1 _13142_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_input63_A io_ibus_inst[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ _19245_/Q _19740_/Q _10354_/S vssd1 vssd1 vccd1 vccd1 _10355_/B sky130_fd_sc_hd__mux2_1
XFILLER_125_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13315__A2 _13120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17950_ _19845_/Q _17090_/X _17952_/S vssd1 vssd1 vccd1 vccd1 _17951_/A sky130_fd_sc_hd__mux2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _18462_/Q _11740_/X _12881_/A _14371_/B vssd1 vssd1 vccd1 vccd1 _13073_/X
+ sky130_fd_sc_hd__a22o_1
X_10285_ _10292_/A _10285_/B vssd1 vssd1 vccd1 vccd1 _10285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16901_ _16374_/X _19412_/Q _16903_/S vssd1 vssd1 vccd1 vccd1 _16902_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12024_ _12011_/X _12014_/Y _12021_/Y _12023_/X vssd1 vssd1 vccd1 vccd1 _12024_/Y
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__09772__A _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17881_ _17881_/A vssd1 vssd1 vccd1 vccd1 _19814_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17462__A0 _17147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12910__B _17098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19620_ _20039_/CLK _19620_/D vssd1 vssd1 vccd1 vccd1 _19620_/Q sky130_fd_sc_hd__dfxtp_1
X_16832_ _16396_/X _19382_/Q _16834_/S vssd1 vssd1 vccd1 vccd1 _16833_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19551_ _19583_/CLK _19551_/D vssd1 vssd1 vccd1 vccd1 _19551_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11526__B _12863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16763_ _16763_/A vssd1 vssd1 vccd1 vccd1 _19351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13975_ _14507_/A vssd1 vssd1 vccd1 vccd1 _14010_/A sky130_fd_sc_hd__buf_2
XANTENNA__18296__S _18302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18502_ _19767_/CLK _18502_/D vssd1 vssd1 vccd1 vccd1 _18502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15714_ _09481_/A _15705_/X _15712_/X _15713_/X vssd1 vssd1 vccd1 vccd1 _18932_/D
+ sky130_fd_sc_hd__o211a_1
X_19482_ _19876_/CLK _19482_/D vssd1 vssd1 vccd1 vccd1 _19482_/Q sky130_fd_sc_hd__dfxtp_1
X_12926_ _19882_/Q _13431_/B vssd1 vssd1 vccd1 vccd1 _12926_/X sky130_fd_sc_hd__and2_1
X_16694_ _16762_/S vssd1 vssd1 vccd1 vccd1 _16703_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__15940__C _15940_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18433_ _19824_/CLK _18433_/D vssd1 vssd1 vccd1 vccd1 _18433_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ _15645_/A vssd1 vssd1 vccd1 vccd1 _18901_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12857_ _12857_/A _12857_/B vssd1 vssd1 vccd1 vccd1 _12857_/Y sky130_fd_sc_hd__nor2_8
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11808_ _18710_/Q vssd1 vssd1 vccd1 vccd1 _12060_/B sky130_fd_sc_hd__clkbuf_4
X_18364_ _18364_/A vssd1 vssd1 vccd1 vccd1 _20013_/D sky130_fd_sc_hd__clkbuf_1
X_15576_ _13046_/A _18903_/Q _15578_/S vssd1 vssd1 vccd1 vccd1 _15577_/A sky130_fd_sc_hd__mux2_1
X_12788_ _12788_/A _12788_/B vssd1 vssd1 vccd1 vccd1 _12789_/B sky130_fd_sc_hd__nand2_2
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17144_/X _19573_/Q _17315_/S vssd1 vssd1 vccd1 vccd1 _17316_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15949__A _15964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11739_ _18753_/Q _14547_/A _13451_/B _19898_/Q vssd1 vssd1 vccd1 vccd1 _11743_/A
+ sky130_fd_sc_hd__a22o_1
X_14527_ _14526_/B _14526_/C _18743_/Q vssd1 vssd1 vccd1 vccd1 _14528_/C sky130_fd_sc_hd__a21oi_1
XFILLER_30_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18295_ _18295_/A vssd1 vssd1 vccd1 vccd1 _19982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17246_ _17147_/X _19542_/Q _17254_/S vssd1 vssd1 vccd1 vccd1 _17247_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14458_ _15715_/B vssd1 vssd1 vccd1 vccd1 _14495_/A sky130_fd_sc_hd__clkbuf_4
X_13409_ input20/X _13318_/X _13368_/X vssd1 vssd1 vccd1 vccd1 _13409_/Y sky130_fd_sc_hd__a21oi_1
X_17177_ _17176_/X _19514_/Q _17177_/S vssd1 vssd1 vccd1 vccd1 _17178_/A sky130_fd_sc_hd__mux2_1
X_14389_ _14390_/A _14390_/B _14388_/X vssd1 vssd1 vccd1 vccd1 _18692_/D sky130_fd_sc_hd__a21oi_1
XFILLER_155_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_152_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19882_/CLK sky130_fd_sc_hd__clkbuf_16
X_16128_ _16128_/A vssd1 vssd1 vccd1 vccd1 _19085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16059_ _11915_/B _12878_/X _13511_/C _14745_/B vssd1 vssd1 vccd1 vccd1 _16076_/S
+ sky130_fd_sc_hd__a31o_1
XFILLER_142_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09682__A _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__C1 _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11868__A2 _14159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_167_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _18867_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17453__A0 _17135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19818_ _19947_/CLK _19818_/D vssd1 vssd1 vccd1 vccd1 _19818_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11717__A _11730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10621__A _10907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19749_ _19974_/CLK _19749_/D vssd1 vssd1 vccd1 vccd1 _19749_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16719__S _16725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09502_ _09502_/A _09516_/A vssd1 vssd1 vccd1 vccd1 _14804_/C sky130_fd_sc_hd__nor2_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12293__A2 _12839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09694__B1 _09547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10923__S0 _10703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09433_ _15457_/A vssd1 vssd1 vccd1 vccd1 _09433_/X sky130_fd_sc_hd__buf_2
XFILLER_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11452__A _11452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _12062_/A vssd1 vssd1 vccd1 vccd1 _12064_/B sky130_fd_sc_hd__inv_2
XFILLER_36_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_105_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19583_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09295_ _18980_/Q _18940_/Q vssd1 vssd1 vccd1 vccd1 _09295_/X sky130_fd_sc_hd__xor2_1
XANTENNA__14763__A _14782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14742__A1 _13750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17692__A0 _17691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17285__S _17293_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16495__A1 _13784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_108_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput160 _12703_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[26] sky130_fd_sc_hd__buf_2
XFILLER_88_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput171 _12205_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_121_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10070_ _18448_/Q _19477_/Q _19514_/Q _19088_/Q _09597_/A _10054_/X vssd1 vssd1 vccd1
+ vccd1 _10070_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11403__S1 _19385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09921__A1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13842__A _17078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13760_ _18486_/Q _13754_/X _13772_/S vssd1 vssd1 vccd1 vccd1 _13761_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10972_ _10972_/A vssd1 vssd1 vccd1 vccd1 _10973_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ _12713_/B vssd1 vssd1 vccd1 vccd1 _15509_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13691_ _18477_/Q _13689_/X _13752_/S vssd1 vssd1 vccd1 vccd1 _13692_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15430_ _12551_/Y _15364_/X _15429_/X _15360_/X vssd1 vssd1 vccd1 vccd1 _15430_/X
+ sky130_fd_sc_hd__a211o_1
X_12642_ _12642_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _12642_/X sky130_fd_sc_hd__or2b_1
XANTENNA__12036__A2 _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_opt_6_0_clock _18998_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_6_0_clock/X sky130_fd_sc_hd__clkbuf_16
XFILLER_157_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15361_ _12413_/Y _15279_/X _15359_/X _15360_/X vssd1 vssd1 vccd1 vccd1 _15361_/X
+ sky130_fd_sc_hd__a211o_1
X_12573_ _12550_/A _12550_/B _12545_/A vssd1 vssd1 vccd1 vccd1 _12574_/B sky130_fd_sc_hd__a21bo_1
XFILLER_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17100_ _17199_/S vssd1 vssd1 vccd1 vccd1 _17113_/S sky130_fd_sc_hd__buf_4
XANTENNA__09767__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ _11524_/A _11634_/A _11634_/B _11642_/B vssd1 vssd1 vccd1 vccd1 _11524_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_12_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14312_ _18668_/Q _18667_/Q _14312_/C vssd1 vssd1 vccd1 vccd1 _14314_/C sky130_fd_sc_hd__and3_2
X_18080_ _18848_/Q _13629_/X _18084_/S vssd1 vssd1 vccd1 vccd1 _18080_/X sky130_fd_sc_hd__mux2_1
X_15292_ _15218_/X _15285_/Y _15291_/Y vssd1 vssd1 vccd1 vccd1 _15293_/C sky130_fd_sc_hd__a21oi_1
X_17031_ _19464_/Q _17030_/X _17040_/S vssd1 vssd1 vccd1 vccd1 _17032_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13289__A _13289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14243_ _14256_/C vssd1 vssd1 vccd1 vccd1 _14279_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_156_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11455_ _11608_/B _11453_/X _11454_/Y vssd1 vssd1 vccd1 vccd1 _11455_/X sky130_fd_sc_hd__a21o_1
X_10406_ _19148_/Q _19409_/Q _19308_/Q _19643_/Q _10129_/S _10398_/A vssd1 vssd1 vccd1
+ vccd1 _10407_/B sky130_fd_sc_hd__mux4_1
XFILLER_125_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14174_ _18630_/Q _14174_/B vssd1 vssd1 vccd1 vccd1 _14180_/C sky130_fd_sc_hd__and2_1
XFILLER_164_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ _09544_/A _11375_/X _11384_/X _10078_/A _12934_/A vssd1 vssd1 vccd1 vccd1
+ _11960_/A sky130_fd_sc_hd__o32a_1
XFILLER_125_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13125_ _18656_/Q _12889_/A _12887_/A _18624_/Q vssd1 vssd1 vccd1 vccd1 _13125_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_84_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 _19771_/CLK sky130_fd_sc_hd__clkbuf_16
X_10337_ _10434_/A _10337_/B vssd1 vssd1 vccd1 vccd1 _10337_/X sky130_fd_sc_hd__or2_1
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18982_ _19523_/CLK _18982_/D vssd1 vssd1 vccd1 vccd1 _18982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17933_ _19837_/Q _17065_/X _17937_/S vssd1 vssd1 vccd1 vccd1 _17934_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _18589_/Q vssd1 vssd1 vccd1 vccd1 _14042_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10268_ _10064_/X _10267_/X _09567_/A vssd1 vssd1 vccd1 vccd1 _10268_/X sky130_fd_sc_hd__o21a_1
XFILLER_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12007_ _12052_/B _12007_/B vssd1 vssd1 vccd1 vccd1 _12008_/D sky130_fd_sc_hd__or2_1
X_17864_ _17864_/A vssd1 vssd1 vccd1 vccd1 _19806_/D sky130_fd_sc_hd__clkbuf_1
X_10199_ _20035_/Q _19873_/Q _19282_/Q _19052_/Q _10313_/S _10182_/X vssd1 vssd1 vccd1
+ vccd1 _10200_/B sky130_fd_sc_hd__mux4_1
XFILLER_94_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_99_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19868_/CLK sky130_fd_sc_hd__clkbuf_16
X_19603_ _20025_/CLK _19603_/D vssd1 vssd1 vccd1 vccd1 _19603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16815_ _16371_/X _19374_/Q _16819_/S vssd1 vssd1 vccd1 vccd1 _16816_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17795_ _17795_/A vssd1 vssd1 vccd1 vccd1 _17804_/S sky130_fd_sc_hd__buf_4
XANTENNA__16539__S _16541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19534_ _19982_/CLK _19534_/D vssd1 vssd1 vccd1 vccd1 _19534_/Q sky130_fd_sc_hd__dfxtp_1
X_16746_ _16746_/A vssd1 vssd1 vccd1 vccd1 _19343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13958_ _18560_/Q _18559_/Q _18558_/Q _13958_/D vssd1 vssd1 vccd1 vccd1 _13964_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19465_ _19633_/CLK _19465_/D vssd1 vssd1 vccd1 vccd1 _19465_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_22_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19792_/CLK sky130_fd_sc_hd__clkbuf_16
X_12909_ _17634_/A vssd1 vssd1 vccd1 vccd1 _12909_/X sky130_fd_sc_hd__clkbuf_2
X_16677_ _16380_/X _19313_/Q _16685_/S vssd1 vssd1 vccd1 vccd1 _16678_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12368__A _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13889_ _12416_/C _13883_/X _12421_/Y _12426_/Y _13885_/X vssd1 vssd1 vccd1 vccd1
+ _18533_/D sky130_fd_sc_hd__o221a_1
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10381__S1 _10163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18416_ _17726_/X _20037_/Q _18418_/S vssd1 vssd1 vccd1 vccd1 _18417_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15628_ _15628_/A vssd1 vssd1 vccd1 vccd1 _18894_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19396_ _19758_/CLK _19396_/D vssd1 vssd1 vccd1 vccd1 _19396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10038__A1 _10028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18347_ _18347_/A vssd1 vssd1 vccd1 vccd1 _20006_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15679__A _15690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16274__S _16280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15559_ _15074_/X _15346_/Y _15243_/A vssd1 vssd1 vccd1 vccd1 _15559_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_37_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19731_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11786__B2 _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12983__B1 _13511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18278_ _19976_/Q _17735_/A _18278_/S vssd1 vssd1 vccd1 vccd1 _18279_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 io_ibus_inst[15] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__13527__A2 _13517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17229_ _17229_/A vssd1 vssd1 vccd1 vccd1 _19534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09396__B _18951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10616__A _15949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput51 io_ibus_inst[25] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_2
Xinput62 io_ibus_inst[6] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10746__C1 _09820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13927__A _14745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09982_ _09969_/X _09971_/X _09973_/X _09981_/X _09876_/A vssd1 vssd1 vccd1 vccd1
+ _09982_/X sky130_fd_sc_hd__a221o_1
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12831__A _12831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11710__A1 _18470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16449__S _16457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09416_ _18948_/Q _18947_/Q vssd1 vssd1 vccd1 vccd1 _14225_/C sky130_fd_sc_hd__or2_1
XFILLER_16_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13215__A1 _13627_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09347_ _18833_/Q vssd1 vssd1 vccd1 vccd1 _09347_/X sky130_fd_sc_hd__buf_4
XANTENNA__16184__S _16184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__B1 _13307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09587__A _11273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09278_ _09481_/A _09481_/B _09481_/C _09481_/D vssd1 vssd1 vccd1 vccd1 _09436_/D
+ sky130_fd_sc_hd__and4bb_1
XFILLER_154_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16912__S _16914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11121__S _11121_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11240_ _11225_/A _11235_/X _11237_/X _11239_/X vssd1 vssd1 vccd1 vccd1 _11240_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11171_ _11441_/S vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10122_ _11467_/S vssd1 vssd1 vccd1 vccd1 _10657_/S sky130_fd_sc_hd__buf_2
XFILLER_79_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17743__S _17749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11357__A _19385_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _10260_/A vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__buf_2
X_14930_ _14928_/X _14929_/X _14938_/S vssd1 vssd1 vccd1 vccd1 _14930_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input26_A io_dbus_rdata[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14861_ _14927_/A vssd1 vssd1 vccd1 vccd1 _14915_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__16359__S _16362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14668__A _15813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16600_ _19279_/Q _13832_/X _16602_/S vssd1 vssd1 vccd1 vccd1 _16601_/A sky130_fd_sc_hd__mux2_1
X_13812_ _13812_/A vssd1 vssd1 vccd1 vccd1 _18502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17580_ _17122_/X _19694_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17581_/A sky130_fd_sc_hd__mux2_1
X_14792_ _14792_/A _14792_/B vssd1 vssd1 vccd1 vccd1 _14795_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16531_ _16531_/A vssd1 vssd1 vccd1 vccd1 _19248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10955_ _11237_/A _10954_/X _10947_/A vssd1 vssd1 vccd1 vccd1 _10955_/X sky130_fd_sc_hd__a21o_1
X_13743_ _13739_/Y _13742_/X _16066_/S vssd1 vssd1 vccd1 vccd1 _13743_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11560__S0 _11566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19250_ _19939_/CLK _19250_/D vssd1 vssd1 vccd1 vccd1 _19250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16462_ _19218_/Q _13842_/X _16468_/S vssd1 vssd1 vccd1 vccd1 _16463_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10886_ _10886_/A _10886_/B vssd1 vssd1 vccd1 vccd1 _10886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13674_ _13681_/B _13673_/Y _13648_/X vssd1 vssd1 vccd1 vccd1 _13674_/Y sky130_fd_sc_hd__a21oi_2
X_18201_ _18201_/A vssd1 vssd1 vccd1 vccd1 _19941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15413_ _15413_/A vssd1 vssd1 vccd1 vccd1 _15413_/X sky130_fd_sc_hd__clkbuf_2
X_19181_ _19966_/CLK _19181_/D vssd1 vssd1 vccd1 vccd1 _19181_/Q sky130_fd_sc_hd__dfxtp_1
X_12625_ _12621_/X _12624_/Y _12814_/S vssd1 vssd1 vccd1 vccd1 _12625_/X sky130_fd_sc_hd__mux2_1
X_16393_ _17729_/A vssd1 vssd1 vccd1 vccd1 _16393_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16094__S _16100_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12916__A _18939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18132_ _18132_/A vssd1 vssd1 vccd1 vccd1 _19911_/D sky130_fd_sc_hd__clkbuf_1
X_12556_ _12556_/A vssd1 vssd1 vccd1 vccd1 _12556_/X sky130_fd_sc_hd__clkbuf_2
X_15344_ _12390_/Y _15279_/X _15343_/X _15275_/X vssd1 vssd1 vccd1 vccd1 _15344_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_11_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ _18846_/Q _09843_/A _09882_/A _11506_/X vssd1 vssd1 vccd1 vccd1 _12842_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_89_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17918__S _17926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18063_ _18843_/Q _13591_/X _18067_/S vssd1 vssd1 vccd1 vccd1 _18063_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16822__S _16830_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12487_ _12032_/X _14763_/C _12486_/Y vssd1 vssd1 vccd1 vccd1 _15397_/A sky130_fd_sc_hd__a21o_4
X_15275_ _15920_/A vssd1 vssd1 vccd1 vccd1 _15275_/X sky130_fd_sc_hd__buf_2
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17014_ _17014_/A vssd1 vssd1 vccd1 vccd1 _17014_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11438_ _11431_/X _11433_/X _11435_/X _11437_/X _09802_/A vssd1 vssd1 vccd1 vccd1
+ _11438_/X sky130_fd_sc_hd__a221o_4
X_14226_ _14226_/A _14226_/B _14226_/C vssd1 vssd1 vccd1 vccd1 _14227_/D sky130_fd_sc_hd__or3_1
XANTENNA_output94_A _12791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14157_ _14191_/A _14164_/C vssd1 vssd1 vccd1 vccd1 _14157_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11369_ _11199_/A _11368_/X _11335_/A vssd1 vssd1 vccd1 vccd1 _11369_/X sky130_fd_sc_hd__a21o_1
XFILLER_153_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13108_ _18842_/Q _13577_/B _13226_/A vssd1 vssd1 vccd1 vccd1 _13108_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14088_ _14088_/A _14088_/B _14088_/C vssd1 vssd1 vccd1 vccd1 _18605_/D sky130_fd_sc_hd__nor3_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18965_ _18992_/CLK _18965_/D vssd1 vssd1 vccd1 vccd1 _18965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13142__B1 _13359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17916_ _17916_/A vssd1 vssd1 vccd1 vccd1 _19829_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15962__A _15966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13039_ _13028_/X _13037_/X _13350_/S vssd1 vssd1 vccd1 vccd1 _13039_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18896_ _18928_/CLK _18896_/D vssd1 vssd1 vccd1 vccd1 _18896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17847_ _17847_/A vssd1 vssd1 vccd1 vccd1 _19798_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16269__S _16269_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17778_ _17691_/X _19768_/Q _17782_/S vssd1 vssd1 vccd1 vccd1 _17779_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10299__A2_N _09843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19517_ _19942_/CLK _19517_/D vssd1 vssd1 vccd1 vccd1 _19517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16729_ _16729_/A vssd1 vssd1 vccd1 vccd1 _19335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15901__S _15901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19448_ _19972_/CLK _19448_/D vssd1 vssd1 vccd1 vccd1 _19448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09201_ _18974_/Q _18975_/Q vssd1 vssd1 vccd1 vccd1 _09256_/A sky130_fd_sc_hd__or2b_1
XFILLER_50_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13748__A2 _13495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19379_ _19379_/CLK _19379_/D vssd1 vssd1 vccd1 vccd1 _19379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11730__A _11730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10431__A1 _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17828__S _17832_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16732__S _16736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16033__A _16044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09965_ _10129_/S vssd1 vssd1 vccd1 vccd1 _10180_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09896_ _19381_/Q _19716_/Q _09903_/A vssd1 vssd1 vccd1 vccd1 _09897_/B sky130_fd_sc_hd__mux2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10042__S0 _10275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09983__S0 _09967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18394__S _18396_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10345__S1 _10223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11542__S0 _11534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10740_ _18438_/Q _19467_/Q _19504_/Q _19078_/Q _10750_/S _10626_/A vssd1 vssd1 vccd1
+ vccd1 _10740_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10671_ _18439_/Q _19468_/Q _19505_/Q _19079_/Q _09652_/A _10656_/A vssd1 vssd1 vccd1
+ vccd1 _10671_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14936__A1 _12298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18127__A1 _13733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16208__A _16208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ _15947_/C _18912_/Q _12517_/S vssd1 vssd1 vccd1 vccd1 _14877_/A sky130_fd_sc_hd__mux2_4
XFILLER_159_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13390_ _18890_/Q _18891_/Q _13390_/C vssd1 vssd1 vccd1 vccd1 _13427_/C sky130_fd_sc_hd__and3_1
XFILLER_167_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12341_ _12341_/A _12416_/D vssd1 vssd1 vccd1 vccd1 _12341_/X sky130_fd_sc_hd__or2_1
XFILLER_166_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15060_ _15169_/A vssd1 vssd1 vccd1 vccd1 _15280_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12272_ _12272_/A _12272_/B vssd1 vssd1 vccd1 vccd1 _12273_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__15361__A1 _12413_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14011_ _18578_/Q _14013_/C _14010_/Y vssd1 vssd1 vccd1 vccd1 _18578_/D sky130_fd_sc_hd__o21a_1
X_11223_ _18837_/Q _09537_/A _11211_/X _11222_/Y vssd1 vssd1 vccd1 vccd1 _11223_/X
+ sky130_fd_sc_hd__a22o_2
XANTENNA__17039__A _17039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ _11154_/A vssd1 vssd1 vccd1 vccd1 _11155_/A sky130_fd_sc_hd__buf_2
XFILLER_161_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7_0_clock_A clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17473__S _17481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10105_ _15970_/C _12857_/B vssd1 vssd1 vccd1 vccd1 _10248_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18750_ _18762_/CLK _18750_/D vssd1 vssd1 vccd1 vccd1 _18750_/Q sky130_fd_sc_hd__dfxtp_1
X_15962_ _15966_/A _15966_/B _15962_/C vssd1 vssd1 vccd1 vccd1 _15962_/X sky130_fd_sc_hd__and3_1
X_11085_ _11388_/A vssd1 vssd1 vccd1 vccd1 _11086_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14872__A0 _15234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17701_ _17717_/A vssd1 vssd1 vccd1 vccd1 _17714_/S sky130_fd_sc_hd__buf_4
XANTENNA__18063__A0 _18843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__A1 _09884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ _10210_/A _10036_/B vssd1 vssd1 vccd1 vccd1 _10036_/Y sky130_fd_sc_hd__nand2_1
X_14913_ _15160_/B _12715_/A _14915_/S vssd1 vssd1 vccd1 vccd1 _14913_/X sky130_fd_sc_hd__mux2_1
X_18681_ _18687_/CLK _18681_/D vssd1 vssd1 vccd1 vccd1 _18681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15893_ _12260_/A _15842_/X _15879_/X input57/X vssd1 vssd1 vccd1 vccd1 _15894_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16089__S _16089_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17632_ _17198_/X _19718_/Q _17632_/S vssd1 vssd1 vccd1 vccd1 _17633_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11815__A _11815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14844_ _14973_/B _14846_/B vssd1 vssd1 vccd1 vccd1 _15384_/A sky130_fd_sc_hd__nor2_2
XFILLER_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17563_ _17619_/A vssd1 vssd1 vccd1 vccd1 _17632_/S sky130_fd_sc_hd__buf_6
X_14775_ _12866_/A _09279_/X _15747_/A _14778_/A _18825_/Q vssd1 vssd1 vccd1 vccd1
+ _14776_/B sky130_fd_sc_hd__a32o_1
XANTENNA__16817__S _16819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11987_ _12078_/C vssd1 vssd1 vccd1 vccd1 _15094_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10336__S1 _10153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19302_ _19637_/CLK _19302_/D vssd1 vssd1 vccd1 vccd1 _19302_/Q sky130_fd_sc_hd__dfxtp_1
X_16514_ _16514_/A vssd1 vssd1 vccd1 vccd1 _19240_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13726_ _13726_/A _19022_/Q vssd1 vssd1 vccd1 vccd1 _13726_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17494_ _17195_/X _19653_/Q _17496_/S vssd1 vssd1 vccd1 vccd1 _17495_/A sky130_fd_sc_hd__mux2_1
X_10938_ _10929_/A _10937_/X _09560_/A vssd1 vssd1 vccd1 vccd1 _10938_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19233_ _20018_/CLK _19233_/D vssd1 vssd1 vccd1 vccd1 _19233_/Q sky130_fd_sc_hd__dfxtp_1
X_16445_ _16445_/A vssd1 vssd1 vccd1 vccd1 _19210_/D sky130_fd_sc_hd__clkbuf_1
X_10869_ _15936_/B _12839_/B vssd1 vssd1 vccd1 vccd1 _11617_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18118__A1 _13710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13657_ _19013_/Q _13657_/B vssd1 vssd1 vccd1 vccd1 _13657_/X sky130_fd_sc_hd__or2_1
XANTENNA__12646__A _18542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19164_ _20016_/CLK _19164_/D vssd1 vssd1 vccd1 vccd1 _19164_/Q sky130_fd_sc_hd__dfxtp_1
X_12608_ _12601_/A _12553_/X _12604_/Y _12607_/Y vssd1 vssd1 vccd1 vccd1 _12608_/X
+ sky130_fd_sc_hd__o22a_2
X_16376_ _16376_/A vssd1 vssd1 vccd1 vccd1 _19183_/D sky130_fd_sc_hd__clkbuf_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _19004_/Q _13588_/B vssd1 vssd1 vccd1 vccd1 _13588_/X sky130_fd_sc_hd__or2_1
XFILLER_12_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18115_ _18115_/A vssd1 vssd1 vccd1 vccd1 _18128_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_158_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15327_ _12364_/Y _15279_/X _15326_/X _15275_/X vssd1 vssd1 vccd1 vccd1 _15327_/X
+ sky130_fd_sc_hd__a211o_1
X_19095_ _19856_/CLK _19095_/D vssd1 vssd1 vccd1 vccd1 _19095_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16552__S _16558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12539_ _12588_/A _12539_/B _12539_/C vssd1 vssd1 vccd1 vccd1 _12540_/A sky130_fd_sc_hd__or3_2
XANTENNA__14861__A _14927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18046_ _18838_/Q _13546_/X _18050_/S vssd1 vssd1 vccd1 vccd1 _18046_/X sky130_fd_sc_hd__mux2_1
X_15258_ _15428_/A vssd1 vssd1 vccd1 vccd1 _15258_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14209_ _18642_/Q _14212_/C vssd1 vssd1 vccd1 vccd1 _14210_/B sky130_fd_sc_hd__and2_1
XFILLER_99_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15189_ _15058_/X _15062_/X _15189_/S vssd1 vssd1 vccd1 vccd1 _15189_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19997_ _19997_/CLK _19997_/D vssd1 vssd1 vccd1 vccd1 _19997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16788__A _16834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17383__S _17387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09750_ _09750_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09750_/X sky130_fd_sc_hd__or2_1
X_18948_ _18958_/CLK _18948_/D vssd1 vssd1 vccd1 vccd1 _18948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18054__A0 _18840_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09681_ _09681_/A vssd1 vssd1 vccd1 vccd1 _09682_/A sky130_fd_sc_hd__clkbuf_4
X_18879_ _19010_/CLK _18879_/D vssd1 vssd1 vccd1 vccd1 _18879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14615__A0 _12452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11429__B1 _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14091__A1 _18606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13940__A _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15631__S _15901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12556__A _12556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13151__S _13203_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11460__A _11462_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13051__C1 _11791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16462__S _16468_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14771__A _14771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18243__A _18265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10168__B1 _10001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10804__A _10858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13106__B1 _12890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17293__S _17293_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ _09765_/A _09947_/X _09837_/A vssd1 vssd1 vccd1 vccd1 _09948_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__14710__S _14716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09879_ _09909_/A _09697_/X _09698_/X _09699_/Y vssd1 vssd1 vccd1 vccd1 _09880_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _12055_/A _12055_/B _12055_/C _09471_/X vssd1 vssd1 vccd1 vccd1 _12196_/A
+ sky130_fd_sc_hd__or4b_2
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13409__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12890_ _12890_/A vssd1 vssd1 vccd1 vccd1 _12890_/X sky130_fd_sc_hd__buf_2
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10891__A1 _09546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11841_/A vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _11772_/A _11772_/B vssd1 vssd1 vccd1 vccd1 _11773_/A sky130_fd_sc_hd__and2_2
X_14560_ _14560_/A _18995_/Q vssd1 vssd1 vccd1 vccd1 _14560_/Y sky130_fd_sc_hd__nand2_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _10723_/A _10723_/B vssd1 vssd1 vccd1 vccd1 _10723_/Y sky130_fd_sc_hd__nor2_1
X_13511_ _13511_/A _13511_/B _13511_/C vssd1 vssd1 vccd1 vccd1 _13511_/X sky130_fd_sc_hd__and3_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14491_ _14493_/B _14493_/C _14465_/X vssd1 vssd1 vccd1 vccd1 _14491_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13061__S _13215_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16230_ _12939_/X _19129_/Q _16236_/S vssd1 vssd1 vccd1 vccd1 _16231_/A sky130_fd_sc_hd__mux2_1
X_10654_ _10654_/A vssd1 vssd1 vccd1 vccd1 _10656_/A sky130_fd_sc_hd__buf_2
XFILLER_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13442_ _17084_/A vssd1 vssd1 vccd1 vccd1 _17726_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17468__S _17470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16161_ _16161_/A vssd1 vssd1 vccd1 vccd1 _19099_/D sky130_fd_sc_hd__clkbuf_1
X_13373_ _19906_/Q _13373_/B vssd1 vssd1 vccd1 vccd1 _13373_/X sky130_fd_sc_hd__and2_1
XANTENNA__16372__S _16378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10585_ _15952_/C _12848_/B vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__or2_1
XFILLER_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15112_ _15110_/X _15111_/X _15202_/S vssd1 vssd1 vccd1 vccd1 _15112_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09775__A _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12324_ _12459_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__nand2_1
X_16092_ _13023_/X _19069_/Q _16100_/S vssd1 vssd1 vccd1 vccd1 _16093_/A sky130_fd_sc_hd__mux2_1
X_12255_ _18766_/Q _18765_/Q _12255_/C vssd1 vssd1 vccd1 vccd1 _12309_/C sky130_fd_sc_hd__and3_1
X_19920_ _19981_/CLK _19920_/D vssd1 vssd1 vccd1 vccd1 _19920_/Q sky130_fd_sc_hd__dfxtp_1
X_15043_ _15038_/X _15041_/X _15199_/S vssd1 vssd1 vccd1 vccd1 _15043_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13896__A1 _12554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_3_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11206_ _11206_/A vssd1 vssd1 vccd1 vccd1 _11287_/A sky130_fd_sc_hd__clkbuf_2
X_19851_ _19949_/CLK _19851_/D vssd1 vssd1 vccd1 vccd1 _19851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_156_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12186_ _12215_/D _12186_/B vssd1 vssd1 vccd1 vccd1 _12186_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_96_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold4_A hold4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18802_ _19912_/CLK _18802_/D vssd1 vssd1 vccd1 vccd1 _18802_/Q sky130_fd_sc_hd__dfxtp_1
X_11137_ _11137_/A _11137_/B vssd1 vssd1 vccd1 vccd1 _11137_/X sky130_fd_sc_hd__or2_1
X_19782_ _19842_/CLK _19782_/D vssd1 vssd1 vccd1 vccd1 _19782_/Q sky130_fd_sc_hd__dfxtp_1
X_16994_ _17075_/A vssd1 vssd1 vccd1 vccd1 _17094_/S sky130_fd_sc_hd__buf_6
XFILLER_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10006__S0 _10275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18733_ _18734_/CLK _18733_/D vssd1 vssd1 vccd1 vccd1 _18733_/Q sky130_fd_sc_hd__dfxtp_1
X_11068_ _11068_/A vssd1 vssd1 vccd1 vccd1 _11335_/A sky130_fd_sc_hd__clkbuf_2
X_15945_ _15945_/A vssd1 vssd1 vccd1 vccd1 _15966_/A sky130_fd_sc_hd__buf_2
XFILLER_95_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17931__S _17937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _10859_/S vssd1 vssd1 vccd1 vccd1 _10749_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18664_ _18734_/CLK _18664_/D vssd1 vssd1 vccd1 vccd1 _18664_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10331__B1 _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15876_ _09261_/B _15875_/X _15820_/X input51/X vssd1 vssd1 vccd1 vccd1 _15877_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17615_ _17173_/X _19710_/Q _17617_/S vssd1 vssd1 vccd1 vccd1 _17616_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14827_ _14869_/A vssd1 vssd1 vccd1 vccd1 _14955_/S sky130_fd_sc_hd__clkbuf_2
X_18595_ _19683_/CLK _18595_/D vssd1 vssd1 vccd1 vccd1 _18595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12084__A0 hold4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17546_ _19679_/Q vssd1 vssd1 vccd1 vccd1 _17547_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14758_ _14758_/A _14758_/B vssd1 vssd1 vccd1 vccd1 _14814_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13709_ _13709_/A _19020_/Q vssd1 vssd1 vccd1 vccd1 _13709_/Y sky130_fd_sc_hd__nand2_1
X_17477_ _17170_/X _19645_/Q _17481_/S vssd1 vssd1 vccd1 vccd1 _17478_/A sky130_fd_sc_hd__mux2_1
X_14689_ _14689_/A vssd1 vssd1 vccd1 vccd1 _18796_/D sky130_fd_sc_hd__clkbuf_1
X_19216_ _20034_/CLK _19216_/D vssd1 vssd1 vccd1 vccd1 _19216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16428_ _16428_/A vssd1 vssd1 vccd1 vccd1 _19202_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12095__B _12583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19147_ _19996_/CLK _19147_/D vssd1 vssd1 vccd1 vccd1 _19147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16359_ _16358_/X _19178_/Q _16362_/S vssd1 vssd1 vccd1 vccd1 _16360_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19078_ _19990_/CLK _19078_/D vssd1 vssd1 vccd1 vccd1 _19078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13336__B1 _09405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18029_ _09444_/B _12163_/B _18028_/X _11915_/B vssd1 vssd1 vccd1 vccd1 _18115_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__10624__A _10624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09802_ _09802_/A vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09960__C1 _09807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13639__A1 _13638_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18027__A0 _09347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09733_ _09950_/S vssd1 vssd1 vccd1 vccd1 _09733_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12311__A1 _12188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17841__S _17843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09664_ _09664_/A vssd1 vssd1 vccd1 vccd1 _10822_/A sky130_fd_sc_hd__buf_2
XANTENNA__10322__B1 _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09595_ _09595_/A vssd1 vssd1 vccd1 vccd1 _10251_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16457__S _16457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14766__A _14766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13092__D input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12075__B1 _12074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13811__A1 _13810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10389__B1 _10001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09595__A _09595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10370_ _20030_/Q _19868_/Q _19277_/Q _19047_/Q _10251_/S _10054_/A vssd1 vssd1 vccd1
+ vccd1 _10370_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12733__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15867__A2 _15856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12040_ _11292_/X _18900_/Q _12179_/S vssd1 vssd1 vccd1 vccd1 _14895_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17317__A _17339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10561__B1 _09539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13991_ _13991_/A _13991_/B _13992_/B vssd1 vssd1 vccd1 vccd1 _18571_/D sky130_fd_sc_hd__nor3_1
XFILLER_74_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _15769_/A vssd1 vssd1 vccd1 vccd1 _15730_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _18552_/Q vssd1 vssd1 vccd1 vccd1 _13936_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_86_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _15661_/A vssd1 vssd1 vccd1 vccd1 _18908_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12873_ _13233_/A vssd1 vssd1 vccd1 vccd1 _13223_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _17411_/A vssd1 vssd1 vccd1 vccd1 _17409_/S sky130_fd_sc_hd__clkbuf_8
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17052__A _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14612_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14613_/A sky130_fd_sc_hd__and2_1
X_18380_ _18380_/A vssd1 vssd1 vccd1 vccd1 _20020_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _11824_/A vssd1 vssd1 vccd1 vccd1 _12887_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15592_ _18878_/Q _18910_/Q _15600_/S vssd1 vssd1 vccd1 vccd1 _15593_/A sky130_fd_sc_hd__mux2_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17167_/X _19580_/Q _17337_/S vssd1 vssd1 vccd1 vccd1 _17332_/A sky130_fd_sc_hd__mux2_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14543_ _18753_/Q _11865_/X _14542_/X _14540_/X vssd1 vssd1 vccd1 vccd1 _18753_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11870_/A vssd1 vssd1 vccd1 vccd1 _11755_/X sky130_fd_sc_hd__buf_2
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_82_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _17262_/A vssd1 vssd1 vccd1 vccd1 _19549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10706_ _10723_/A _10706_/B vssd1 vssd1 vccd1 vccd1 _10706_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14474_ _14476_/B _14476_/C _14465_/X vssd1 vssd1 vccd1 vccd1 _14474_/Y sky130_fd_sc_hd__a21oi_1
X_11686_ _11686_/A vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19001_ _19001_/CLK _19001_/D vssd1 vssd1 vccd1 vccd1 _19001_/Q sky130_fd_sc_hd__dfxtp_1
X_16213_ _13423_/X _19123_/Q _16217_/S vssd1 vssd1 vccd1 vccd1 _16214_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13566__B1 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13425_ _13425_/A vssd1 vssd1 vccd1 vccd1 _18451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10637_ _19240_/Q _19735_/Q _10637_/S vssd1 vssd1 vccd1 vccd1 _10637_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17193_ _17192_/X _19519_/Q _17193_/S vssd1 vssd1 vccd1 vccd1 _17194_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13030__A2 _12943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15938__C _15938_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10475__S0 _10208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16144_ _13463_/X _19093_/Q _16144_/S vssd1 vssd1 vccd1 vccd1 _16145_/A sky130_fd_sc_hd__mux2_1
X_13356_ _13356_/A vssd1 vssd1 vccd1 vccd1 _18447_/D sky130_fd_sc_hd__clkbuf_1
X_10568_ _20026_/Q _19864_/Q _19273_/Q _19043_/Q _10529_/S _10011_/A vssd1 vssd1 vccd1
+ vccd1 _10568_/X sky130_fd_sc_hd__mux4_1
XFILLER_143_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11552__A1_N _18864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17926__S _17926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12307_ _18465_/Q _12372_/B vssd1 vssd1 vccd1 vccd1 _12307_/X sky130_fd_sc_hd__or2_1
X_16075_ _16075_/A _16075_/B vssd1 vssd1 vccd1 vccd1 _16075_/X sky130_fd_sc_hd__or2_1
X_10499_ _19146_/Q _19407_/Q _19306_/Q _19641_/Q _10543_/S _10497_/A vssd1 vssd1 vccd1
+ vccd1 _10500_/B sky130_fd_sc_hd__mux4_1
XANTENNA__16830__S _16830_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13287_ _13664_/A _13288_/B vssd1 vssd1 vccd1 vccd1 _13289_/B sky130_fd_sc_hd__nor2_1
X_15026_ _15169_/A vssd1 vssd1 vccd1 vccd1 _15190_/S sky130_fd_sc_hd__clkbuf_2
X_19903_ _19910_/CLK _19903_/D vssd1 vssd1 vccd1 vccd1 _19903_/Q sky130_fd_sc_hd__dfxtp_1
X_12238_ _15254_/A _12238_/B vssd1 vssd1 vccd1 vccd1 _12242_/A sky130_fd_sc_hd__xnor2_1
XFILLER_123_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13755__A _17098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19834_ _19972_/CLK _19834_/D vssd1 vssd1 vccd1 vccd1 _19834_/Q sky130_fd_sc_hd__dfxtp_1
X_12169_ _13518_/A vssd1 vssd1 vccd1 vccd1 _12347_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19765_ _20023_/CLK _19765_/D vssd1 vssd1 vccd1 vccd1 _19765_/Q sky130_fd_sc_hd__dfxtp_1
X_16977_ _16977_/A vssd1 vssd1 vccd1 vccd1 _16986_/S sky130_fd_sc_hd__buf_4
XFILLER_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput5 io_dbus_rdata[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15970__A _15978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18716_ _18744_/CLK _18716_/D vssd1 vssd1 vccd1 vccd1 _18716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15928_ _15928_/A vssd1 vssd1 vccd1 vccd1 _15928_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19696_ _20018_/CLK _19696_/D vssd1 vssd1 vccd1 vccd1 _19696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18647_ _18688_/CLK _18647_/D vssd1 vssd1 vccd1 vccd1 _18647_/Q sky130_fd_sc_hd__dfxtp_1
X_15859_ _15859_/A vssd1 vssd1 vccd1 vccd1 _18980_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14586__A _14595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09380_ _11705_/A _14227_/B _11700_/B vssd1 vssd1 vccd1 vccd1 _13510_/A sky130_fd_sc_hd__o21ai_1
XFILLER_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18578_ _18819_/CLK _18578_/D vssd1 vssd1 vccd1 vccd1 _18578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17529_ _17529_/A vssd1 vssd1 vccd1 vccd1 _19670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10619__A _11186_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15806__A1_N _15805_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13557__A0 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12834__A _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10769__S1 _10663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17571__S _17573_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ _09957_/A vssd1 vssd1 vccd1 vccd1 _09750_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09647_ _09647_/A vssd1 vssd1 vccd1 vccd1 _09660_/A sky130_fd_sc_hd__buf_4
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09578_ _10508_/A vssd1 vssd1 vccd1 vccd1 _10458_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_104_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ _09868_/A _11539_/X _09690_/X vssd1 vssd1 vccd1 vccd1 _11540_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11271__A1 _10983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15537__A1 _18862_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13548__A0 _13546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11471_ _19333_/Q _19604_/Q _19828_/Q _19572_/Q _10821_/S _10597_/A vssd1 vssd1 vccd1
+ vccd1 _11471_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ _19675_/Q _19441_/Q _18506_/Q _19771_/Q _10388_/S _10153_/A vssd1 vssd1 vccd1
+ vccd1 _10422_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13210_ _18469_/Q _11740_/X _12944_/A _18693_/Q _13209_/X vssd1 vssd1 vccd1 vccd1
+ _13210_/X sky130_fd_sc_hd__a221o_1
XANTENNA__09529__S _15127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10457__S0 _10180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ _18636_/Q _14190_/B vssd1 vssd1 vccd1 vccd1 _14197_/C sky130_fd_sc_hd__and2_2
XFILLER_152_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12771__A1 _18483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10353_ _19676_/Q _19442_/Q _18507_/Q _19772_/Q _10356_/S _09636_/A vssd1 vssd1 vccd1
+ vccd1 _10353_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13141_ _18876_/Q vssd1 vssd1 vccd1 vccd1 _13603_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16650__S _16652_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13072_ _18686_/Q vssd1 vssd1 vccd1 vccd1 _14371_/B sky130_fd_sc_hd__clkbuf_2
X_10284_ _19343_/Q _19614_/Q _19838_/Q _19582_/Q _10279_/X _10283_/X vssd1 vssd1 vccd1
+ vccd1 _10285_/B sky130_fd_sc_hd__mux4_1
XANTENNA_input56_A io_ibus_inst[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16900_ _16900_/A vssd1 vssd1 vccd1 vccd1 _19411_/D sky130_fd_sc_hd__clkbuf_1
X_12023_ _12020_/X _12016_/X _12168_/S _13650_/A vssd1 vssd1 vccd1 vccd1 _12023_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_29_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17880_ _19814_/Q _17093_/X _17880_/S vssd1 vssd1 vccd1 vccd1 _17881_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_opt_2_0_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16831_ _16831_/A vssd1 vssd1 vccd1 vccd1 _19381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17481__S _17481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19550_ _19936_/CLK _19550_/D vssd1 vssd1 vccd1 vccd1 _19550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16762_ _19351_/Q _13857_/X _16762_/S vssd1 vssd1 vccd1 vccd1 _16763_/A sky130_fd_sc_hd__mux2_1
X_13974_ _13991_/A _13974_/B _13976_/B vssd1 vssd1 vccd1 vccd1 _18565_/D sky130_fd_sc_hd__nor3_1
XFILLER_47_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18501_ _19767_/CLK _18501_/D vssd1 vssd1 vccd1 vccd1 _18501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15713_ _17208_/A vssd1 vssd1 vccd1 vccd1 _15713_/X sky130_fd_sc_hd__clkbuf_2
X_19481_ _19587_/CLK _19481_/D vssd1 vssd1 vccd1 vccd1 _19481_/Q sky130_fd_sc_hd__dfxtp_1
X_12925_ _12925_/A vssd1 vssd1 vccd1 vccd1 _18424_/D sky130_fd_sc_hd__clkbuf_1
X_16693_ _16749_/A vssd1 vssd1 vccd1 vccd1 _16762_/S sky130_fd_sc_hd__buf_6
XFILLER_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18432_ _19567_/CLK _18432_/D vssd1 vssd1 vccd1 vccd1 _18432_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15644_ _18901_/Q _18522_/Q _15644_/S vssd1 vssd1 vccd1 vccd1 _15645_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16973__A0 _16374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15776__A1 _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ _12857_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12856_/Y sky130_fd_sc_hd__nor2_4
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12638__B _14907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _14544_/B _11774_/A _11803_/X _15738_/B vssd1 vssd1 vccd1 vccd1 _18746_/D
+ sky130_fd_sc_hd__a22o_1
X_18363_ _17649_/X _20013_/Q _18363_/S vssd1 vssd1 vccd1 vccd1 _18364_/A sky130_fd_sc_hd__mux2_1
X_15575_ _15575_/A vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__clkbuf_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _12742_/A _12742_/B _12763_/B _12741_/A vssd1 vssd1 vccd1 vccd1 _12788_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_109_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17314_ _17314_/A vssd1 vssd1 vccd1 vccd1 _19572_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _18743_/Q _14526_/B _14526_/C vssd1 vssd1 vccd1 vccd1 _14528_/B sky130_fd_sc_hd__and3_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _12946_/A vssd1 vssd1 vccd1 vccd1 _13451_/B sky130_fd_sc_hd__buf_2
X_18294_ _17652_/X _19982_/Q _18302_/S vssd1 vssd1 vccd1 vccd1 _18295_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15949__B _15949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17245_ _17267_/A vssd1 vssd1 vccd1 vccd1 _17254_/S sky130_fd_sc_hd__buf_2
XFILLER_30_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10873__S _10921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14457_ _14459_/B _14459_/C _14456_/Y vssd1 vssd1 vccd1 vccd1 _18718_/D sky130_fd_sc_hd__o21a_1
X_11669_ _12153_/B _12153_/C vssd1 vssd1 vccd1 vccd1 _19880_/D sky130_fd_sc_hd__nand2_1
X_13408_ _13408_/A vssd1 vssd1 vccd1 vccd1 _18450_/D sky130_fd_sc_hd__clkbuf_1
X_17176_ _17713_/A vssd1 vssd1 vccd1 vccd1 _17176_/X sky130_fd_sc_hd__clkbuf_2
X_14388_ _18692_/Q _18691_/Q _14391_/D _14094_/A vssd1 vssd1 vccd1 vccd1 _14388_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_143_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16127_ _13323_/X _19085_/Q _16133_/S vssd1 vssd1 vccd1 vccd1 _16128_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13339_ _13188_/X _13683_/B _13338_/X _13289_/A vssd1 vssd1 vccd1 vccd1 _13339_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09963__A _15976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16058_ _16058_/A vssd1 vssd1 vccd1 vccd1 _19057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15009_ _14944_/X _14947_/X _15014_/S vssd1 vssd1 vccd1 vccd1 _15009_/X sky130_fd_sc_hd__mux2_1
X_19817_ _19947_/CLK _19817_/D vssd1 vssd1 vccd1 vccd1 _19817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15904__S _15946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19748_ _19810_/CLK _19748_/D vssd1 vssd1 vccd1 vccd1 _19748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09501_ _09502_/A _09501_/B vssd1 vssd1 vccd1 vccd1 _14804_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19679_ _20033_/CLK _19679_/D vssd1 vssd1 vccd1 vccd1 _19679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12829__A _12829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13424__S _13464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10923__S1 _10663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09432_ _15914_/S vssd1 vssd1 vccd1 vccd1 _15457_/A sky130_fd_sc_hd__buf_4
XANTENNA__15767__A1 _14749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09363_ _12064_/A _09361_/X _09362_/X _18746_/Q vssd1 vssd1 vccd1 vccd1 _12062_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_162_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09294_ _18936_/Q _18976_/Q vssd1 vssd1 vccd1 vccd1 _09294_/X sky130_fd_sc_hd__and2b_1
XFILLER_36_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14763__B _15553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_3_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__S0 _10141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15875__A _15875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13950__B1 _13949_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16470__S _16472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09873__A _09873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput150 _12485_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[17] sky130_fd_sc_hd__buf_2
XFILLER_133_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput161 _12728_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[27] sky130_fd_sc_hd__buf_2
XANTENNA__12505__A1 _18472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput172 _12235_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[8] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_30_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10611__S0 _10655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15455__B1 _15453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ _11131_/A vssd1 vssd1 vccd1 vccd1 _11252_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12710_ _12709_/Y _18924_/Q _12782_/S vssd1 vssd1 vccd1 vccd1 _12713_/B sky130_fd_sc_hd__mux2_4
XFILLER_55_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_3_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _20012_/CLK sky130_fd_sc_hd__clkbuf_16
X_13690_ _13690_/A vssd1 vssd1 vccd1 vccd1 _13752_/S sky130_fd_sc_hd__buf_2
XFILLER_70_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12641_ _12641_/A vssd1 vssd1 vccd1 vccd1 _15463_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11244__A1 _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15360_ _15920_/A vssd1 vssd1 vccd1 vccd1 _15360_/X sky130_fd_sc_hd__clkbuf_2
X_12572_ _12572_/A _12572_/B vssd1 vssd1 vccd1 vccd1 _12574_/A sky130_fd_sc_hd__and2_2
XFILLER_11_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14311_ _14316_/B _14317_/D _14310_/Y vssd1 vssd1 vccd1 vccd1 _18669_/D sky130_fd_sc_hd__o21a_1
X_11523_ _11586_/A _11629_/A _11586_/C _10352_/A _11522_/Y vssd1 vssd1 vccd1 vccd1
+ _11634_/B sky130_fd_sc_hd__a311o_2
XFILLER_156_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15291_ _15291_/A _15291_/B vssd1 vssd1 vccd1 vccd1 _15291_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17030_ _17030_/A vssd1 vssd1 vccd1 vccd1 _17030_/X sky130_fd_sc_hd__clkbuf_2
X_14242_ _18649_/Q _18648_/Q _14242_/C _14242_/D vssd1 vssd1 vccd1 vccd1 _14256_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_156_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11454_ _11223_/X _12827_/B _11292_/X _12826_/B vssd1 vssd1 vccd1 vccd1 _11454_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10405_ _19340_/Q _19611_/Q _19835_/Q _19579_/Q _09995_/A _09610_/A vssd1 vssd1 vccd1
+ vccd1 _10405_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15785__A input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11385_ _18834_/Q vssd1 vssd1 vccd1 vccd1 _12934_/A sky130_fd_sc_hd__inv_2
X_14173_ _14189_/A _14173_/B _14174_/B vssd1 vssd1 vccd1 vccd1 _18629_/D sky130_fd_sc_hd__nor3_1
XFILLER_124_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ _18800_/Q _13071_/X _12879_/A _12283_/A _13123_/X vssd1 vssd1 vccd1 vccd1
+ _13124_/X sky130_fd_sc_hd__a221o_2
X_10336_ _19150_/Q _19411_/Q _19310_/Q _19645_/Q _10152_/X _10153_/X vssd1 vssd1 vccd1
+ vccd1 _10337_/B sky130_fd_sc_hd__mux4_1
XFILLER_139_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18981_ _19526_/CLK _18981_/D vssd1 vssd1 vccd1 vccd1 _18981_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_output162_A _12752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17932_ _17932_/A vssd1 vssd1 vccd1 vccd1 _19836_/D sky130_fd_sc_hd__clkbuf_1
X_10267_ _18447_/Q _19476_/Q _19513_/Q _19087_/Q _10059_/S _10261_/X vssd1 vssd1 vccd1
+ vccd1 _10267_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _18621_/Q _11794_/X _13053_/X _13054_/X vssd1 vssd1 vccd1 vccd1 _13055_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12006_ _18520_/Q _15633_/D vssd1 vssd1 vccd1 vccd1 _12007_/B sky130_fd_sc_hd__nor2_1
XFILLER_94_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17863_ _19806_/Q _17068_/X _17865_/S vssd1 vssd1 vccd1 vccd1 _17864_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10602__S0 _10655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10198_ _10369_/A _10197_/X _10107_/X vssd1 vssd1 vccd1 vccd1 _10198_/X sky130_fd_sc_hd__o21a_1
XFILLER_120_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19602_ _19829_/CLK _19602_/D vssd1 vssd1 vccd1 vccd1 _19602_/Q sky130_fd_sc_hd__dfxtp_1
X_16814_ _16814_/A vssd1 vssd1 vccd1 vccd1 _19373_/D sky130_fd_sc_hd__clkbuf_1
X_17794_ _17794_/A vssd1 vssd1 vccd1 vccd1 _19775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16745_ _19343_/Q _13832_/X _16747_/S vssd1 vssd1 vccd1 vccd1 _16746_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19533_ _20015_/CLK _19533_/D vssd1 vssd1 vccd1 vccd1 _19533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13957_ _13991_/A _13957_/B _13957_/C vssd1 vssd1 vccd1 vccd1 _18559_/D sky130_fd_sc_hd__nor3_1
XFILLER_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11553__A _11553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19464_ _19637_/CLK _19464_/D vssd1 vssd1 vccd1 vccd1 _19464_/Q sky130_fd_sc_hd__dfxtp_1
X_12908_ _16992_/A vssd1 vssd1 vccd1 vccd1 _17634_/A sky130_fd_sc_hd__clkbuf_2
X_16676_ _16676_/A vssd1 vssd1 vccd1 vccd1 _16685_/S sky130_fd_sc_hd__buf_4
XANTENNA__15749__A1 _15847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13888_ _13883_/X _12401_/Y _12402_/X _13946_/A vssd1 vssd1 vccd1 vccd1 _18532_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18415_ _18415_/A vssd1 vssd1 vccd1 vccd1 _20036_/D sky130_fd_sc_hd__clkbuf_1
X_15627_ _13737_/A _18926_/Q _15901_/S vssd1 vssd1 vccd1 vccd1 _15628_/A sky130_fd_sc_hd__mux2_1
X_12839_ _12833_/A _12839_/B vssd1 vssd1 vccd1 vccd1 _12840_/A sky130_fd_sc_hd__and2b_2
X_19395_ _19758_/CLK _19395_/D vssd1 vssd1 vccd1 vccd1 _19395_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18346_ _17729_/X _20006_/Q _18346_/S vssd1 vssd1 vccd1 vccd1 _18347_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ _14965_/A _15205_/X _15557_/X vssd1 vssd1 vccd1 vccd1 _15558_/X sky130_fd_sc_hd__a21o_1
XFILLER_148_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14509_ _14510_/B _14510_/C _14508_/Y vssd1 vssd1 vccd1 vccd1 _18736_/D sky130_fd_sc_hd__o21a_1
XFILLER_159_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18277_ _18277_/A vssd1 vssd1 vccd1 vccd1 _19975_/D sky130_fd_sc_hd__clkbuf_1
X_15489_ _15489_/A _15489_/B _15489_/C vssd1 vssd1 vccd1 vccd1 _15489_/X sky130_fd_sc_hd__and3_1
XANTENNA__12384__A _12385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14185__B1 _14160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17228_ _17122_/X _19534_/Q _17232_/S vssd1 vssd1 vccd1 vccd1 _17229_/A sky130_fd_sc_hd__mux2_1
Xinput30 io_dbus_rdata[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_6
XFILLER_174_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput41 io_ibus_inst[16] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_6
Xinput52 io_ibus_inst[26] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_6
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput63 io_ibus_inst[7] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_6
X_17159_ _17159_/A vssd1 vssd1 vccd1 vccd1 _19508_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11094__S0 _11158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09981_ _10270_/A _09979_/X _09980_/X vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10351__B _12854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11710__A2 _12943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11463__A _15936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09415_ _09381_/Y _11695_/A _09410_/X _09414_/X vssd1 vssd1 vccd1 vccd1 _09415_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_41_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10079__A _18857_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _18834_/Q vssd1 vssd1 vccd1 vccd1 _09425_/B sky130_fd_sc_hd__buf_4
XFILLER_166_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12974__A1 _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09277_ _09248_/X _09310_/C _09276_/X vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11170_ _15925_/C _12831_/B _11609_/A vssd1 vssd1 vccd1 vccd1 _11606_/A sky130_fd_sc_hd__o21ai_1
XFILLER_161_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_7_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ _11468_/S vssd1 vssd1 vccd1 vccd1 _11467_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_121_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15140__A2 _15138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__A _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ _10398_/A vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14860_ _14860_/A vssd1 vssd1 vccd1 vccd1 _15424_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13811_ _18502_/Q _13810_/X _13820_/S vssd1 vssd1 vccd1 vccd1 _13812_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input19_A io_dbus_rdata[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ _14791_/A _15740_/B vssd1 vssd1 vccd1 vccd1 _14791_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16530_ _19248_/Q _13835_/X _16530_/S vssd1 vssd1 vccd1 vccd1 _16531_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_151_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _18687_/CLK sky130_fd_sc_hd__clkbuf_16
X_13742_ _13531_/A _19024_/Q _09341_/X _13741_/X vssd1 vssd1 vccd1 vccd1 _13742_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_56_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10899__S0 _10892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ _19233_/Q _19728_/Q _10954_/S vssd1 vssd1 vccd1 vccd1 _10954_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11560__S1 _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16461_ _16461_/A vssd1 vssd1 vccd1 vccd1 _19217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16375__S _16378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13673_ _13664_/A _13672_/C _13306_/X vssd1 vssd1 vccd1 vccd1 _13673_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10885_ _19202_/Q _19793_/Q _19955_/Q _19170_/Q _10704_/A _10048_/A vssd1 vssd1 vccd1
+ vccd1 _10886_/B sky130_fd_sc_hd__mux4_1
X_18200_ _17726_/X _19941_/Q _18202_/S vssd1 vssd1 vccd1 vccd1 _18201_/A sky130_fd_sc_hd__mux2_1
X_15412_ _15438_/A _15412_/B _15412_/C vssd1 vssd1 vccd1 vccd1 _15412_/X sky130_fd_sc_hd__and3_1
X_19180_ _19965_/CLK _19180_/D vssd1 vssd1 vccd1 vccd1 _19180_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09778__A _10162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12624_ _12624_/A _12647_/B vssd1 vssd1 vccd1 vccd1 _12624_/Y sky130_fd_sc_hd__nor2_1
X_16392_ _16392_/A vssd1 vssd1 vccd1 vccd1 _19188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_166_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19880_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18131_ _18130_/X _19911_/Q _18134_/S vssd1 vssd1 vccd1 vccd1 _18132_/A sky130_fd_sc_hd__mux2_1
X_15343_ _15329_/X _15331_/X _15341_/X _15342_/X vssd1 vssd1 vccd1 vccd1 _15343_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12555_ _12551_/A _12554_/Y _12697_/S vssd1 vssd1 vccd1 vccd1 _12555_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11506_ _11491_/X _11496_/X _09820_/A _11505_/X vssd1 vssd1 vccd1 vccd1 _11506_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_18062_ _18062_/A vssd1 vssd1 vccd1 vccd1 _19890_/D sky130_fd_sc_hd__clkbuf_1
X_15274_ _15243_/X _15263_/X _15273_/X _15258_/X vssd1 vssd1 vccd1 vccd1 _15274_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ _12537_/A _12849_/B _12318_/B vssd1 vssd1 vccd1 vccd1 _12486_/Y sky130_fd_sc_hd__o21ai_1
X_17013_ _17013_/A vssd1 vssd1 vccd1 vccd1 _19458_/D sky130_fd_sc_hd__clkbuf_1
X_14225_ _18943_/Q _18938_/Q _14225_/C _14225_/D vssd1 vssd1 vccd1 vccd1 _14226_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11437_ _11111_/A _11436_/X _09788_/A vssd1 vssd1 vccd1 vccd1 _11437_/X sky130_fd_sc_hd__o21a_1
XANTENNA__16404__A _16472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output87_A _12645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10823__S0 _10872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13747__B _19025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14156_ _18624_/Q _18623_/Q _18622_/Q _14156_/D vssd1 vssd1 vccd1 vccd1 _14164_/C
+ sky130_fd_sc_hd__and4_1
X_11368_ _19225_/Q _19720_/Q _11410_/S vssd1 vssd1 vccd1 vccd1 _11368_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _18559_/Q _13070_/A _13104_/X _13105_/X _13106_/X vssd1 vssd1 vccd1 vccd1
+ _13577_/B sky130_fd_sc_hd__a2111o_4
X_10319_ _10319_/A vssd1 vssd1 vccd1 vccd1 _10319_/X sky130_fd_sc_hd__buf_4
XFILLER_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14086_/B _14086_/C _18605_/Q vssd1 vssd1 vccd1 vccd1 _14088_/C sky130_fd_sc_hd__a21oi_1
X_18964_ _18967_/CLK _18964_/D vssd1 vssd1 vccd1 vccd1 _18964_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _11164_/A _11294_/X _11296_/Y _11298_/Y vssd1 vssd1 vccd1 vccd1 _11299_/X
+ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_104_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19839_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17915_ _19829_/Q _17039_/X _17915_/S vssd1 vssd1 vccd1 vccd1 _17916_/A sky130_fd_sc_hd__mux2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13175_/A vssd1 vssd1 vccd1 vccd1 _13350_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_85_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15962__B _15966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18895_ _18928_/CLK _18895_/D vssd1 vssd1 vccd1 vccd1 _18895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17846_ _19798_/Q _17042_/X _17854_/S vssd1 vssd1 vccd1 vccd1 _17847_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17777_ _17777_/A vssd1 vssd1 vccd1 vccd1 _19767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14989_ _15444_/A vssd1 vssd1 vccd1 vccd1 _15438_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14642__A1 _11898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19747_/CLK sky130_fd_sc_hd__clkbuf_16
X_19516_ _19942_/CLK _19516_/D vssd1 vssd1 vccd1 vccd1 _19516_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11000__S0 _11048_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16728_ _19335_/Q _13806_/X _16736_/S vssd1 vssd1 vccd1 vccd1 _16729_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16659_ _16355_/X _19305_/Q _16663_/S vssd1 vssd1 vccd1 vccd1 _16660_/A sky130_fd_sc_hd__mux2_1
X_19447_ _19940_/CLK _19447_/D vssd1 vssd1 vccd1 vccd1 _19447_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16285__S _16291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09200_ _09190_/X _12003_/C _11939_/A vssd1 vssd1 vccd1 vccd1 _14791_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__09688__A _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12405__B1 _12404_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19378_ _19940_/CLK _19378_/D vssd1 vssd1 vccd1 vccd1 _19378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18329_ _17704_/X _19998_/Q _18335_/S vssd1 vssd1 vccd1 vccd1 _18330_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10967__B1 _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15629__S _15901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18005__S _18009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12842__A _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09964_ _10493_/S vssd1 vssd1 vccd1 vccd1 _10129_/S sky130_fd_sc_hd__buf_2
XFILLER_131_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09895_ _09895_/A vssd1 vssd1 vccd1 vccd1 _11554_/A sky130_fd_sc_hd__buf_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09983__S1 _09612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12892__B1 _12886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11542__S1 _09660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14708__S _14716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09598__A _09668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _10670_/A _10670_/B vssd1 vssd1 vccd1 vccd1 _10670_/X sky130_fd_sc_hd__or2_1
XFILLER_41_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ _18940_/Q _18985_/Q vssd1 vssd1 vccd1 vccd1 _09696_/A sky130_fd_sc_hd__or2b_1
XANTENNA__16923__S _16931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12340_ _12340_/A _12340_/B _12340_/C vssd1 vssd1 vccd1 vccd1 _12416_/D sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_98_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19966_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_154_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12271_ _12220_/A _12220_/B _12246_/A _12270_/X vssd1 vssd1 vccd1 vccd1 _12272_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_153_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16224__A _16691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14010_ _14010_/A _14010_/B vssd1 vssd1 vccd1 vccd1 _14010_/Y sky130_fd_sc_hd__nor2_1
X_11222_ _11291_/A _11222_/B vssd1 vssd1 vccd1 vccd1 _11222_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19855_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17754__S _17760_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11153_ _11153_/A vssd1 vssd1 vccd1 vccd1 _11154_/A sky130_fd_sc_hd__clkbuf_4
X_10104_ _10104_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _10104_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15961_ _19014_/Q _15954_/X _15955_/X _15960_/Y vssd1 vssd1 vccd1 vccd1 _19014_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11084_ _11340_/A vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17700_ _17700_/A vssd1 vssd1 vccd1 vccd1 _17700_/X sky130_fd_sc_hd__clkbuf_2
X_10035_ _19249_/Q _19744_/Q _10037_/S vssd1 vssd1 vccd1 vccd1 _10036_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18063__A1 _13591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14912_ _14912_/A vssd1 vssd1 vccd1 vccd1 _15160_/B sky130_fd_sc_hd__buf_2
XFILLER_76_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17055__A _17055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15892_ _15892_/A vssd1 vssd1 vccd1 vccd1 _18990_/D sky130_fd_sc_hd__clkbuf_1
X_18680_ _18687_/CLK _18680_/D vssd1 vssd1 vccd1 vccd1 _18680_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_36_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _20021_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17631_ _17631_/A vssd1 vssd1 vccd1 vccd1 _19717_/D sky130_fd_sc_hd__clkbuf_1
X_14843_ _15544_/A vssd1 vssd1 vccd1 vccd1 _15489_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output125_A _12856_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17562_ _17738_/B _17635_/A vssd1 vssd1 vccd1 vccd1 _17619_/A sky130_fd_sc_hd__or2_4
X_14774_ _14774_/A vssd1 vssd1 vccd1 vccd1 _18824_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11986_ _12174_/A _11981_/Y _11985_/X vssd1 vssd1 vccd1 vccd1 _12078_/C sky130_fd_sc_hd__o21a_1
X_16513_ _19240_/Q _13810_/X _16519_/S vssd1 vssd1 vccd1 vccd1 _16514_/A sky130_fd_sc_hd__mux2_1
X_19301_ _19636_/CLK _19301_/D vssd1 vssd1 vccd1 vccd1 _19301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13725_ _19022_/Q _13725_/B vssd1 vssd1 vccd1 vccd1 _13725_/X sky130_fd_sc_hd__or2_1
X_17493_ _17493_/A vssd1 vssd1 vccd1 vccd1 _19652_/D sky130_fd_sc_hd__clkbuf_1
X_10937_ _18433_/Q _19462_/Q _19499_/Q _19073_/Q _10703_/A _10709_/A vssd1 vssd1 vccd1
+ vccd1 _10937_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_152_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11831__A _11831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16444_ _19210_/Q _13816_/X _16446_/S vssd1 vssd1 vccd1 vccd1 _16445_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14388__B1 _14094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19232_ _20017_/CLK _19232_/D vssd1 vssd1 vccd1 vccd1 _19232_/Q sky130_fd_sc_hd__dfxtp_1
X_13656_ _13656_/A vssd1 vssd1 vccd1 vccd1 _13656_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10868_ _09702_/X _10850_/X _10867_/X _09843_/A _18844_/Q vssd1 vssd1 vccd1 vccd1
+ _12839_/B sky130_fd_sc_hd__a32o_4
XANTENNA__17929__S _17937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19163_ _20012_/CLK _19163_/D vssd1 vssd1 vccd1 vccd1 _19163_/Q sky130_fd_sc_hd__dfxtp_1
X_12607_ _12530_/X _12605_/Y _12606_/X _12583_/X vssd1 vssd1 vccd1 vccd1 _12607_/Y
+ sky130_fd_sc_hd__o31ai_2
X_16375_ _16374_/X _19183_/Q _16378_/S vssd1 vssd1 vccd1 vccd1 _16376_/A sky130_fd_sc_hd__mux2_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13587_ _13656_/A vssd1 vssd1 vccd1 vccd1 _13587_/X sky130_fd_sc_hd__clkbuf_2
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _19925_/Q _19539_/Q _19989_/Q _19108_/Q _10906_/S _10625_/A vssd1 vssd1 vccd1
+ vccd1 _10799_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18114_ _18858_/Q _13704_/X _18118_/S vssd1 vssd1 vccd1 vccd1 _18114_/X sky130_fd_sc_hd__mux2_1
X_15326_ _15243_/X _15314_/X _15325_/X _15258_/X vssd1 vssd1 vccd1 vccd1 _15326_/X
+ sky130_fd_sc_hd__o211a_1
X_19094_ _19975_/CLK _19094_/D vssd1 vssd1 vccd1 vccd1 _19094_/Q sky130_fd_sc_hd__dfxtp_1
X_12538_ _12634_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12539_/C sky130_fd_sc_hd__nor2_1
XFILLER_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18045_ _18045_/A vssd1 vssd1 vccd1 vccd1 _19885_/D sky130_fd_sc_hd__clkbuf_1
X_15257_ _15205_/X _15248_/X _15256_/X _15238_/X vssd1 vssd1 vccd1 vccd1 _15257_/X
+ sky130_fd_sc_hd__a211o_1
X_12469_ _12469_/A _12469_/B vssd1 vssd1 vccd1 vccd1 _12470_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__12662__A _15487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14208_ _14315_/A _14208_/B _14212_/C vssd1 vssd1 vccd1 vccd1 _18641_/D sky130_fd_sc_hd__nor3_1
XANTENNA__13363__A1 _13005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15188_ _15057_/X _15054_/X _15202_/S vssd1 vssd1 vccd1 vccd1 _15188_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11278__A _11278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14139_ _14142_/B _14142_/C _14102_/X vssd1 vssd1 vccd1 vccd1 _14139_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15104__A2 _15100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19996_ _19996_/CLK _19996_/D vssd1 vssd1 vccd1 vccd1 _19996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_77_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18947_ _18958_/CLK _18947_/D vssd1 vssd1 vccd1 vccd1 _18947_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14589__A _14595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18054__A1 _13563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ _19525_/Q vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18878_ _18878_/CLK _18878_/D vssd1 vssd1 vccd1 vccd1 _18878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17829_ _17829_/A vssd1 vssd1 vccd1 vccd1 _19790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14615__A1 _11724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15812__B1 _15798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11429__A1 _11291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11429__B2 _12895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15213__A _15393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15040__A1 _14966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17839__S _17843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16743__S _16747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11288__S0 _11125_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13668__A _18104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16044__A _16044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10168__A1 _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15883__A _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09881__A _09881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09947_ _18452_/Q _19481_/Q _19518_/Q _19092_/Q _09939_/X _09940_/X vssd1 vssd1 vccd1
+ vccd1 _09947_/X sky130_fd_sc_hd__mux4_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11117__B1 _11095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10820__A _10820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _09849_/X _09862_/X _09877_/X _09540_/X _18862_/Q vssd1 vssd1 vccd1 vccd1
+ _15978_/C sky130_fd_sc_hd__a32o_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16918__S _16918_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _15875_/A vssd1 vssd1 vccd1 vccd1 _11860_/A sky130_fd_sc_hd__buf_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11812_/B vssd1 vssd1 vccd1 vccd1 _17096_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _13510_/A _13510_/B vssd1 vssd1 vccd1 vccd1 _13511_/C sky130_fd_sc_hd__nor2_1
XFILLER_14_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _19669_/Q _19435_/Q _18500_/Q _19765_/Q _10764_/S _09606_/A vssd1 vssd1 vccd1
+ vccd1 _10723_/B sky130_fd_sc_hd__mux4_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14490_ _18729_/Q _14487_/B _14489_/Y vssd1 vssd1 vccd1 vccd1 _18729_/D sky130_fd_sc_hd__o21a_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13441_ _13223_/X _13426_/Y _13440_/X vssd1 vssd1 vccd1 vccd1 _17084_/A sky130_fd_sc_hd__o21ai_2
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17749__S _17749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10653_ _10653_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11279__S0 _11125_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16160_ _12978_/X _19099_/Q _16162_/S vssd1 vssd1 vccd1 vccd1 _16161_/A sky130_fd_sc_hd__mux2_1
X_13372_ _13188_/X _18858_/Q _12957_/X vssd1 vssd1 vccd1 vccd1 _13372_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10584_ _09883_/A _10570_/X _10582_/X _09913_/A _10583_/Y vssd1 vssd1 vccd1 vccd1
+ _12848_/B sky130_fd_sc_hd__o32a_4
XFILLER_70_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09892__S0 _09733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15111_ _15014_/X _15009_/X _15121_/S vssd1 vssd1 vccd1 vccd1 _15111_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12323_ _12323_/A _12323_/B _12323_/C _15291_/A vssd1 vssd1 vccd1 vccd1 _12406_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_127_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16091_ _16148_/S vssd1 vssd1 vccd1 vccd1 _16100_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_170_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15042_ _15094_/A vssd1 vssd1 vccd1 vccd1 _15199_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_170_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12254_ _12231_/A _12255_/C _18766_/Q vssd1 vssd1 vccd1 vccd1 _12254_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17484__S _17492_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11205_ _11283_/A _11205_/B vssd1 vssd1 vccd1 vccd1 _11205_/X sky130_fd_sc_hd__or2_1
XFILLER_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19850_ _19948_/CLK _19850_/D vssd1 vssd1 vccd1 vccd1 _19850_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10206__S _10469_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12185_ _12185_/A _12185_/B vssd1 vssd1 vccd1 vccd1 _12186_/B sky130_fd_sc_hd__and2_1
X_18801_ _19883_/CLK _18801_/D vssd1 vssd1 vccd1 vccd1 _18801_/Q sky130_fd_sc_hd__dfxtp_1
X_11136_ _18430_/Q _19459_/Q _19496_/Q _19070_/Q _10995_/X _11050_/A vssd1 vssd1 vccd1
+ vccd1 _11137_/B sky130_fd_sc_hd__mux4_1
X_19781_ _20039_/CLK _19781_/D vssd1 vssd1 vccd1 vccd1 _19781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16993_ _16993_/A _17954_/B vssd1 vssd1 vccd1 vccd1 _17075_/A sky130_fd_sc_hd__nor2_4
XFILLER_110_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18732_ _18734_/CLK _18732_/D vssd1 vssd1 vccd1 vccd1 _18732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11067_ _11283_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11067_/Y sky130_fd_sc_hd__nor2_1
X_15944_ _19008_/Q _15927_/X _15928_/X _15943_/Y vssd1 vssd1 vccd1 vccd1 _19008_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12320__A2 _12841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10867__C1 _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _10290_/A vssd1 vssd1 vccd1 vccd1 _10093_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15875_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15875_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18663_ _18731_/CLK _18663_/D vssd1 vssd1 vccd1 vccd1 _18663_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10331__A1 _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16828__S _16830_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17614_ _17614_/A vssd1 vssd1 vccd1 vccd1 _19709_/D sky130_fd_sc_hd__clkbuf_1
X_14826_ _14826_/A vssd1 vssd1 vccd1 vccd1 _15458_/A sky130_fd_sc_hd__buf_2
X_18594_ _18660_/CLK _18594_/D vssd1 vssd1 vccd1 vccd1 _18594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17545_ _17545_/A vssd1 vssd1 vccd1 vccd1 _19678_/D sky130_fd_sc_hd__clkbuf_1
X_14757_ _11660_/A _09520_/B _14756_/X vssd1 vssd1 vccd1 vccd1 _14764_/B sky130_fd_sc_hd__o21ai_1
X_11969_ _14865_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _12871_/A sky130_fd_sc_hd__and2_2
XFILLER_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13708_ _19020_/Q _13708_/B vssd1 vssd1 vccd1 vccd1 _13708_/X sky130_fd_sc_hd__or2_1
X_17476_ _17476_/A vssd1 vssd1 vccd1 vccd1 _19644_/D sky130_fd_sc_hd__clkbuf_1
X_14688_ _18796_/Q _13553_/X _14694_/S vssd1 vssd1 vccd1 vccd1 _14689_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10190__S0 _10449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19215_ _20030_/CLK _19215_/D vssd1 vssd1 vccd1 vccd1 _19215_/Q sky130_fd_sc_hd__dfxtp_1
X_16427_ _19202_/Q _13790_/X _16435_/S vssd1 vssd1 vccd1 vccd1 _16428_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15968__A _15982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13033__B1 _11794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13639_ _11724_/X _13638_/Y _13689_/S vssd1 vssd1 vccd1 vccd1 _13639_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10177__A _15974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16563__S _16569_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19146_ _19995_/CLK _19146_/D vssd1 vssd1 vccd1 vccd1 _19146_/Q sky130_fd_sc_hd__dfxtp_1
X_16358_ _17694_/A vssd1 vssd1 vccd1 vccd1 _16358_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09966__A _10180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15309_ _15282_/X _15415_/B _15308_/X _15238_/X vssd1 vssd1 vccd1 vccd1 _15309_/X
+ sky130_fd_sc_hd__a211o_1
X_19077_ _19990_/CLK _19077_/D vssd1 vssd1 vccd1 vccd1 _19077_/Q sky130_fd_sc_hd__dfxtp_1
X_16289_ _13443_/X _19156_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _16290_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12392__A _12416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13919__C _18606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18028_ _11845_/X _13511_/C _13518_/A vssd1 vssd1 vccd1 vccd1 _18028_/X sky130_fd_sc_hd__a21o_1
XFILLER_173_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17394__S _17398_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15907__S _15946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09801_ _19388_/Q vssd1 vssd1 vccd1 vccd1 _09802_/A sky130_fd_sc_hd__inv_2
XFILLER_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19979_ _19979_/CLK _19979_/D vssd1 vssd1 vccd1 vccd1 _19979_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14836__A1 _14966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18027__A1 _14554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09732_ _10094_/S vssd1 vssd1 vccd1 vccd1 _09950_/S sky130_fd_sc_hd__buf_2
XFILLER_68_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09663_ _11122_/A vssd1 vssd1 vccd1 vccd1 _09664_/A sky130_fd_sc_hd__buf_2
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09594_ _10447_/S vssd1 vssd1 vccd1 vccd1 _09595_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15261__A1 _18842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13272__B1 _12984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13162__S _13203_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__B1 _09837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17569__S _17573_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18254__A _18265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14782__A _14782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__A _09876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10389__A1 _10013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16513__A1 _13810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14524__B1 _14507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_100_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10236__S1 _10013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10561__A1 _09849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10561__B2 _18850_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ _18571_/Q _18570_/Q _13990_/C vssd1 vssd1 vccd1 vccd1 _13992_/B sky130_fd_sc_hd__and3_1
XFILLER_105_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _12941_/A vssd1 vssd1 vccd1 vccd1 _18425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16648__S _16652_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13861__A _14385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15660_ _18908_/Q _12340_/A _15666_/S vssd1 vssd1 vccd1 vccd1 _15661_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12872_ _19487_/Q vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__inv_2
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _18772_/Q _13629_/X _14615_/S vssd1 vssd1 vccd1 vccd1 _14612_/B sky130_fd_sc_hd__mux2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _18801_/Q _11841_/A _11817_/X _18768_/Q _11822_/X vssd1 vssd1 vccd1 vccd1
+ _11823_/X sky130_fd_sc_hd__a221o_2
XFILLER_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15591_ _15602_/A vssd1 vssd1 vccd1 vccd1 _15600_/S sky130_fd_sc_hd__buf_2
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17330_/A vssd1 vssd1 vccd1 vccd1 _19579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11381__A _11425_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14542_ input68/X _14544_/B vssd1 vssd1 vccd1 vccd1 _14542_/X sky130_fd_sc_hd__or2_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _18775_/Q vssd1 vssd1 vccd1 vccd1 _12508_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _17170_/X _19549_/Q _17265_/S vssd1 vssd1 vccd1 vccd1 _17262_/A sky130_fd_sc_hd__mux2_1
X_10705_ _19927_/Q _19541_/Q _19991_/Q _19110_/Q _10764_/S _09606_/A vssd1 vssd1 vccd1
+ vccd1 _10706_/B sky130_fd_sc_hd__mux4_1
XANTENNA__17479__S _17481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15788__A _15879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14473_ _18723_/Q _14470_/B _14472_/Y vssd1 vssd1 vccd1 vccd1 _18723_/D sky130_fd_sc_hd__o21a_1
X_11685_ _14227_/B _11790_/B vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__nor2_4
X_16212_ _16212_/A vssd1 vssd1 vccd1 vccd1 _19122_/D sky130_fd_sc_hd__clkbuf_1
X_19000_ _19001_/CLK _19000_/D vssd1 vssd1 vccd1 vccd1 _19000_/Q sky130_fd_sc_hd__dfxtp_2
X_13424_ _13423_/X _18451_/Q _13464_/S vssd1 vssd1 vccd1 vccd1 _13425_/A sky130_fd_sc_hd__mux2_1
X_10636_ _09777_/A _10628_/Y _10630_/Y _10633_/Y _10635_/Y vssd1 vssd1 vccd1 vccd1
+ _10636_/X sky130_fd_sc_hd__o32a_1
XFILLER_139_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17192_ _17729_/A vssd1 vssd1 vccd1 vccd1 _17192_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09865__S0 _09635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16143_ _16143_/A vssd1 vssd1 vccd1 vccd1 _19092_/D sky130_fd_sc_hd__clkbuf_1
X_13355_ _13354_/X _18447_/Q _13366_/S vssd1 vssd1 vccd1 vccd1 _13356_/A sky130_fd_sc_hd__mux2_1
X_10567_ _10567_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _10567_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10475__S1 _10473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__A _10919_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ _12479_/S _12304_/X _12305_/X _12056_/X vssd1 vssd1 vccd1 vccd1 _12306_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16074_ _16074_/A vssd1 vssd1 vccd1 vccd1 _19062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13286_ _18885_/Q vssd1 vssd1 vccd1 vccd1 _13664_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10498_ _19338_/Q _19609_/Q _19833_/Q _19577_/Q _10319_/A _10497_/X vssd1 vssd1 vccd1
+ vccd1 _10498_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10444__B _12851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15025_ _15021_/X _15024_/X _15198_/S vssd1 vssd1 vccd1 vccd1 _15025_/X sky130_fd_sc_hd__mux2_1
X_19902_ _19910_/CLK _19902_/D vssd1 vssd1 vccd1 vccd1 _19902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15835__A2_N _15834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12237_ _15234_/A _12323_/A _12322_/A vssd1 vssd1 vccd1 vccd1 _12238_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10227__S1 _10013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__S0 _11409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19833_ _19864_/CLK _19833_/D vssd1 vssd1 vccd1 vccd1 _19833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13755__B _17098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12168_ _18763_/Q _12167_/Y _12168_/S vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17942__S _17948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11119_ _18840_/Q vssd1 vssd1 vccd1 vccd1 _11119_/Y sky130_fd_sc_hd__inv_2
X_19764_ _19764_/CLK _19764_/D vssd1 vssd1 vccd1 vccd1 _19764_/Q sky130_fd_sc_hd__dfxtp_1
X_16976_ _16976_/A vssd1 vssd1 vccd1 vccd1 _19445_/D sky130_fd_sc_hd__clkbuf_1
X_12099_ _18458_/Q _12472_/A vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__or2_1
XFILLER_49_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18715_ _19883_/CLK _18715_/D vssd1 vssd1 vccd1 vccd1 _18715_/Q sky130_fd_sc_hd__dfxtp_1
Xinput6 io_dbus_rdata[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15927_ _15954_/A vssd1 vssd1 vccd1 vccd1 _15927_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15970__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19695_ _20017_/CLK _19695_/D vssd1 vssd1 vccd1 vccd1 _19695_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16558__S _16558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13771__A _17007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18646_ _18688_/CLK _18646_/D vssd1 vssd1 vccd1 vccd1 _18646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15858_ _15861_/A _17208_/B vssd1 vssd1 vccd1 vccd1 _15859_/A sky130_fd_sc_hd__and2_1
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14809_ _14993_/B vssd1 vssd1 vccd1 vccd1 _15004_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18577_ _19909_/CLK _18577_/D vssd1 vssd1 vccd1 vccd1 _18577_/Q sky130_fd_sc_hd__dfxtp_1
X_15789_ _15789_/A vssd1 vssd1 vccd1 vccd1 _15789_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13921__D _14099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11291__A _11291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17528_ _19670_/Q vssd1 vssd1 vccd1 vccd1 _17529_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17459_ _17144_/X _19637_/Q _17459_/S vssd1 vssd1 vccd1 vccd1 _17460_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16293__S _16295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09856__S0 _11532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12834__B _12844_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19129_ _19389_/CLK _19129_/D vssd1 vssd1 vccd1 vccd1 _19129_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15210__B _15219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14107__A _14143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10240__B1 _09913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13946__A _13946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__S0 _09586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12850__A _12851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13157__S _13359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17852__S _17854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09715_ _09946_/A vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__buf_2
XFILLER_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16468__S _16468_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09646_ _09646_/A vssd1 vssd1 vccd1 vccd1 _09647_/A sky130_fd_sc_hd__buf_2
XFILLER_71_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09577_ _10549_/A vssd1 vssd1 vccd1 vccd1 _10508_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16992__A _16992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10154__S0 _10152_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14716__S _14716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11470_ _09607_/A _11467_/X _11469_/X vssd1 vssd1 vccd1 vccd1 _11470_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10421_ _15960_/B vssd1 vssd1 vccd1 vccd1 _10444_/A sky130_fd_sc_hd__inv_2
XANTENNA__10457__S1 _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16931__S _16931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13140_ _13140_/A vssd1 vssd1 vccd1 vccd1 _18434_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12771__A2 _12012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10352_ _10352_/A _10352_/B vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__nor2_1
XFILLER_136_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10782__A1 _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17328__A _17339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ _13269_/A vssd1 vssd1 vccd1 vccd1 _13071_/X sky130_fd_sc_hd__clkbuf_2
X_10283_ _10283_/A vssd1 vssd1 vccd1 vccd1 _10283_/X sky130_fd_sc_hd__buf_2
XANTENNA__12760__A _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12022_ _12188_/A vssd1 vssd1 vccd1 vccd1 _13650_/A sky130_fd_sc_hd__buf_2
XANTENNA__13720__A1 _12422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input49_A io_ibus_inst[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16830_ _16393_/X _19381_/Q _16830_/S vssd1 vssd1 vccd1 vccd1 _16831_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16761_ _16761_/A vssd1 vssd1 vccd1 vccd1 _19350_/D sky130_fd_sc_hd__clkbuf_1
X_13973_ _18565_/Q _18564_/Q _13973_/C vssd1 vssd1 vccd1 vccd1 _13976_/B sky130_fd_sc_hd__and3_1
XANTENNA__16378__S _16378_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13484__B1 _13368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18500_ _19861_/CLK _18500_/D vssd1 vssd1 vccd1 vccd1 _18500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12924_ _12909_/X _18424_/Q _13003_/S vssd1 vssd1 vccd1 vccd1 _12925_/A sky130_fd_sc_hd__mux2_1
X_15712_ _18932_/Q _15740_/B vssd1 vssd1 vccd1 vccd1 _15712_/X sky130_fd_sc_hd__or2_1
X_16692_ _16692_/A _17882_/B vssd1 vssd1 vccd1 vccd1 _16749_/A sky130_fd_sc_hd__nor2_2
X_19480_ _19942_/CLK _19480_/D vssd1 vssd1 vccd1 vccd1 _19480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10393__S0 _10141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15225__A1 _18840_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18431_ _19950_/CLK _18431_/D vssd1 vssd1 vccd1 vccd1 _18431_/Q sky130_fd_sc_hd__dfxtp_1
X_12855_ _12857_/A _12855_/B vssd1 vssd1 vccd1 vccd1 _12855_/Y sky130_fd_sc_hd__nor2_4
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15643_ _15643_/A vssd1 vssd1 vccd1 vccd1 _18900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11806_ _15783_/B vssd1 vssd1 vccd1 vccd1 _15738_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18362_ _18362_/A vssd1 vssd1 vccd1 vccd1 _20012_/D sky130_fd_sc_hd__clkbuf_1
X_15574_ _13554_/A _18902_/Q _15578_/S vssd1 vssd1 vccd1 vccd1 _15575_/A sky130_fd_sc_hd__mux2_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12786_/A vssd1 vssd1 vccd1 vccd1 _12788_/A sky130_fd_sc_hd__inv_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _17141_/X _19572_/Q _17315_/S vssd1 vssd1 vccd1 vccd1 _17314_/A sky130_fd_sc_hd__mux2_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14525_ _14526_/B _14526_/C _14524_/Y vssd1 vssd1 vccd1 vccd1 _18742_/D sky130_fd_sc_hd__o21a_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _18599_/Q _11732_/X _11733_/X _18631_/Q _11736_/X vssd1 vssd1 vccd1 vccd1
+ _13245_/B sky130_fd_sc_hd__a221o_2
XANTENNA__10696__S1 _10010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18293_ _18350_/S vssd1 vssd1 vccd1 vccd1 _18302_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17002__S _17008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17244_ _17244_/A vssd1 vssd1 vccd1 vccd1 _19541_/D sky130_fd_sc_hd__clkbuf_1
X_14456_ _14459_/B _14459_/C _14427_/X vssd1 vssd1 vccd1 vccd1 _14456_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11668_ _11975_/A _11975_/B _11975_/C _11975_/D vssd1 vssd1 vccd1 vccd1 _12153_/C
+ sky130_fd_sc_hd__or4_2
X_13407_ _13406_/X _18450_/Q _13464_/S vssd1 vssd1 vccd1 vccd1 _13408_/A sky130_fd_sc_hd__mux2_1
X_17175_ _17175_/A vssd1 vssd1 vccd1 vccd1 _19513_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17937__S _17937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10619_ _11186_/S vssd1 vssd1 vccd1 vccd1 _10892_/A sky130_fd_sc_hd__buf_2
XFILLER_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14387_ _18692_/Q vssd1 vssd1 vccd1 vccd1 _14390_/A sky130_fd_sc_hd__inv_2
X_11599_ _11599_/A _11599_/B vssd1 vssd1 vccd1 vccd1 _11600_/B sky130_fd_sc_hd__nand2_1
X_16126_ _16126_/A vssd1 vssd1 vccd1 vccd1 _19084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13338_ _13360_/A _18855_/Q vssd1 vssd1 vccd1 vccd1 _13338_/X sky130_fd_sc_hd__or2_1
XFILLER_143_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16057_ _13501_/X _19057_/Q _16057_/S vssd1 vssd1 vccd1 vccd1 _16058_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09963__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ _13269_/A vssd1 vssd1 vccd1 vccd1 _13269_/X sky130_fd_sc_hd__buf_2
XFILLER_170_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ _15405_/A vssd1 vssd1 vccd1 vccd1 _15428_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13711__A1 _13710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__B1 _09913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19816_ _19816_/CLK _19816_/D vssd1 vssd1 vccd1 vccd1 _19816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19747_ _19747_/CLK _19747_/D vssd1 vssd1 vccd1 vccd1 _19747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16959_ _16959_/A vssd1 vssd1 vccd1 vccd1 _19437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14597__A _14648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09500_ _11961_/B _09500_/B vssd1 vssd1 vccd1 vccd1 _11956_/B sky130_fd_sc_hd__or2_1
XFILLER_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19678_ _20032_/CLK _19678_/D vssd1 vssd1 vccd1 vccd1 _19678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09431_ _15624_/A vssd1 vssd1 vccd1 vccd1 _15914_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18629_ _18731_/CLK _18629_/D vssd1 vssd1 vccd1 vccd1 _18629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17701__A _17717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09362_ _18752_/Q _18747_/Q vssd1 vssd1 vccd1 vccd1 _09362_/X sky130_fd_sc_hd__and2_1
XANTENNA__14975__B1 _15940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09293_ _18937_/Q vssd1 vssd1 vccd1 vccd1 _09322_/A sky130_fd_sc_hd__inv_2
XFILLER_32_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12450__A1 _12338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16317__A _16400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10439__S1 _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17148__A _17180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput140 _12836_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[9] sky130_fd_sc_hd__buf_2
Xoutput151 _12510_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[18] sky130_fd_sc_hd__buf_2
XFILLER_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput162 _12752_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[28] sky130_fd_sc_hd__buf_2
XFILLER_82_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13395__B _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput173 _12259_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[9] sky130_fd_sc_hd__buf_2
XFILLER_114_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11908__B _14771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17582__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10611__S1 _09607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16652__A0 _16345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15455__A1 _12599_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16198__S _16206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10970_ _11325_/A vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__buf_2
XFILLER_56_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ _10369_/A vssd1 vssd1 vccd1 vccd1 _09973_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _12640_/A _12640_/B vssd1 vssd1 vccd1 vccd1 _12729_/A sky130_fd_sc_hd__and2_2
XFILLER_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ _12571_/A _14863_/A vssd1 vssd1 vccd1 vccd1 _12572_/B sky130_fd_sc_hd__or2_1
XANTENNA__16227__A _16295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14310_ _14316_/B _14317_/D _14203_/X vssd1 vssd1 vccd1 vccd1 _14310_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13350__S _13350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ _11522_/A vssd1 vssd1 vccd1 vccd1 _11522_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12992__A2 _12889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15290_ _15284_/X _15285_/Y _15289_/X _15268_/X vssd1 vssd1 vccd1 vccd1 _15293_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14241_ _18649_/Q _14241_/B vssd1 vssd1 vccd1 vccd1 _14244_/B sky130_fd_sc_hd__nor2_1
X_11453_ _11408_/X _11607_/A _11611_/A vssd1 vssd1 vccd1 vccd1 _11453_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16661__S _16663_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__A _10275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ _10400_/X _10402_/X _10403_/X _10191_/A _09565_/A vssd1 vssd1 vccd1 vccd1
+ _10409_/B sky130_fd_sc_hd__o221a_1
XFILLER_109_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14172_ _18629_/Q _18628_/Q _14172_/C vssd1 vssd1 vccd1 vccd1 _14174_/B sky130_fd_sc_hd__and3_1
X_11384_ _11377_/Y _11379_/Y _11381_/Y _11383_/Y _19526_/Q vssd1 vssd1 vccd1 vccd1
+ _11384_/X sky130_fd_sc_hd__o221a_1
XFILLER_124_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13123_ _18464_/Q _12982_/A _11847_/A _14378_/B _13122_/X vssd1 vssd1 vccd1 vccd1
+ _13123_/X sky130_fd_sc_hd__a221o_1
XANTENNA__17058__A _17058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10335_ _10335_/A _10335_/B vssd1 vssd1 vccd1 vccd1 _10335_/X sky130_fd_sc_hd__or2_1
XFILLER_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18980_ _19526_/CLK _18980_/D vssd1 vssd1 vccd1 vccd1 _18980_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12490__A _15397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _19836_/Q _17062_/X _17937_/S vssd1 vssd1 vccd1 vccd1 _17932_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _18557_/Q _13054_/B vssd1 vssd1 vccd1 vccd1 _13054_/X sky130_fd_sc_hd__or2_1
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10266_ _10266_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10266_/X sky130_fd_sc_hd__or2_1
XFILLER_87_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output155_A _12585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17492__S _17492_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ _18520_/Q _15633_/D vssd1 vssd1 vccd1 vccd1 _12052_/B sky130_fd_sc_hd__and2_1
X_17862_ _17862_/A vssd1 vssd1 vccd1 vccd1 _19805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10602__S1 _10654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ _18450_/Q _19479_/Q _19516_/Q _19090_/Q _10313_/S _10182_/X vssd1 vssd1 vccd1
+ vccd1 _10197_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19601_ _19856_/CLK _19601_/D vssd1 vssd1 vccd1 vccd1 _19601_/Q sky130_fd_sc_hd__dfxtp_1
X_16813_ _16368_/X _19373_/Q _16819_/S vssd1 vssd1 vccd1 vccd1 _16814_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17793_ _17713_/X _19775_/Q _17793_/S vssd1 vssd1 vccd1 vccd1 _17794_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19532_ _19982_/CLK _19532_/D vssd1 vssd1 vccd1 vccd1 _19532_/Q sky130_fd_sc_hd__dfxtp_1
X_16744_ _16744_/A vssd1 vssd1 vccd1 vccd1 _19342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14210__A _14239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ _18559_/Q _13956_/B _13956_/C vssd1 vssd1 vccd1 vccd1 _13957_/C sky130_fd_sc_hd__and3_1
XANTENNA__12141__A2_N _12830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19463_ _20018_/CLK _19463_/D vssd1 vssd1 vccd1 vccd1 _19463_/Q sky130_fd_sc_hd__dfxtp_1
X_12907_ _12874_/X _12898_/X _12902_/X input1/X _12906_/X vssd1 vssd1 vccd1 vccd1
+ _16992_/A sky130_fd_sc_hd__a32o_4
X_16675_ _16675_/A vssd1 vssd1 vccd1 vccd1 _19312_/D sky130_fd_sc_hd__clkbuf_1
X_13887_ _12377_/A _12377_/B _14447_/B vssd1 vssd1 vccd1 vccd1 _18531_/D sky130_fd_sc_hd__a21o_1
XFILLER_35_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18414_ _17723_/X _20036_/Q _18418_/S vssd1 vssd1 vccd1 vccd1 _18415_/A sky130_fd_sc_hd__mux2_1
X_12838_ _12838_/A vssd1 vssd1 vccd1 vccd1 _12838_/X sky130_fd_sc_hd__clkbuf_1
X_15626_ _15626_/A vssd1 vssd1 vccd1 vccd1 _18893_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19394_ _19758_/CLK _19394_/D vssd1 vssd1 vccd1 vccd1 _19394_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10118__S0 _09595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18345_ _18345_/A vssd1 vssd1 vccd1 vccd1 _20005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ _15236_/A _15555_/X _15556_/Y _15400_/A vssd1 vssd1 vccd1 vccd1 _15557_/X
+ sky130_fd_sc_hd__a31o_1
X_12769_ _12769_/A _12793_/B vssd1 vssd1 vccd1 vccd1 _12769_/X sky130_fd_sc_hd__or2_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12983__A2 _11845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14508_ _14510_/B _14510_/C _14507_/X vssd1 vssd1 vccd1 vccd1 _14508_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_159_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18276_ _19975_/Q _17732_/A _18278_/S vssd1 vssd1 vccd1 vccd1 _18277_/A sky130_fd_sc_hd__mux2_1
X_15488_ _15142_/A _15483_/Y _15487_/Y vssd1 vssd1 vccd1 vccd1 _15489_/C sky130_fd_sc_hd__a21oi_1
XFILLER_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 io_dbus_rdata[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_4
X_17227_ _17227_/A vssd1 vssd1 vccd1 vccd1 _19533_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15976__A _15978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14439_ _18707_/Q _18706_/Q _14439_/C vssd1 vssd1 vccd1 vccd1 _14440_/C sky130_fd_sc_hd__and3_1
Xinput31 io_dbus_rdata[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
Xinput42 io_ibus_inst[17] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_2
Xinput53 io_ibus_inst[27] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 io_ibus_inst[8] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_6
XANTENNA__18320__A0 _17691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17158_ _17157_/X _19508_/Q _17161_/S vssd1 vssd1 vccd1 vccd1 _17159_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11094__S1 _11022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16109_ _13180_/X _19077_/Q _16111_/S vssd1 vssd1 vccd1 vccd1 _16110_/A sky130_fd_sc_hd__mux2_1
X_09980_ _09980_/A vssd1 vssd1 vccd1 vccd1 _09980_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17089_ _17089_/A vssd1 vssd1 vccd1 vccd1 _19482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11728__B _15715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_147_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11463__B _12839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09414_ _15779_/A _09411_/Y _09412_/X _15777_/A vssd1 vssd1 vccd1 vccd1 _09414_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14948__A0 _15474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09345_ _09345_/A vssd1 vssd1 vccd1 vccd1 _15633_/A sky130_fd_sc_hd__buf_2
XFILLER_34_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _14755_/A _09514_/A _09276_/C vssd1 vssd1 vccd1 vccd1 _09276_/X sky130_fd_sc_hd__or3_4
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14790__A _15762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09884__A _09884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10120_ _10107_/X _10111_/Y _10114_/Y _10117_/Y _10119_/Y vssd1 vssd1 vccd1 vccd1
+ _10120_/X sky130_fd_sc_hd__o32a_1
XFILLER_122_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10051_ _10587_/A vssd1 vssd1 vccd1 vccd1 _10398_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15979__A2 _14803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13345__S _13366_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13810_ _17046_/A vssd1 vssd1 vccd1 vccd1 _13810_/X sky130_fd_sc_hd__clkbuf_2
X_14790_ _15762_/A vssd1 vssd1 vccd1 vccd1 _15740_/B sky130_fd_sc_hd__buf_2
XFILLER_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ _19024_/Q _13472_/X _13740_/Y _11717_/X vssd1 vssd1 vccd1 vccd1 _13741_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10953_ _19361_/Q _19696_/Q _10953_/S vssd1 vssd1 vccd1 vccd1 _10953_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16460_ _19217_/Q _13838_/X _16468_/S vssd1 vssd1 vccd1 vccd1 _16461_/A sky130_fd_sc_hd__mux2_1
X_13672_ _18885_/Q _18886_/Q _13672_/C vssd1 vssd1 vccd1 vccd1 _13681_/B sky130_fd_sc_hd__or3_1
X_10884_ _10727_/A _10883_/X _10712_/A vssd1 vssd1 vccd1 vccd1 _10884_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12623_ _18540_/Q _18541_/Q _12623_/C vssd1 vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__and3_1
X_15411_ _15159_/X _15406_/Y _15410_/Y vssd1 vssd1 vccd1 vccd1 _15412_/C sky130_fd_sc_hd__a21oi_1
X_16391_ _16390_/X _19188_/Q _16394_/S vssd1 vssd1 vccd1 vccd1 _16392_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18130_ _18863_/Q _13742_/X _18130_/S vssd1 vssd1 vccd1 vccd1 _18130_/X sky130_fd_sc_hd__mux2_1
X_15342_ _15428_/A vssd1 vssd1 vccd1 vccd1 _15342_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12554_ _12554_/A _12576_/C vssd1 vssd1 vccd1 vccd1 _12554_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_129_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11505_ _09793_/A _11498_/Y _11500_/Y _11502_/Y _11504_/Y vssd1 vssd1 vccd1 vccd1
+ _11505_/X sky130_fd_sc_hd__o32a_1
XFILLER_129_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15796__A _15807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18061_ _18060_/X _19890_/Q _18061_/S vssd1 vssd1 vccd1 vccd1 _18062_/A sky130_fd_sc_hd__mux2_1
X_15273_ _15205_/X _15440_/B _15272_/X _15238_/X vssd1 vssd1 vccd1 vccd1 _15273_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10209__S _10209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16391__S _16394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12485_ _12501_/A _12415_/X _12481_/X _12484_/Y vssd1 vssd1 vccd1 vccd1 _12485_/X
+ sky130_fd_sc_hd__o22a_4
XANTENNA__16150__C_N _15735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14224_ _15779_/A _15777_/A _18942_/Q _18941_/Q vssd1 vssd1 vccd1 vccd1 _14226_/B
+ sky130_fd_sc_hd__or4_1
X_17012_ _19458_/Q _17010_/X _17024_/S vssd1 vssd1 vccd1 vccd1 _17013_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11436_ _19192_/Q _19783_/Q _19945_/Q _19160_/Q _10960_/A _11388_/A vssd1 vssd1 vccd1
+ vccd1 _11436_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10728__A1 _09664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11829__A _14552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ _14245_/A vssd1 vssd1 vccd1 vccd1 _14191_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11367_ _19353_/Q _19688_/Q _11367_/S vssd1 vssd1 vccd1 vccd1 _11367_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10823__S1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13106_ _18591_/Q _13057_/A _12890_/A _18723_/Q vssd1 vssd1 vccd1 vccd1 _13106_/X
+ sky130_fd_sc_hd__a22o_1
X_10318_ _10543_/S vssd1 vssd1 vccd1 vccd1 _10319_/A sky130_fd_sc_hd__buf_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14086_ _18605_/Q _14086_/B _14086_/C vssd1 vssd1 vccd1 vccd1 _14088_/B sky130_fd_sc_hd__and3_1
X_18963_ _18967_/CLK _18963_/D vssd1 vssd1 vccd1 vccd1 _18963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _11309_/A _11297_/X _09772_/A vssd1 vssd1 vccd1 vccd1 _11298_/Y sky130_fd_sc_hd__o21ai_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _17914_/A vssd1 vssd1 vccd1 vccd1 _19828_/D sky130_fd_sc_hd__clkbuf_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _18839_/Q _13551_/B _13349_/S vssd1 vssd1 vccd1 vccd1 _13037_/X sky130_fd_sc_hd__mux2_1
X_10249_ _15968_/B _12856_/B vssd1 vssd1 vccd1 vccd1 _11635_/A sky130_fd_sc_hd__xnor2_1
XFILLER_121_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15962__C _15962_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18894_ _18928_/CLK _18894_/D vssd1 vssd1 vccd1 vccd1 _18894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17845_ _17867_/A vssd1 vssd1 vccd1 vccd1 _17854_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_120_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17950__S _17952_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17776_ _17688_/X _19767_/Q _17782_/S vssd1 vssd1 vccd1 vccd1 _17777_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14988_ _15041_/S vssd1 vssd1 vccd1 vccd1 _15055_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_75_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19515_ _20034_/CLK _19515_/D vssd1 vssd1 vccd1 vccd1 _19515_/Q sky130_fd_sc_hd__dfxtp_1
X_16727_ _16749_/A vssd1 vssd1 vccd1 vccd1 _16736_/S sky130_fd_sc_hd__clkbuf_4
X_13939_ _13947_/D vssd1 vssd1 vccd1 vccd1 _13945_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14875__A _14931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19446_ _19873_/CLK _19446_/D vssd1 vssd1 vccd1 vccd1 _19446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16658_ _16658_/A vssd1 vssd1 vccd1 vccd1 _19304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15609_ _13306_/X _18918_/Q _15611_/S vssd1 vssd1 vccd1 vccd1 _15610_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12405__A1 _11904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19377_ _19873_/CLK _19377_/D vssd1 vssd1 vccd1 vccd1 _19377_/Q sky130_fd_sc_hd__dfxtp_1
X_16589_ _19274_/Q _13816_/X _16591_/S vssd1 vssd1 vccd1 vccd1 _16590_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_73_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18328_ _18328_/A vssd1 vssd1 vccd1 vccd1 _19997_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10967__A1 _09702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10967__B2 _18842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18259_ _19967_/Q _17707_/A _18263_/S vssd1 vssd1 vccd1 vccd1 _18260_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12842__B _12844_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19980_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09963_ _15976_/C _12862_/B vssd1 vssd1 vccd1 vccd1 _11644_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09209__A _19488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13954__A _14094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09894_ _09887_/Y _09889_/Y _09891_/Y _09893_/Y _11574_/A vssd1 vssd1 vccd1 vccd1
+ _09894_/X sky130_fd_sc_hd__o221a_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15830__A1 hold4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15830__B2 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09328_ _18984_/Q vssd1 vssd1 vccd1 vccd1 _09328_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09259_ _18987_/Q vssd1 vssd1 vccd1 vccd1 _09261_/A sky130_fd_sc_hd__buf_4
XFILLER_138_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12270_ _12244_/X _12241_/X _12243_/B vssd1 vssd1 vccd1 vccd1 _12270_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16224__B _16691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11221_ _11214_/Y _11216_/Y _11218_/Y _11220_/Y _09549_/A vssd1 vssd1 vccd1 vccd1
+ _11222_/B sky130_fd_sc_hd__o221a_1
XANTENNA__13372__A2 _18858_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10553__A _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11152_ _11145_/Y _11147_/Y _11149_/Y _11151_/Y _11166_/A vssd1 vssd1 vccd1 vccd1
+ _11152_/X sky130_fd_sc_hd__o221a_1
XFILLER_150_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10103_ _09884_/X _10091_/X _10102_/X _09913_/X _10079_/Y vssd1 vssd1 vccd1 vccd1
+ _12856_/B sky130_fd_sc_hd__o32a_4
XFILLER_1_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13124__A2 _13071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13864__A _14577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15960_ _15964_/A _15960_/B vssd1 vssd1 vccd1 vccd1 _15960_/Y sky130_fd_sc_hd__nor2_1
X_11083_ _11111_/A vssd1 vssd1 vccd1 vccd1 _11340_/A sky130_fd_sc_hd__buf_2
XFILLER_49_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input31_A io_dbus_rdata[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _19680_/Q _19446_/Q _18511_/Q _19776_/Q _10277_/S _10082_/A vssd1 vssd1 vccd1
+ vccd1 _10034_/X sky130_fd_sc_hd__mux4_1
X_14911_ _14908_/X _14910_/X _15032_/S vssd1 vssd1 vccd1 vccd1 _14911_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15891_ _15897_/A _15891_/B vssd1 vssd1 vccd1 vccd1 _15892_/A sky130_fd_sc_hd__and2_1
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17630_ _17195_/X _19717_/Q _17632_/S vssd1 vssd1 vccd1 vccd1 _17631_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14842_ _15444_/A vssd1 vssd1 vccd1 vccd1 _15544_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15821__A1 hold2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15821__B2 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17561_ _17561_/A vssd1 vssd1 vccd1 vccd1 _19686_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12635__A1 _09466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14773_ _14780_/A _14773_/B vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__and2_1
X_11985_ _09495_/A _11984_/X _09319_/A vssd1 vssd1 vccd1 vccd1 _11985_/X sky130_fd_sc_hd__a21o_1
XANTENNA_output118_A _12849_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19300_ _19989_/CLK _19300_/D vssd1 vssd1 vccd1 vccd1 _19300_/Q sky130_fd_sc_hd__dfxtp_1
X_16512_ _16512_/A vssd1 vssd1 vccd1 vccd1 _19239_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17071__A _17071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10936_ _10936_/A _10936_/B vssd1 vssd1 vccd1 vccd1 _10936_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13724_ _13737_/C _13723_/Y _13700_/X vssd1 vssd1 vccd1 vccd1 _13724_/Y sky130_fd_sc_hd__a21oi_1
X_17492_ _17192_/X _19652_/Q _17492_/S vssd1 vssd1 vccd1 vccd1 _17493_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19231_ _19726_/CLK _19231_/D vssd1 vssd1 vccd1 vccd1 _19231_/Q sky130_fd_sc_hd__dfxtp_1
X_16443_ _16443_/A vssd1 vssd1 vccd1 vccd1 _19209_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10867_ _09776_/A _10858_/X _10862_/X _10866_/X _09819_/A vssd1 vssd1 vccd1 vccd1
+ _10867_/X sky130_fd_sc_hd__a311o_2
X_13655_ _13672_/C _13654_/Y _13648_/X vssd1 vssd1 vccd1 vccd1 _13655_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_20_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09301__B _18938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19162_ _19979_/CLK _19162_/D vssd1 vssd1 vccd1 vccd1 _19162_/Q sky130_fd_sc_hd__dfxtp_1
X_12606_ _18779_/Q _12628_/C vssd1 vssd1 vccd1 vccd1 _12606_/X sky130_fd_sc_hd__and2_1
X_16374_ _17710_/A vssd1 vssd1 vccd1 vccd1 _16374_/X sky130_fd_sc_hd__clkbuf_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _13586_/A vssd1 vssd1 vccd1 vccd1 _18463_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13060__A1 _18653_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _18436_/Q _19465_/Q _19502_/Q _19076_/Q _10797_/X _10793_/X vssd1 vssd1 vccd1
+ vccd1 _10798_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18113_ _18113_/A vssd1 vssd1 vccd1 vccd1 _19905_/D sky130_fd_sc_hd__clkbuf_1
X_12537_ _12537_/A vssd1 vssd1 vccd1 vccd1 _12634_/A sky130_fd_sc_hd__clkbuf_2
X_15325_ _15282_/X _15315_/X _15323_/X _15324_/X vssd1 vssd1 vccd1 vccd1 _15325_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19093_ _19747_/CLK _19093_/D vssd1 vssd1 vccd1 vccd1 _19093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12943__A _12943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16415__A _16472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18044_ hold5/X _19885_/Q _18044_/S vssd1 vssd1 vccd1 vccd1 _18045_/A sky130_fd_sc_hd__mux2_1
X_12468_ _12437_/A _15373_/B _12442_/A _12442_/B vssd1 vssd1 vccd1 vccd1 _12469_/B
+ sky130_fd_sc_hd__a22o_1
X_15256_ _15323_/A _15256_/B _15256_/C vssd1 vssd1 vccd1 vccd1 _15256_/X sky130_fd_sc_hd__and3_1
XFILLER_126_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11419_ _11058_/A _11412_/Y _11414_/Y _11418_/Y _09872_/A vssd1 vssd1 vccd1 vccd1
+ _11419_/X sky130_fd_sc_hd__o311a_1
X_14207_ _18641_/Q _18640_/Q _14207_/C vssd1 vssd1 vccd1 vccd1 _14212_/C sky130_fd_sc_hd__and3_2
X_15187_ _15489_/A _15182_/X _15186_/Y _15005_/X vssd1 vssd1 vccd1 vccd1 _15187_/X
+ sky130_fd_sc_hd__a211o_1
X_12399_ _12399_/A _12424_/C vssd1 vssd1 vccd1 vccd1 _12399_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14138_ _18618_/Q _14134_/C _14137_/Y vssd1 vssd1 vccd1 vccd1 _18618_/D sky130_fd_sc_hd__o21a_1
X_19995_ _19995_/CLK _19995_/D vssd1 vssd1 vccd1 vccd1 _19995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10582__C1 _09806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13774__A _17010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14069_ _14070_/B _14070_/C _14068_/Y vssd1 vssd1 vccd1 vccd1 _18598_/D sky130_fd_sc_hd__o21a_1
XFILLER_98_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18946_ _18967_/CLK _18946_/D vssd1 vssd1 vccd1 vccd1 _18946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16150__A _16474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18877_ _18878_/CLK _18877_/D vssd1 vssd1 vccd1 vccd1 _18877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17828_ _19790_/Q _17017_/X _17832_/S vssd1 vssd1 vccd1 vccd1 _17829_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17759_ _17759_/A vssd1 vssd1 vccd1 vccd1 _19759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12837__B _12837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19429_ _20015_/CLK _19429_/D vssd1 vssd1 vccd1 vccd1 _19429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10638__A _10638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13051__B2 _18461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__S1 _11077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13949__A _13967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18016__S _18020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__A _12857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13339__C1 _13289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_150_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _18677_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10799__S0 _10906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09946_ _09946_/A _09946_/B vssd1 vssd1 vccd1 vccd1 _09946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_165_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _18960_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09877_ _09864_/X _09866_/X _09868_/X _09870_/X _09876_/X vssd1 vssd1 vccd1 vccd1
+ _09877_/X sky130_fd_sc_hd__a221o_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16995__A _17094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _12060_/A _11770_/B _15777_/A vssd1 vssd1 vccd1 vccd1 _11812_/B sky130_fd_sc_hd__or3b_2
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10706_/Y _10713_/Y _10715_/Y _10720_/Y _09551_/A vssd1 vssd1 vccd1 vccd1
+ _10721_/X sky130_fd_sc_hd__o221a_2
XANTENNA__15567__A0 _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16934__S _16942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13440_ _13307_/X _13429_/X _13430_/Y _13439_/Y _09532_/A vssd1 vssd1 vccd1 vccd1
+ _13440_/X sky130_fd_sc_hd__a221o_1
X_10652_ _10652_/A _12847_/B vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_103_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _20032_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11279__S1 _11065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13371_ _13699_/A _13390_/C vssd1 vssd1 vccd1 vccd1 _13371_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ _18850_/Q vssd1 vssd1 vccd1 vccd1 _10583_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09892__S1 _09768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15110_ _15011_/X _15022_/X _15113_/S vssd1 vssd1 vccd1 vccd1 _15110_/X sky130_fd_sc_hd__mux2_1
X_12322_ _12322_/A vssd1 vssd1 vccd1 vccd1 _12459_/A sky130_fd_sc_hd__buf_2
XANTENNA__10800__B1 _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16090_ _16090_/A vssd1 vssd1 vccd1 vccd1 _19068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13578__B _19003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17765__S _17771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15041_ _15039_/X _15040_/Y _15041_/S vssd1 vssd1 vccd1 vccd1 _15041_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12253_ _14744_/B vssd1 vssd1 vccd1 vccd1 _12344_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10283__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_118_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19973_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11204_ _19132_/Q _19393_/Q _19292_/Q _19627_/Q _11063_/X _11065_/X vssd1 vssd1 vccd1
+ vccd1 _11205_/B sky130_fd_sc_hd__mux4_1
XFILLER_135_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12184_ _12184_/A _12150_/A vssd1 vssd1 vccd1 vccd1 _12185_/B sky130_fd_sc_hd__or2b_1
XFILLER_162_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18800_ _19883_/CLK _18800_/D vssd1 vssd1 vccd1 vccd1 _18800_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_21_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11135_ _11252_/A _11135_/B vssd1 vssd1 vccd1 vccd1 _11135_/X sky130_fd_sc_hd__or2_1
X_19780_ _19842_/CLK _19780_/D vssd1 vssd1 vccd1 vccd1 _19780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16992_ _16992_/A vssd1 vssd1 vccd1 vccd1 _16992_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12305__B1 _12301_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18731_ _18731_/CLK _18731_/D vssd1 vssd1 vccd1 vccd1 _18731_/Q sky130_fd_sc_hd__dfxtp_1
X_15943_ _15964_/A _15943_/B vssd1 vssd1 vccd1 vccd1 _15943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11066_ _19920_/Q _19534_/Q _19984_/Q _19103_/Q _11063_/X _11065_/X vssd1 vssd1 vccd1
+ vccd1 _11067_/B sky130_fd_sc_hd__mux4_1
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11318__S _11367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10017_ _10380_/A vssd1 vssd1 vccd1 vccd1 _10290_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18662_ _18731_/CLK _18662_/D vssd1 vssd1 vccd1 vccd1 _18662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15874_ _15874_/A vssd1 vssd1 vccd1 vccd1 _18985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17613_ _17170_/X _19709_/Q _17617_/S vssd1 vssd1 vccd1 vccd1 _17614_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14825_ _15048_/A vssd1 vssd1 vccd1 vccd1 _14826_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12608__A1 _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18593_ _18724_/CLK _18593_/D vssd1 vssd1 vccd1 vccd1 _18593_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12938__A _16998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17005__S _17008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17544_ _19678_/Q vssd1 vssd1 vccd1 vccd1 _17545_/A sky130_fd_sc_hd__clkbuf_1
X_14756_ _14756_/A _14756_/B vssd1 vssd1 vccd1 vccd1 _14756_/X sky130_fd_sc_hd__or2_1
XFILLER_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11968_ _11967_/Y _18897_/Q _12039_/A vssd1 vssd1 vccd1 vccd1 _12870_/B sky130_fd_sc_hd__mux2_4
XANTENNA__10714__S0 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13707_ _13714_/A _13714_/C vssd1 vssd1 vccd1 vccd1 _13707_/Y sky130_fd_sc_hd__xnor2_1
X_17475_ _17167_/X _19644_/Q _17481_/S vssd1 vssd1 vccd1 vccd1 _17476_/A sky130_fd_sc_hd__mux2_1
X_10919_ _19233_/Q _19728_/Q _10919_/S vssd1 vssd1 vccd1 vccd1 _10920_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10458__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14687_ _14687_/A vssd1 vssd1 vccd1 vccd1 _18795_/D sky130_fd_sc_hd__clkbuf_1
X_11899_ _11773_/A _11898_/X _11812_/B vssd1 vssd1 vccd1 vccd1 _11899_/X sky130_fd_sc_hd__a21bo_1
X_19214_ _19935_/CLK _19214_/D vssd1 vssd1 vccd1 vccd1 _19214_/Q sky130_fd_sc_hd__dfxtp_1
X_16426_ _16472_/S vssd1 vssd1 vccd1 vccd1 _16435_/S sky130_fd_sc_hd__buf_4
XFILLER_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13638_ _13646_/C _13638_/B vssd1 vssd1 vccd1 vccd1 _13638_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__10177__B _12860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19145_ _19641_/CLK _19145_/D vssd1 vssd1 vccd1 vccd1 _19145_/Q sky130_fd_sc_hd__dfxtp_1
X_16357_ _16357_/A vssd1 vssd1 vccd1 vccd1 _19177_/D sky130_fd_sc_hd__clkbuf_1
X_13569_ _13569_/A vssd1 vssd1 vccd1 vccd1 _18461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15308_ _15323_/A _15308_/B _15308_/C vssd1 vssd1 vccd1 vccd1 _15308_/X sky130_fd_sc_hd__and3_1
X_19076_ _19633_/CLK _19076_/D vssd1 vssd1 vccd1 vccd1 _19076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16288_ _16288_/A vssd1 vssd1 vccd1 vccd1 _19155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15984__A _17098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18027_ _09347_/X _14554_/X _18050_/S vssd1 vssd1 vccd1 vccd1 _18027_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13336__A2 _09402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14533__B2 _14548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15239_ _15205_/X _15229_/X _15236_/X _15238_/X vssd1 vssd1 vccd1 vccd1 _15239_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13741__C1 _11717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09800_ _09750_/A _09786_/X _09809_/A vssd1 vssd1 vccd1 vccd1 _09800_/X sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_82_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _20028_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19978_ _19978_/CLK _19978_/D vssd1 vssd1 vccd1 vccd1 _19978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09731_ _10277_/S vssd1 vssd1 vccd1 vccd1 _10094_/S sky130_fd_sc_hd__buf_2
X_18929_ _18967_/CLK _18929_/D vssd1 vssd1 vccd1 vccd1 _18929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09662_ _11199_/A vssd1 vssd1 vccd1 vccd1 _11122_/A sky130_fd_sc_hd__buf_2
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_97_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19644_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09593_ _10493_/S vssd1 vssd1 vccd1 vccd1 _10447_/S sky130_fd_sc_hd__buf_2
XANTENNA__12848__A _12851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15261__A2 _09433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10705__S0 _10764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_clock clkbuf_opt_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _18851_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16754__S _16758_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11822__A2 _13290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14772__B2 _13531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12583__A _12583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11130__S0 _11270_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19633_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11199__A _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10546__C1 _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_195_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09929_ _09929_/A _09929_/B vssd1 vssd1 vccd1 vccd1 _09929_/X sky130_fd_sc_hd__or2_1
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12919__B1_N _16846_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16929__S _16931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11197__S0 _11125_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12940_ _12939_/X _18425_/Q _13003_/S vssd1 vssd1 vccd1 vccd1 _12941_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10944__S0 _10892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _12871_/A _12871_/B vssd1 vssd1 vccd1 vccd1 _12871_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__10977__S _10977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15252__A2 _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _14610_/A vssd1 vssd1 vccd1 vccd1 _18771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _19892_/Q _13290_/B _12944_/A _18689_/Q _11821_/X vssd1 vssd1 vccd1 vccd1
+ _11822_/X sky130_fd_sc_hd__a221o_1
XFILLER_27_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15590_ _15590_/A vssd1 vssd1 vccd1 vccd1 _18877_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _18752_/Q _11865_/X _14538_/X _14540_/X vssd1 vssd1 vccd1 vccd1 _18752_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11753_ _18600_/Q _11683_/X _11687_/X _18632_/Q _11752_/X vssd1 vssd1 vccd1 vccd1
+ _13257_/A sky130_fd_sc_hd__a221o_2
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10704_/A vssd1 vssd1 vccd1 vccd1 _10764_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17260_/A vssd1 vssd1 vccd1 vccd1 _19548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11684_ _11697_/A _11697_/B _11697_/C _15775_/A vssd1 vssd1 vccd1 vccd1 _11790_/B
+ sky130_fd_sc_hd__or4b_4
X_14472_ _14472_/A _14476_/C vssd1 vssd1 vccd1 vccd1 _14472_/Y sky130_fd_sc_hd__nor2_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _13406_/X _19122_/Q _16217_/S vssd1 vssd1 vccd1 vccd1 _16212_/A sky130_fd_sc_hd__mux2_1
X_10635_ _10680_/A _10634_/X _09777_/A vssd1 vssd1 vccd1 vccd1 _10635_/Y sky130_fd_sc_hd__o21ai_1
X_13423_ _17723_/A vssd1 vssd1 vccd1 vccd1 _13423_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17191_ _17191_/A vssd1 vssd1 vccd1 vccd1 _19518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09865__S1 _09851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13354_ _17710_/A vssd1 vssd1 vccd1 vccd1 _13354_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16142_ _13443_/X _19092_/Q _16144_/S vssd1 vssd1 vccd1 vccd1 _16143_/A sky130_fd_sc_hd__mux2_1
X_10566_ _19209_/Q _19800_/Q _19962_/Q _19177_/Q _10521_/X _10522_/X vssd1 vssd1 vccd1
+ vccd1 _10567_/B sky130_fd_sc_hd__mux4_1
XFILLER_128_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ _12279_/A _12279_/B _12279_/C _12301_/X vssd1 vssd1 vccd1 vccd1 _12305_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_155_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13285_ _13285_/A vssd1 vssd1 vccd1 vccd1 _18443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16073_ _19062_/Q _16072_/X _16073_/S vssd1 vssd1 vccd1 vccd1 _16074_/A sky130_fd_sc_hd__mux2_1
X_10497_ _10497_/A vssd1 vssd1 vccd1 vccd1 _10497_/X sky130_fd_sc_hd__buf_2
XANTENNA__12526__A0 _12521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15024_ _15022_/X _15023_/X _15114_/S vssd1 vssd1 vccd1 vccd1 _15024_/X sky130_fd_sc_hd__mux2_1
X_12236_ _11903_/A _12835_/B _12260_/C _18990_/Q vssd1 vssd1 vccd1 vccd1 _15254_/A
+ sky130_fd_sc_hd__a22o_1
X_19901_ _19910_/CLK _19901_/D vssd1 vssd1 vccd1 vccd1 _19901_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11424__S1 _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19832_ _20040_/CLK _19832_/D vssd1 vssd1 vccd1 vccd1 _19832_/Q sky130_fd_sc_hd__dfxtp_1
X_12167_ _12167_/A _12167_/B vssd1 vssd1 vccd1 vccd1 _12167_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__13755__C _16846_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14213__A _14239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11118_ _09791_/A _11113_/X _11115_/Y _11117_/Y _09803_/A vssd1 vssd1 vccd1 vccd1
+ _11118_/X sky130_fd_sc_hd__o221a_1
X_19763_ _19796_/CLK _19763_/D vssd1 vssd1 vccd1 vccd1 _19763_/Q sky130_fd_sc_hd__dfxtp_1
X_16975_ _16377_/X _19445_/Q _16975_/S vssd1 vssd1 vccd1 vccd1 _16976_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12098_ _12503_/A _12096_/X _12097_/X _12056_/X vssd1 vssd1 vccd1 vccd1 _12098_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11048__S _11048_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18714_ _19883_/CLK _18714_/D vssd1 vssd1 vccd1 vccd1 _18714_/Q sky130_fd_sc_hd__dfxtp_1
X_15926_ _19001_/Q _15921_/X _15925_/X vssd1 vssd1 vccd1 vccd1 _19001_/D sky130_fd_sc_hd__a21o_1
X_11049_ _19359_/Q _19694_/Q _11049_/S vssd1 vssd1 vccd1 vccd1 _11050_/B sky130_fd_sc_hd__mux2_1
X_19694_ _19726_/CLK _19694_/D vssd1 vssd1 vccd1 vccd1 _19694_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15970__C _15970_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 io_dbus_rdata[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_6
XANTENNA__10935__S0 _10703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18645_ _18653_/CLK _18645_/D vssd1 vssd1 vccd1 vccd1 _18645_/Q sky130_fd_sc_hd__dfxtp_1
X_15857_ _12082_/X _15856_/X _15843_/X input44/X vssd1 vssd1 vccd1 vccd1 _17208_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16440__A1 _13810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14808_ _14808_/A _14822_/C _14808_/C vssd1 vssd1 vccd1 vccd1 _14993_/B sky130_fd_sc_hd__and3_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12057__A2 _12046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18576_ _20005_/CLK _18576_/D vssd1 vssd1 vccd1 vccd1 _18576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15788_ _15879_/A vssd1 vssd1 vccd1 vccd1 _15788_/X sky130_fd_sc_hd__buf_2
X_17527_ _17527_/A vssd1 vssd1 vccd1 vccd1 _19669_/D sky130_fd_sc_hd__clkbuf_1
X_14739_ _14739_/A vssd1 vssd1 vccd1 vccd1 _18819_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16574__S _16580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__A _10449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09977__A _10411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17458_ _17458_/A vssd1 vssd1 vccd1 vccd1 _19636_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16409_ _19194_/Q _13765_/X _16413_/S vssd1 vssd1 vccd1 vccd1 _16410_/A sky130_fd_sc_hd__mux2_1
X_17389_ _17411_/A vssd1 vssd1 vccd1 vccd1 _17398_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10916__A _15934_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09856__S1 _09660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19128_ _19389_/CLK _19128_/D vssd1 vssd1 vccd1 vccd1 _19128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10240__A1 _09884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19059_ _19882_/CLK _19059_/D vssd1 vssd1 vccd1 vccd1 _19059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12517__A0 _15958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11415__S1 _11208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12850__B _12850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09714_ _10294_/A vssd1 vssd1 vccd1 vccd1 _09946_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09645_ _09568_/X _09616_/Y _09634_/Y _09641_/Y _09644_/Y vssd1 vssd1 vccd1 vccd1
+ _09645_/X sky130_fd_sc_hd__o32a_1
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09576_ _10670_/A vssd1 vssd1 vccd1 vccd1 _10549_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09449__B1 _09279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16484__S _16486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18265__A _18265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10154__S1 _10153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11103__S0 _11293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13202__A _17681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ _09547_/A _10409_/Y _10418_/X _10078_/X _10419_/Y vssd1 vssd1 vccd1 vccd1
+ _15960_/B sky130_fd_sc_hd__o32a_2
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10351_ _10351_/A _12854_/B vssd1 vssd1 vccd1 vccd1 _10352_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10037__S _10037_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18204__S _18206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ _13070_/A vssd1 vssd1 vccd1 vccd1 _13070_/X sky130_fd_sc_hd__clkbuf_2
X_10282_ _10294_/A _10276_/X _10278_/Y _10281_/Y vssd1 vssd1 vccd1 vccd1 _10282_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12021_ _12016_/X _12168_/S _12020_/X vssd1 vssd1 vccd1 vccd1 _12021_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_3_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16659__S _16663_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14968__A _15553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16760_ _19350_/Q _13854_/X _16762_/S vssd1 vssd1 vccd1 vccd1 _16761_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13484__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13972_ _18564_/Q _13973_/C _18565_/Q vssd1 vssd1 vccd1 vccd1 _13974_/B sky130_fd_sc_hd__a21oi_1
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15711_ _09481_/B _15705_/X _15710_/X _14540_/X vssd1 vssd1 vccd1 vccd1 _18931_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10298__B2 _09823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ _13502_/S vssd1 vssd1 vccd1 vccd1 _13003_/S sky130_fd_sc_hd__buf_4
X_16691_ _16691_/A _16691_/B _16298_/C vssd1 vssd1 vccd1 vccd1 _17882_/B sky130_fd_sc_hd__or3b_2
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16422__A1 _13784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15225__A2 _09433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10393__S1 _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18430_ _19567_/CLK _18430_/D vssd1 vssd1 vccd1 vccd1 _18430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15642_ _18900_/Q _18521_/Q _15644_/S vssd1 vssd1 vccd1 vccd1 _15643_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13236__A1 _13223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12854_ _12857_/A _12854_/B vssd1 vssd1 vccd1 vccd1 _12854_/Y sky130_fd_sc_hd__nor2_2
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _15762_/A vssd1 vssd1 vccd1 vccd1 _15783_/B sky130_fd_sc_hd__clkbuf_1
X_18361_ _17646_/X _20012_/Q _18363_/S vssd1 vssd1 vccd1 vccd1 _18362_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16394__S _16394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output100_A _12186_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15573_ _15573_/A vssd1 vssd1 vccd1 vccd1 _18869_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _12785_/A vssd1 vssd1 vccd1 vccd1 _12789_/A sky130_fd_sc_hd__clkinv_2
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13811__S _13820_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17312_ _17312_/A vssd1 vssd1 vccd1 vccd1 _19571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09797__A _10382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14524_ _14526_/B _14526_/C _14507_/X vssd1 vssd1 vccd1 vccd1 _14524_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18292_ _18292_/A vssd1 vssd1 vccd1 vccd1 _19981_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11736_ _18663_/Q _11815_/A _11855_/B _18731_/Q vssd1 vssd1 vccd1 vccd1 _11736_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17243_ _17144_/X _19541_/Q _17243_/S vssd1 vssd1 vccd1 vccd1 _17244_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14736__A1 _13727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14455_ _18717_/Q _14452_/B _14454_/Y vssd1 vssd1 vccd1 vccd1 _18717_/D sky130_fd_sc_hd__o21a_1
X_11667_ _11667_/A _14805_/A _11667_/C vssd1 vssd1 vccd1 vccd1 _11975_/D sky130_fd_sc_hd__and3_1
X_13406_ _17720_/A vssd1 vssd1 vccd1 vccd1 _13406_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17174_ _17173_/X _19513_/Q _17177_/S vssd1 vssd1 vccd1 vccd1 _17175_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10618_ _10618_/A vssd1 vssd1 vccd1 vccd1 _11186_/S sky130_fd_sc_hd__clkbuf_4
X_11598_ _11598_/A vssd1 vssd1 vccd1 vccd1 _11599_/B sky130_fd_sc_hd__inv_2
X_14386_ _14386_/A vssd1 vssd1 vccd1 vccd1 _18691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16489__A1 _13774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16125_ _13302_/X _19084_/Q _16133_/S vssd1 vssd1 vccd1 vccd1 _16126_/A sky130_fd_sc_hd__mux2_1
X_10549_ _10549_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10549_/X sky130_fd_sc_hd__or2_1
X_13337_ _14510_/B _11776_/X _13333_/X _13336_/X vssd1 vssd1 vccd1 vccd1 _13683_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_109_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16056_ _16056_/A vssd1 vssd1 vccd1 vccd1 _19056_/D sky130_fd_sc_hd__clkbuf_1
X_13268_ _13268_/A _13268_/B _13288_/B vssd1 vssd1 vccd1 vccd1 _13268_/X sky130_fd_sc_hd__or3_1
XFILLER_124_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13172__A0 _18846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__A1 _09884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15007_ _15048_/A _15007_/B vssd1 vssd1 vccd1 vccd1 _15405_/A sky130_fd_sc_hd__nor2_1
XFILLER_124_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12219_ _12150_/A _12215_/X _12216_/X _12218_/Y vssd1 vssd1 vccd1 vccd1 _12220_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13199_ input6/X _13091_/A _13094_/A vssd1 vssd1 vccd1 vccd1 _13199_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11183__C1 _09817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19815_ _19816_/CLK _19815_/D vssd1 vssd1 vccd1 vccd1 _19815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16569__S _16569_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16958_ _16352_/X _19437_/Q _16964_/S vssd1 vssd1 vccd1 vccd1 _16959_/A sky130_fd_sc_hd__mux2_1
X_19746_ _20036_/CLK _19746_/D vssd1 vssd1 vccd1 vccd1 _19746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15909_ _15909_/A vssd1 vssd1 vccd1 vccd1 _18996_/D sky130_fd_sc_hd__clkbuf_1
X_19677_ _19935_/CLK _19677_/D vssd1 vssd1 vccd1 vccd1 _19677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16889_ _16889_/A vssd1 vssd1 vccd1 vccd1 _19406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09430_ _13926_/A _15719_/A vssd1 vssd1 vccd1 vccd1 _15624_/A sky130_fd_sc_hd__nor2_8
X_18628_ _18660_/CLK _18628_/D vssd1 vssd1 vccd1 vccd1 _18628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09361_ _18753_/Q _18748_/Q _18749_/Q _18754_/Q vssd1 vssd1 vccd1 vccd1 _09361_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14975__A1 _12871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18559_ _18741_/CLK _18559_/D vssd1 vssd1 vccd1 vccd1 _18559_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11333__S0 _11409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_143_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09292_ _09292_/A _09292_/B _09292_/C _14819_/A vssd1 vssd1 vccd1 vccd1 _09292_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_21_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17913__A1 _17036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14727__A1 _11898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13022__A _17010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13957__A _13991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12861__A _12861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16333__A _16400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18024__S _18024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput130 _12863_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[29] sky130_fd_sc_hd__buf_2
XFILLER_133_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput141 _11908_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wr_en sky130_fd_sc_hd__buf_2
XANTENNA__17863__S _17865_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput152 _12534_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[19] sky130_fd_sc_hd__buf_2
XFILLER_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput163 _12776_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[29] sky130_fd_sc_hd__buf_2
XFILLER_115_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10072__S0 _09918_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_68_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17164__A _17180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09628_ _10462_/A vssd1 vssd1 vccd1 vccd1 _10369_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09559_ _09559_/A vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _12571_/A _14863_/A vssd1 vssd1 vccd1 vccd1 _12572_/A sky130_fd_sc_hd__nand2_1
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12441__A2 _12389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09410__A _09410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11521_ _15966_/C _12855_/B vssd1 vssd1 vccd1 vccd1 _11522_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16942__S _16942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14028__A _14044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14240_ _18648_/Q _14236_/A _14239_/Y vssd1 vssd1 vccd1 vccd1 _18648_/D sky130_fd_sc_hd__o21a_1
X_11452_ _11452_/A _12825_/B vssd1 vssd1 vccd1 vccd1 _11611_/A sky130_fd_sc_hd__nor2_1
XFILLER_172_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14194__A2 _14197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15391__A1 _18850_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10403_ _19675_/Q _19441_/Q _18506_/Q _19771_/Q _10319_/X _10320_/X vssd1 vssd1 vccd1
+ vccd1 _10403_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10204__A1 _09849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10204__B2 _18859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13867__A _15807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14171_ _18628_/Q _14172_/C _18629_/Q vssd1 vssd1 vccd1 vccd1 _14173_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__17339__A _17339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11383_ _11414_/A _11382_/X _09681_/A vssd1 vssd1 vccd1 vccd1 _11383_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11952__A1 _09522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _19342_/Q _19613_/Q _19837_/Q _19581_/Q _10152_/X _10153_/X vssd1 vssd1 vccd1
+ vccd1 _10335_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16340__A0 _16339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input61_A io_ibus_inst[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ _19891_/Q _13451_/B vssd1 vssd1 vccd1 vccd1 _13122_/X sky130_fd_sc_hd__and2_1
XFILLER_140_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17930_ _17930_/A vssd1 vssd1 vccd1 vccd1 _19835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13053_ _13053_/A _13053_/B vssd1 vssd1 vccd1 vccd1 _13053_/X sky130_fd_sc_hd__or2_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _19936_/Q _19550_/Q _20000_/Q _19119_/Q _09657_/A _10261_/X vssd1 vssd1 vccd1
+ vccd1 _10266_/B sky130_fd_sc_hd__mux4_1
XFILLER_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11165__C1 _11095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ _12004_/A _12004_/B _12004_/C _12004_/D vssd1 vssd1 vccd1 vccd1 _15633_/D
+ sky130_fd_sc_hd__or4_2
X_17861_ _19805_/Q _17065_/X _17865_/S vssd1 vssd1 vccd1 vccd1 _17862_/A sky130_fd_sc_hd__mux2_1
X_10196_ _10200_/A _10196_/B vssd1 vssd1 vccd1 vccd1 _10196_/X sky130_fd_sc_hd__or2_1
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output148_A _12427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16812_ _16812_/A vssd1 vssd1 vccd1 vccd1 _19372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17074__A _17074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19600_ _19957_/CLK _19600_/D vssd1 vssd1 vccd1 vccd1 _19600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17792_ _17792_/A vssd1 vssd1 vccd1 vccd1 _19774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19531_ _19981_/CLK _19531_/D vssd1 vssd1 vccd1 vccd1 _19531_/Q sky130_fd_sc_hd__dfxtp_1
X_16743_ _19342_/Q _13829_/X _16747_/S vssd1 vssd1 vccd1 vccd1 _16744_/A sky130_fd_sc_hd__mux2_1
X_13955_ _13956_/B _13956_/C _18559_/Q vssd1 vssd1 vccd1 vccd1 _13957_/B sky130_fd_sc_hd__a21oi_1
XFILLER_59_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10366__S1 _10054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19462_ _19856_/CLK _19462_/D vssd1 vssd1 vccd1 vccd1 _19462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12906_ _12906_/A vssd1 vssd1 vccd1 vccd1 _12906_/X sky130_fd_sc_hd__clkbuf_4
X_16674_ _16377_/X _19312_/Q _16674_/S vssd1 vssd1 vccd1 vccd1 _16675_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _12340_/B _13883_/X _12346_/Y _12351_/X _13885_/X vssd1 vssd1 vccd1 vccd1
+ _18530_/D sky130_fd_sc_hd__o221a_1
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18413_ _18413_/A vssd1 vssd1 vccd1 vccd1 _20035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15625_ _18893_/Q _18925_/Q _15901_/S vssd1 vssd1 vccd1 vccd1 _15626_/A sky130_fd_sc_hd__mux2_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12833_/A _12837_/B vssd1 vssd1 vccd1 vccd1 _12838_/A sky130_fd_sc_hd__and2b_4
X_19393_ _19981_/CLK _19393_/D vssd1 vssd1 vccd1 vccd1 _19393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18344_ _17726_/X _20005_/Q _18346_/S vssd1 vssd1 vccd1 vccd1 _18345_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _15552_/Y _15181_/A _14970_/B vssd1 vssd1 vccd1 vccd1 _15556_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _18546_/Q _18547_/Q _12768_/C vssd1 vssd1 vccd1 vccd1 _12793_/B sky130_fd_sc_hd__and3_1
XANTENNA__12665__B _15487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17948__S _17948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__A _18939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14507_ _14507_/A vssd1 vssd1 vccd1 vccd1 _14507_/X sky130_fd_sc_hd__buf_4
XFILLER_159_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18275_ _18275_/A vssd1 vssd1 vccd1 vccd1 _19974_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11719_ _13747_/A vssd1 vssd1 vccd1 vccd1 _14552_/A sky130_fd_sc_hd__buf_2
X_15487_ _15487_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _15487_/Y sky130_fd_sc_hd__nor2_1
X_12699_ _12338_/A _12697_/X _12698_/Y vssd1 vssd1 vccd1 vccd1 _12699_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17226_ _17119_/X _19533_/Q _17232_/S vssd1 vssd1 vccd1 vccd1 _17227_/A sky130_fd_sc_hd__mux2_1
Xinput10 io_dbus_rdata[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_4
X_14438_ _18706_/Q _14439_/C _18707_/Q vssd1 vssd1 vccd1 vccd1 _14440_/B sky130_fd_sc_hd__a21oi_1
Xinput21 io_dbus_rdata[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_2
XANTENNA__15976__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput32 io_dbus_rdata[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_2
Xinput43 io_ibus_inst[18] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
Xinput54 io_ibus_inst[28] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_8
X_17157_ _17694_/A vssd1 vssd1 vccd1 vccd1 _17157_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput65 io_ibus_inst[9] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_6
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14369_ _18677_/Q _14369_/B _14373_/D vssd1 vssd1 vccd1 vccd1 _14371_/C sky130_fd_sc_hd__and3_1
XFILLER_116_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16153__A _16221_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16108_ _16108_/A vssd1 vssd1 vccd1 vccd1 _19076_/D sky130_fd_sc_hd__clkbuf_1
X_17088_ _19482_/Q _17087_/X _17088_/S vssd1 vssd1 vccd1 vccd1 _17089_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16039_ _16039_/A vssd1 vssd1 vccd1 vccd1 _19048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18084__A0 _18849_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10903__C1 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19729_ _19731_/CLK _19729_/D vssd1 vssd1 vccd1 vccd1 _19729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11236__S _11295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _18957_/Q vssd1 vssd1 vccd1 vccd1 _15777_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14948__A1 _15219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12856__A _12857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09344_ _09442_/A _09442_/B vssd1 vssd1 vccd1 vccd1 _09345_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09275_ _09275_/A _11948_/B _09275_/C _09274_/X vssd1 vssd1 vccd1 vccd1 _09292_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_138_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16762__S _16762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10293__S0 _10037_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16998__A _16998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17593__S _17595_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13687__A1 _18476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _10050_/A vssd1 vssd1 vccd1 vccd1 _10587_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09405__A _09405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13740_ _14560_/A _19024_/Q vssd1 vssd1 vccd1 vccd1 _13740_/Y sky130_fd_sc_hd__nand2_1
X_10952_ _10952_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _10952_/X sky130_fd_sc_hd__or2_1
XFILLER_71_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13671_ _13671_/A vssd1 vssd1 vccd1 vccd1 _18474_/D sky130_fd_sc_hd__clkbuf_1
X_10883_ _18434_/Q _19463_/Q _19500_/Q _19074_/Q _10919_/S _10596_/A vssd1 vssd1 vccd1
+ vccd1 _10883_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16238__A _16295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15410_ _15410_/A _15410_/B vssd1 vssd1 vccd1 vccd1 _15410_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12622_ _12601_/A _12623_/C _18541_/Q vssd1 vssd1 vccd1 vccd1 _12624_/A sky130_fd_sc_hd__a21oi_1
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16390_ _17726_/A vssd1 vssd1 vccd1 vccd1 _16390_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15341_ _15282_/X _15332_/X _15340_/X _15324_/X vssd1 vssd1 vccd1 vccd1 _15341_/X
+ sky130_fd_sc_hd__a211o_1
X_12553_ _12790_/A vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16672__S _16674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14981__A _15016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11504_ _10858_/A _11503_/X _09793_/A vssd1 vssd1 vccd1 vccd1 _11504_/Y sky130_fd_sc_hd__o21ai_1
X_18060_ _18842_/Q _13579_/X _18067_/S vssd1 vssd1 vccd1 vccd1 _18060_/X sky130_fd_sc_hd__mux2_1
X_15272_ _15323_/A _15272_/B _15272_/C vssd1 vssd1 vccd1 vccd1 _15272_/X sky130_fd_sc_hd__and3_1
XFILLER_157_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12484_ _12422_/X _12482_/Y _12532_/C _12425_/X vssd1 vssd1 vccd1 vccd1 _12484_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_8_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13375__B1 _11843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17011_ _17094_/S vssd1 vssd1 vccd1 vccd1 _17024_/S sky130_fd_sc_hd__buf_2
XFILLER_138_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14223_ _18960_/Q _18959_/Q _18940_/Q _16474_/B vssd1 vssd1 vccd1 vccd1 _14226_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11435_ _11435_/A _11435_/B vssd1 vssd1 vccd1 vccd1 _11435_/X sky130_fd_sc_hd__or2_1
XFILLER_172_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11366_ _11414_/A _11366_/B vssd1 vssd1 vccd1 vccd1 _11366_/Y sky130_fd_sc_hd__nor2_1
X_14154_ _14189_/A _14154_/B _14154_/C vssd1 vssd1 vccd1 vccd1 _18623_/D sky130_fd_sc_hd__nor3_1
XFILLER_152_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13127__B1 _13082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10317_ _19150_/Q _19411_/Q _19310_/Q _19645_/Q _10354_/S _10185_/X vssd1 vssd1 vccd1
+ vccd1 _10317_/X sky130_fd_sc_hd__mux4_1
X_13105_ _18655_/Q _13081_/A _11824_/A _18623_/Q vssd1 vssd1 vccd1 vccd1 _13105_/X
+ sky130_fd_sc_hd__a22o_1
X_14085_ _14086_/B _14086_/C _14084_/Y vssd1 vssd1 vccd1 vccd1 _18604_/D sky130_fd_sc_hd__o21a_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18962_ _18992_/CLK _18962_/D vssd1 vssd1 vccd1 vccd1 _18962_/Q sky130_fd_sc_hd__dfxtp_1
X_11297_ _19658_/Q _19424_/Q _18489_/Q _19754_/Q _11155_/A _11172_/A vssd1 vssd1 vccd1
+ vccd1 _11297_/X sky130_fd_sc_hd__mux4_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12006__A _18520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ _19828_/Q _17036_/X _17915_/S vssd1 vssd1 vccd1 vccd1 _17914_/A sky130_fd_sc_hd__mux2_1
X_10248_ _10248_/A _10047_/Y vssd1 vssd1 vccd1 vccd1 _10248_/X sky130_fd_sc_hd__or2b_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _19488_/Q vssd1 vssd1 vccd1 vccd1 _13349_/S sky130_fd_sc_hd__clkbuf_2
X_18893_ _18926_/CLK _18893_/D vssd1 vssd1 vccd1 vccd1 _18893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11845__A _13290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17008__S _17008_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17844_ _17844_/A vssd1 vssd1 vccd1 vccd1 _19797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15317__A _15393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10179_ _10246_/A _10179_/B vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17775_ _17775_/A vssd1 vssd1 vccd1 vccd1 _19766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14987_ _14978_/X _14985_/X _14986_/X vssd1 vssd1 vccd1 vccd1 _15546_/B sky130_fd_sc_hd__o21a_1
XFILLER_93_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10339__S1 _10223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16726_ _16726_/A vssd1 vssd1 vccd1 vccd1 _19334_/D sky130_fd_sc_hd__clkbuf_1
X_19514_ _20035_/CLK _19514_/D vssd1 vssd1 vccd1 vccd1 _19514_/Q sky130_fd_sc_hd__dfxtp_1
X_13938_ _18554_/Q _18553_/Q _18552_/Q _13938_/D vssd1 vssd1 vccd1 vccd1 _13947_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_75_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19445_ _19839_/CLK _19445_/D vssd1 vssd1 vccd1 vccd1 _19445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16657_ _16352_/X _19304_/Q _16663_/S vssd1 vssd1 vccd1 vccd1 _16658_/A sky130_fd_sc_hd__mux2_1
X_13869_ _13879_/A vssd1 vssd1 vccd1 vccd1 _14529_/A sky130_fd_sc_hd__buf_6
XFILLER_23_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15608_ _15608_/A vssd1 vssd1 vccd1 vccd1 _18885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19376_ _20035_/CLK _19376_/D vssd1 vssd1 vccd1 vccd1 _19376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16588_ _16588_/A vssd1 vssd1 vccd1 vccd1 _19273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12405__A2 _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_16_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18327_ _17700_/X _19997_/Q _18335_/S vssd1 vssd1 vccd1 vccd1 _18328_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11613__B1 _11462_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15539_ _15539_/A _15542_/A vssd1 vssd1 vccd1 vccd1 _15539_/X sky130_fd_sc_hd__or2_1
XANTENNA__10196__A _10200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _18258_/A vssd1 vssd1 vccd1 vccd1 _19966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ _17209_/A vssd1 vssd1 vccd1 vccd1 _19526_/D sky130_fd_sc_hd__clkbuf_1
X_18189_ _17710_/X _19936_/Q _18191_/S vssd1 vssd1 vccd1 vccd1 _18190_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ _09884_/X _09949_/X _09960_/X _09913_/X _09961_/Y vssd1 vssd1 vccd1 vccd1
+ _12862_/B sky130_fd_sc_hd__o32a_4
XANTENNA__18302__S _18302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13669__A1 _13667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18057__A0 _18841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09968__S0 _09967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ _09750_/A _09892_/X _09809_/X vssd1 vssd1 vccd1 vccd1 _09893_/Y sky130_fd_sc_hd__o21ai_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10578__S1 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13181__S _13203_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15594__A1 _18911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09327_ _18985_/Q _12004_/A vssd1 vssd1 vccd1 vccd1 _09699_/A sky130_fd_sc_hd__or2_1
XFILLER_166_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09895__A _09895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ _09311_/A vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_166_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09189_ _09189_/A vssd1 vssd1 vccd1 vccd1 _12003_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11220_ _11287_/A _11219_/X _11058_/X vssd1 vssd1 vccd1 vccd1 _11220_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_153_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16224__C _16298_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11151_ _11088_/A _11150_/X _11095_/X vssd1 vssd1 vccd1 vccd1 _11151_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_161_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14740__S _14742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10102_ _09809_/A _10093_/Y _10097_/Y _10101_/Y _09807_/X vssd1 vssd1 vccd1 vccd1
+ _10102_/X sky130_fd_sc_hd__o311a_1
XANTENNA__09834__S _09898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13864__B _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ _09848_/A _11060_/X _11081_/Y _09537_/A _18840_/Q vssd1 vssd1 vccd1 vccd1
+ _15925_/C sky130_fd_sc_hd__a32o_4
X_10033_ _10007_/Y _10015_/Y _10030_/Y _10032_/Y _09823_/A vssd1 vssd1 vccd1 vccd1
+ _10033_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14910_ _15177_/B _12664_/A _14915_/S vssd1 vssd1 vccd1 vccd1 _14910_/X sky130_fd_sc_hd__mux2_1
X_15890_ _14750_/B _15875_/X _15879_/X input55/X vssd1 vssd1 vccd1 vccd1 _15891_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input24_A io_dbus_rdata[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ _14990_/C _14846_/B vssd1 vssd1 vccd1 vccd1 _15444_/A sky130_fd_sc_hd__or2_1
XFILLER_64_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13880__A _15833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17560_ _19686_/Q vssd1 vssd1 vccd1 vccd1 _17561_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14772_ _11660_/A _09279_/X _15747_/A _14778_/A _13531_/A vssd1 vssd1 vccd1 vccd1
+ _14773_/B sky130_fd_sc_hd__a32o_1
XFILLER_63_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11984_ _18970_/Q _11983_/X _12084_/S vssd1 vssd1 vccd1 vccd1 _11984_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16511_ _19239_/Q _13806_/X _16519_/S vssd1 vssd1 vccd1 vccd1 _16512_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13723_ _18893_/Q _13723_/B vssd1 vssd1 vccd1 vccd1 _13723_/Y sky130_fd_sc_hd__nand2_1
X_10935_ _19922_/Q _19536_/Q _19986_/Q _19105_/Q _10703_/A _10663_/A vssd1 vssd1 vccd1
+ vccd1 _10936_/B sky130_fd_sc_hd__mux4_1
X_17491_ _17491_/A vssd1 vssd1 vccd1 vccd1 _19651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19230_ _19726_/CLK _19230_/D vssd1 vssd1 vccd1 vccd1 _19230_/Q sky130_fd_sc_hd__dfxtp_1
X_16442_ _19209_/Q _13813_/X _16446_/S vssd1 vssd1 vccd1 vccd1 _16443_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13654_ _18884_/Q _13654_/B vssd1 vssd1 vccd1 vccd1 _13654_/Y sky130_fd_sc_hd__nand2_1
X_10866_ _10843_/A _10863_/X _10865_/X _09793_/A vssd1 vssd1 vccd1 vccd1 _10866_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13596__A0 _13591_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19161_ _19720_/CLK _19161_/D vssd1 vssd1 vccd1 vccd1 _19161_/Q sky130_fd_sc_hd__dfxtp_1
X_12605_ _18779_/Q _12628_/C vssd1 vssd1 vccd1 vccd1 _12605_/Y sky130_fd_sc_hd__nor2_1
X_16373_ _16373_/A vssd1 vssd1 vccd1 vccd1 _19182_/D sky130_fd_sc_hd__clkbuf_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _18463_/Q _13583_/X _13617_/S vssd1 vssd1 vccd1 vccd1 _13586_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10797_ _10953_/S vssd1 vssd1 vccd1 vccd1 _10797_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_157_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18112_ _18111_/X _19905_/Q _18112_/S vssd1 vssd1 vccd1 vccd1 _18113_/A sky130_fd_sc_hd__mux2_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15324_ _15400_/A vssd1 vssd1 vccd1 vccd1 _15324_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19092_ _19587_/CLK _19092_/D vssd1 vssd1 vccd1 vccd1 _19092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12536_ _12536_/A _12536_/B vssd1 vssd1 vccd1 vccd1 _12539_/B sky130_fd_sc_hd__nor2_1
XFILLER_129_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18043_ _18837_/Q hold7/A _18050_/S vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__mux2_1
XANTENNA__14545__C1 _14540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15255_ _15218_/X _15250_/Y _15254_/Y vssd1 vssd1 vccd1 vccd1 _15256_/C sky130_fd_sc_hd__a21oi_1
X_12467_ _12467_/A vssd1 vssd1 vccd1 vccd1 _15373_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14216__A _14239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13899__A1 _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output92_A _12766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ _18640_/Q _14207_/C _18641_/Q vssd1 vssd1 vccd1 vccd1 _14208_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11418_ _11131_/A _11415_/X _11417_/X vssd1 vssd1 vccd1 vccd1 _11418_/Y sky130_fd_sc_hd__o21ai_1
X_15186_ _15489_/A _15491_/B vssd1 vssd1 vccd1 vccd1 _15186_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12398_ _18771_/Q vssd1 vssd1 vccd1 vccd1 _12399_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14137_ _14146_/A _14142_/C vssd1 vssd1 vccd1 vccd1 _14137_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11349_ _19226_/Q _19721_/Q _11441_/S vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__mux2_1
X_19994_ _19994_/CLK _19994_/D vssd1 vssd1 vccd1 vccd1 _19994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14068_ _14070_/B _14070_/C _14059_/X vssd1 vssd1 vccd1 vccd1 _14068_/Y sky130_fd_sc_hd__a21oi_1
X_18945_ _18974_/CLK _18945_/D vssd1 vssd1 vccd1 vccd1 _18945_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16150__B _16150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17961__S _17965_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13019_ _13359_/B _13019_/B vssd1 vssd1 vccd1 vccd1 _13019_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18876_ _18878_/CLK _18876_/D vssd1 vssd1 vccd1 vccd1 _18876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17827_ _17827_/A vssd1 vssd1 vccd1 vccd1 _19789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13790__A _17026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15812__A2 _11860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17758_ _17662_/X _19759_/Q _17760_/S vssd1 vssd1 vccd1 vccd1 _17759_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16709_ _16709_/A vssd1 vssd1 vccd1 vccd1 _19326_/D sky130_fd_sc_hd__clkbuf_1
X_17689_ _17688_/X _19735_/Q _17698_/S vssd1 vssd1 vccd1 vccd1 _17690_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19428_ _19758_/CLK _19428_/D vssd1 vssd1 vccd1 vccd1 _19428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19359_ _19758_/CLK _19359_/D vssd1 vssd1 vccd1 vccd1 _19359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15328__A1 _18846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12853__B _12853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__A _10654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15790__A1_N _15785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_13_0_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19379_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10799__S1 _10625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13965__A _13991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18032__S _18044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09945_ _19941_/Q _19555_/Q _20005_/Q _19124_/Q _09950_/S _09940_/X vssd1 vssd1 vccd1
+ vccd1 _09946_/B sky130_fd_sc_hd__mux4_1
XFILLER_98_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09876_ _09876_/A vssd1 vssd1 vccd1 vccd1 _09876_/X sky130_fd_sc_hd__buf_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10720_ _11477_/A _10718_/X _10719_/X vssd1 vssd1 vccd1 vccd1 _10720_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09402__B _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_191_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _10652_/A _12847_/B vssd1 vssd1 vccd1 vccd1 _10653_/A sky130_fd_sc_hd__and2_1
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10582_ _09796_/A _10572_/Y _10576_/Y _10581_/Y _09806_/A vssd1 vssd1 vccd1 vccd1
+ _10582_/X sky130_fd_sc_hd__o311a_1
XANTENNA__12250__B1 _12246_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13370_ _18890_/Q vssd1 vssd1 vccd1 vccd1 _13699_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12321_ _12406_/A vssd1 vssd1 vccd1 vccd1 _15306_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14036__A _14044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ _14966_/A _14957_/S _14832_/A vssd1 vssd1 vccd1 vccd1 _15040_/Y sky130_fd_sc_hd__a21boi_1
X_12252_ _18463_/Q _12372_/B vssd1 vssd1 vccd1 vccd1 _12252_/X sky130_fd_sc_hd__or2_1
XFILLER_135_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11203_ _11283_/A _11197_/X _11199_/X _11202_/X vssd1 vssd1 vccd1 vccd1 _11203_/X
+ sky130_fd_sc_hd__o22a_1
X_12183_ _12183_/A _14909_/A vssd1 vssd1 vccd1 vccd1 _12185_/A sky130_fd_sc_hd__or2b_1
XFILLER_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11134_ _19919_/Q _19533_/Q _19983_/Q _19102_/Q _10995_/X _10996_/X vssd1 vssd1 vccd1
+ vccd1 _11135_/B sky130_fd_sc_hd__mux4_1
X_16991_ _16991_/A vssd1 vssd1 vccd1 vccd1 _19452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15942_ _15942_/A vssd1 vssd1 vccd1 vccd1 _15964_/A sky130_fd_sc_hd__buf_2
X_11065_ _11073_/A vssd1 vssd1 vccd1 vccd1 _11065_/X sky130_fd_sc_hd__clkbuf_4
X_18730_ _18731_/CLK _18730_/D vssd1 vssd1 vccd1 vccd1 _18730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10016_ _10172_/A vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__buf_2
XANTENNA__10867__A1 _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18661_ _18731_/CLK _18661_/D vssd1 vssd1 vccd1 vccd1 _18661_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output130_A _12863_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15873_ _15881_/A _16844_/B vssd1 vssd1 vccd1 vccd1 _15874_/A sky130_fd_sc_hd__and2_1
XANTENNA__16397__S _16400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13814__S _13820_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17612_ _17612_/A vssd1 vssd1 vccd1 vccd1 _19708_/D sky130_fd_sc_hd__clkbuf_1
X_14824_ _14973_/A _14973_/B vssd1 vssd1 vccd1 vccd1 _15048_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18592_ _18724_/CLK _18592_/D vssd1 vssd1 vccd1 vccd1 _18592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17543_ _17543_/A vssd1 vssd1 vccd1 vccd1 _19677_/D sky130_fd_sc_hd__clkbuf_1
X_14755_ _14755_/A _14761_/C vssd1 vssd1 vccd1 vccd1 _14764_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11967_ _11967_/A vssd1 vssd1 vccd1 vccd1 _11967_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10714__S1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11292__A1 _18836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13706_ _18479_/Q _13526_/A _13701_/Y _13705_/X vssd1 vssd1 vccd1 vccd1 _18479_/D
+ sky130_fd_sc_hd__o22a_1
X_17474_ _17474_/A vssd1 vssd1 vccd1 vccd1 _19643_/D sky130_fd_sc_hd__clkbuf_1
X_10918_ _10918_/A _10918_/B vssd1 vssd1 vccd1 vccd1 _11605_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_1_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19979_/CLK sky130_fd_sc_hd__clkbuf_16
X_14686_ _18795_/Q _13546_/X _14694_/S vssd1 vssd1 vccd1 vccd1 _14687_/A sky130_fd_sc_hd__mux2_1
X_11898_ _11731_/X _11896_/X _11897_/Y _11723_/X _19018_/Q vssd1 vssd1 vccd1 vccd1
+ _11898_/X sky130_fd_sc_hd__a32o_4
X_19213_ _19836_/CLK _19213_/D vssd1 vssd1 vccd1 vccd1 _19213_/Q sky130_fd_sc_hd__dfxtp_1
X_16425_ _16425_/A vssd1 vssd1 vccd1 vccd1 _19201_/D sky130_fd_sc_hd__clkbuf_1
X_13637_ _18881_/Q _13637_/B vssd1 vssd1 vccd1 vccd1 _13638_/B sky130_fd_sc_hd__nand2_1
XFILLER_158_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10849_ _10858_/A _10846_/X _10848_/X _09794_/A vssd1 vssd1 vccd1 vccd1 _10849_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13033__A2 _12889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16426__A _16472_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17021__S _17024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19144_ _20025_/CLK _19144_/D vssd1 vssd1 vccd1 vccd1 _19144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16356_ _16355_/X _19177_/Q _16362_/S vssd1 vssd1 vccd1 vccd1 _16357_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13568_ _18461_/Q _13567_/X _13575_/S vssd1 vssd1 vccd1 vccd1 _13569_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15307_ _15305_/X _15301_/Y _15306_/Y vssd1 vssd1 vccd1 vccd1 _15308_/C sky130_fd_sc_hd__a21oi_1
X_19075_ _19637_/CLK _19075_/D vssd1 vssd1 vccd1 vccd1 _19075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12519_ _12519_/A vssd1 vssd1 vccd1 vccd1 _15397_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16287_ _13423_/X _19155_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _16288_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13499_ _12874_/X _13484_/Y _13498_/X vssd1 vssd1 vccd1 vccd1 _17093_/A sky130_fd_sc_hd__o21ai_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18026_ _18053_/A vssd1 vssd1 vccd1 vccd1 _18050_/S sky130_fd_sc_hd__clkbuf_2
X_15238_ _15400_/A vssd1 vssd1 vccd1 vccd1 _15238_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15984__B _16846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14533__A2 _13650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15169_ _15169_/A vssd1 vssd1 vccd1 vccd1 _15298_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10555__B1 _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19977_ _19978_/CLK _19977_/D vssd1 vssd1 vccd1 vccd1 _19977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09730_ _10166_/S vssd1 vssd1 vccd1 vccd1 _10277_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18928_ _18928_/CLK _18928_/D vssd1 vssd1 vccd1 vccd1 _18928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09661_ _10972_/A vssd1 vssd1 vccd1 vccd1 _11199_/A sky130_fd_sc_hd__clkinv_2
XFILLER_83_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18859_ _19010_/CLK _18859_/D vssd1 vssd1 vccd1 vccd1 _18859_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09592_ _10586_/S vssd1 vssd1 vccd1 vccd1 _10493_/S sky130_fd_sc_hd__buf_2
XANTENNA__16100__S _16100_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12848__B _12848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13272__A2 _13269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12864__A _12866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14772__A2 _09279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09936__C1 _09876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_138_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09928_ _19941_/Q _19555_/Q _20005_/Q _19124_/Q _09659_/S _09647_/A vssd1 vssd1 vccd1
+ vccd1 _09929_/B sky130_fd_sc_hd__mux4_1
XFILLER_131_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11197__S1 _11077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10849__A1 _10858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _19157_/Q _19418_/Q _19317_/Q _19652_/Q _09855_/A _09642_/A vssd1 vssd1 vccd1
+ vccd1 _09860_/B sky130_fd_sc_hd__mux4_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _14957_/S _12870_/B vssd1 vssd1 vccd1 vccd1 _12871_/B sky130_fd_sc_hd__nor2_4
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _18465_/Q _11870_/A _11671_/A _18712_/Q vssd1 vssd1 vccd1 vccd1 _11821_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16945__S _16953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _17208_/A vssd1 vssd1 vccd1 vccd1 _14540_/X sky130_fd_sc_hd__buf_2
XANTENNA__11274__A1 _11258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _18664_/Q _13081_/A _12890_/A _18732_/Q vssd1 vssd1 vccd1 vccd1 _11752_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10703_/A vssd1 vssd1 vccd1 vccd1 _10704_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14471_ _14471_/A vssd1 vssd1 vccd1 vccd1 _14476_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11683_ _13057_/A vssd1 vssd1 vccd1 vccd1 _11683_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16210_/A vssd1 vssd1 vccd1 vccd1 _19121_/D sky130_fd_sc_hd__clkbuf_1
X_13422_ _17081_/A vssd1 vssd1 vccd1 vccd1 _17723_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10634_ _18440_/Q _19469_/Q _19506_/Q _19080_/Q _09726_/A _10626_/X vssd1 vssd1 vccd1
+ vccd1 _10634_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17190_ _17189_/X _19518_/Q _17193_/S vssd1 vssd1 vccd1 vccd1 _17191_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17776__S _17782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16141_ _16141_/A vssd1 vssd1 vccd1 vccd1 _19091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13353_ _17068_/A vssd1 vssd1 vccd1 vccd1 _17710_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10565_ _10567_/A _10564_/X _09777_/A vssd1 vssd1 vccd1 vccd1 _10565_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12304_ _12340_/A _12340_/C vssd1 vssd1 vccd1 vccd1 _12304_/X sky130_fd_sc_hd__xor2_1
X_16072_ _16072_/A _16072_/B vssd1 vssd1 vccd1 vccd1 _16072_/X sky130_fd_sc_hd__or2_1
X_13284_ _13283_/X _18443_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _13285_/A sky130_fd_sc_hd__mux2_1
X_10496_ _10492_/X _10494_/X _10495_/X _10553_/A _09563_/A vssd1 vssd1 vccd1 vccd1
+ _10502_/B sky130_fd_sc_hd__o221a_1
XFILLER_154_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09927__C1 _09862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15023_ _14937_/X _14924_/X _15023_/S vssd1 vssd1 vccd1 vccd1 _15023_/X sky130_fd_sc_hd__mux2_1
X_19900_ _19900_/CLK _19900_/D vssd1 vssd1 vccd1 vccd1 _19900_/Q sky130_fd_sc_hd__dfxtp_1
X_12235_ _11997_/X _12233_/X _12234_/X vssd1 vssd1 vccd1 vccd1 _12235_/X sky130_fd_sc_hd__a21o_2
XFILLER_154_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10537__B1 _09913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19831_ _19976_/CLK _19831_/D vssd1 vssd1 vccd1 vccd1 _19831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12166_ _12135_/X _12164_/X _12165_/X vssd1 vssd1 vccd1 vccd1 _12167_/B sky130_fd_sc_hd__o21ai_1
XFILLER_110_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold2_A hold2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ _11088_/A _11116_/X _11095_/X vssd1 vssd1 vccd1 vccd1 _11117_/Y sky130_fd_sc_hd__o21ai_1
X_19762_ _20023_/CLK _19762_/D vssd1 vssd1 vccd1 vccd1 _19762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16974_ _16974_/A vssd1 vssd1 vccd1 vccd1 _19444_/D sky130_fd_sc_hd__clkbuf_1
X_12097_ _12193_/A _12279_/B _12279_/C _12094_/X vssd1 vssd1 vccd1 vccd1 _12097_/X
+ sky130_fd_sc_hd__o31a_1
X_18713_ _18993_/CLK _18713_/D vssd1 vssd1 vccd1 vccd1 _18713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15925_ _15940_/A _15955_/A _15925_/C vssd1 vssd1 vccd1 vccd1 _15925_/X sky130_fd_sc_hd__and3_1
X_11048_ _19231_/Q _19726_/Q _11048_/S vssd1 vssd1 vccd1 vccd1 _11048_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19693_ _19693_/CLK _19693_/D vssd1 vssd1 vccd1 vccd1 _19693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 io_dbus_rdata[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_4
XFILLER_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10935__S1 _10663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15856_ _15856_/A vssd1 vssd1 vccd1 vccd1 _15856_/X sky130_fd_sc_hd__buf_2
XFILLER_37_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18644_ _18653_/CLK _18644_/D vssd1 vssd1 vccd1 vccd1 _18644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09323__A _09468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14807_ _14813_/B _14807_/B _14807_/C _14807_/D vssd1 vssd1 vccd1 vccd1 _14808_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_149_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15787_ _19880_/D _15787_/B vssd1 vssd1 vccd1 vccd1 _15879_/A sky130_fd_sc_hd__nor2_2
XANTENNA__16855__S _16859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18575_ _19023_/CLK _18575_/D vssd1 vssd1 vccd1 vccd1 _18575_/Q sky130_fd_sc_hd__dfxtp_1
X_12999_ _12936_/A _12994_/X _12996_/Y _12998_/X vssd1 vssd1 vccd1 vccd1 _12999_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12462__A0 _15952_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17526_ _19669_/Q vssd1 vssd1 vccd1 vccd1 _17527_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_45_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14738_ _18819_/Q _13733_/X _14738_/S vssd1 vssd1 vccd1 vccd1 _14739_/A sky130_fd_sc_hd__mux2_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17457_ _17141_/X _19636_/Q _17459_/S vssd1 vssd1 vccd1 vccd1 _17458_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14669_ _14669_/A vssd1 vssd1 vccd1 vccd1 _18788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16408_ _16408_/A vssd1 vssd1 vccd1 vccd1 _19193_/D sky130_fd_sc_hd__clkbuf_1
X_17388_ _17388_/A vssd1 vssd1 vccd1 vccd1 _19605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10916__B _12837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17686__S _17698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_164_clock clkbuf_opt_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _18958_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16339_ _17675_/A vssd1 vssd1 vccd1 vccd1 _16339_/X sky130_fd_sc_hd__clkbuf_2
X_19127_ _19976_/CLK _19127_/D vssd1 vssd1 vccd1 vccd1 _19127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19058_ _19062_/CLK _19058_/D vssd1 vssd1 vccd1 vccd1 _19058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18009_ _19871_/Q _17071_/X _18009_/S vssd1 vssd1 vccd1 vccd1 _18010_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15219__B _15219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10651__B _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_102_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19936_/CLK sky130_fd_sc_hd__clkbuf_16
X_09713_ _10434_/A vssd1 vssd1 vccd1 vccd1 _10294_/A sky130_fd_sc_hd__buf_2
XFILLER_56_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14690__A1 _14548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11763__A _11831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ _09868_/A _09643_/X _09568_/X vssd1 vssd1 vccd1 vccd1 _09644_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10700__B1 _09912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09575_ _10723_/A vssd1 vssd1 vccd1 vccd1 _10670_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_117_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19023_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17450__A _17496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_64_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11103__S1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18281__A _18337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11003__A _11003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10350_ _10351_/A _12854_/B vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__and2_1
XFILLER_3_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10281_ _10290_/A _10280_/X _10162_/X vssd1 vssd1 vccd1 vccd1 _10281_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16005__S _16009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14314__A _18670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12020_ _18759_/Q vssd1 vssd1 vccd1 vccd1 _12020_/X sky130_fd_sc_hd__buf_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13971_ _18564_/Q _13973_/C _13970_/Y vssd1 vssd1 vccd1 vccd1 _18564_/D sky130_fd_sc_hd__o21a_1
XFILLER_120_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14681__A1 _11801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15710_ _18931_/Q _15740_/B vssd1 vssd1 vccd1 vccd1 _15710_/X sky130_fd_sc_hd__or2_1
XFILLER_58_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12922_ _13386_/A vssd1 vssd1 vccd1 vccd1 _13502_/S sky130_fd_sc_hd__buf_4
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16690_ _16690_/A vssd1 vssd1 vccd1 vccd1 _19319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15641_ _15641_/A vssd1 vssd1 vccd1 vccd1 _18899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12853_ _12857_/A _12853_/B vssd1 vssd1 vccd1 vccd1 _12853_/Y sky130_fd_sc_hd__nor2_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _14771_/B vssd1 vssd1 vccd1 vccd1 _15762_/A sky130_fd_sc_hd__buf_2
X_18360_ _18360_/A vssd1 vssd1 vccd1 vccd1 _20011_/D sky130_fd_sc_hd__clkbuf_1
X_15572_ _13535_/A _18901_/Q _15578_/S vssd1 vssd1 vccd1 vccd1 _15573_/A sky130_fd_sc_hd__mux2_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12784_/A _15542_/B vssd1 vssd1 vccd1 vccd1 _12785_/A sky130_fd_sc_hd__xnor2_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17311_ _17138_/X _19571_/Q _17315_/S vssd1 vssd1 vccd1 vccd1 _17312_/A sky130_fd_sc_hd__mux2_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _18741_/Q _14520_/B _14522_/Y vssd1 vssd1 vccd1 vccd1 _18741_/D sky130_fd_sc_hd__o21a_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11735_ _13082_/A vssd1 vssd1 vccd1 vccd1 _11855_/B sky130_fd_sc_hd__buf_2
X_18291_ _17649_/X _19981_/Q _18291_/S vssd1 vssd1 vccd1 vccd1 _18292_/A sky130_fd_sc_hd__mux2_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 _19972_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17242_/A vssd1 vssd1 vccd1 vccd1 _19540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14454_ _14472_/A _14459_/C vssd1 vssd1 vccd1 vccd1 _14454_/Y sky130_fd_sc_hd__nor2_1
X_11666_ _11660_/A _14805_/A _11657_/Y vssd1 vssd1 vccd1 vccd1 _11975_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__15933__A1 _15053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13405_ _17078_/A vssd1 vssd1 vccd1 vccd1 _17720_/A sky130_fd_sc_hd__clkbuf_2
X_17173_ _17710_/A vssd1 vssd1 vccd1 vccd1 _17173_/X sky130_fd_sc_hd__clkbuf_2
X_10617_ _10960_/A vssd1 vssd1 vccd1 vccd1 _10618_/A sky130_fd_sc_hd__clkbuf_4
X_14385_ _14385_/A _14385_/B _14390_/B vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__and3_1
XFILLER_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10758__B1 _09912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11597_ _10761_/B _11616_/B _10759_/X vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__a21o_1
XFILLER_10_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16124_ _16135_/A vssd1 vssd1 vccd1 vccd1 _16133_/S sky130_fd_sc_hd__buf_6
XFILLER_116_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13336_ _14086_/B _09402_/D _09405_/B _18636_/Q _13335_/X vssd1 vssd1 vccd1 vccd1
+ _13336_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_96_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19935_/CLK sky130_fd_sc_hd__clkbuf_16
X_10548_ _19145_/Q _19406_/Q _19305_/Q _19640_/Q _09652_/A _10497_/A vssd1 vssd1 vccd1
+ vccd1 _10549_/B sky130_fd_sc_hd__mux4_1
XFILLER_155_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16055_ _13481_/X _19056_/Q _16057_/S vssd1 vssd1 vccd1 vccd1 _16056_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13267_ _18883_/Q _18884_/Q _13267_/C vssd1 vssd1 vccd1 vccd1 _13288_/B sky130_fd_sc_hd__and3_1
X_10479_ _19932_/Q _19546_/Q _19996_/Q _19115_/Q _09729_/A _10473_/X vssd1 vssd1 vccd1
+ vccd1 _10480_/B sky130_fd_sc_hd__mux4_1
XFILLER_29_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15006_ _14977_/X _15546_/B _15003_/X _15005_/X vssd1 vssd1 vccd1 vccd1 _15006_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13172__A1 _13609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10605__S0 _10724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12218_ _12185_/A _12217_/Y _12182_/B vssd1 vssd1 vccd1 vccd1 _12218_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13198_ _13188_/X _13619_/B _13197_/X _13289_/A vssd1 vssd1 vccd1 vccd1 _13198_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19814_ _19846_/CLK _19814_/D vssd1 vssd1 vccd1 vccd1 _19814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12149_ _12122_/B _12124_/B _12120_/X vssd1 vssd1 vccd1 vccd1 _12184_/A sky130_fd_sc_hd__a21oi_2
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10930__B1 _09873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19745_ _19939_/CLK _19745_/D vssd1 vssd1 vccd1 vccd1 _19745_/Q sky130_fd_sc_hd__dfxtp_1
X_16957_ _16957_/A vssd1 vssd1 vccd1 vccd1 _19436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16949__A0 _16339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ _18996_/Q _15907_/X _15914_/S vssd1 vssd1 vccd1 vccd1 _15909_/A sky130_fd_sc_hd__mux2_1
X_19676_ _19836_/CLK _19676_/D vssd1 vssd1 vccd1 vccd1 _19676_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_34_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19664_/CLK sky130_fd_sc_hd__clkbuf_16
X_16888_ _16355_/X _19406_/Q _16892_/S vssd1 vssd1 vccd1 vccd1 _16889_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18627_ _18660_/CLK _18627_/D vssd1 vssd1 vccd1 vccd1 _18627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16585__S _16591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15839_ input39/X _15834_/X _15789_/X _09280_/Y vssd1 vssd1 vccd1 vccd1 _15840_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _18755_/Q _18751_/Q _18789_/Q _18756_/Q vssd1 vssd1 vccd1 vccd1 _12064_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14975__A2 _15482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18558_ _18741_/CLK _18558_/D vssd1 vssd1 vccd1 vccd1 _18558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12986__A1 _12134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__S1 _11208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17509_ _17509_/A vssd1 vssd1 vccd1 vccd1 _19660_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_49_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19959_/CLK sky130_fd_sc_hd__clkbuf_16
X_09291_ _09315_/B vssd1 vssd1 vccd1 vccd1 _14819_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18489_ _19948_/CLK _18489_/D vssd1 vssd1 vccd1 vccd1 _18489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13303__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11097__S0 _11023_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18305__S _18313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10844__S0 _10859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput120 _12824_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[1] sky130_fd_sc_hd__buf_2
XANTENNA__14134__A _14143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput131 _12825_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[2] sky130_fd_sc_hd__buf_2
Xoutput142 _11918_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_115_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput153 _13864_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_82_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput164 _12028_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10072__S1 _10057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15860__B1 _15788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09627_ _10557_/A vssd1 vssd1 vccd1 vccd1 _10462_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16495__S _16497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17180__A _17180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09558_ _11003_/A vssd1 vssd1 vccd1 vccd1 _09559_/A sky130_fd_sc_hd__buf_2
XFILLER_102_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09489_ _09489_/A vssd1 vssd1 vccd1 vccd1 _19486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14309__A _18669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ _11589_/A _11626_/A _11589_/C _10445_/A _11519_/X vssd1 vssd1 vccd1 vccd1
+ _11586_/C sky130_fd_sc_hd__a311o_1
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ _11960_/A _12823_/B _11967_/A _11450_/X vssd1 vssd1 vccd1 vccd1 _11607_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17117__A0 _17115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18215__S _18219_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10402_ _10448_/A _10401_/X _10557_/A vssd1 vssd1 vccd1 vccd1 _10402_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10835__S0 _11467_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14170_ _18628_/Q _14172_/C _14169_/Y vssd1 vssd1 vccd1 vccd1 _18628_/D sky130_fd_sc_hd__o21a_1
XFILLER_164_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11382_ _20010_/Q _19848_/Q _19257_/Q _19027_/Q _11124_/A _11077_/A vssd1 vssd1 vccd1
+ vccd1 _11382_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ _18688_/Q vssd1 vssd1 vccd1 vccd1 _14378_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10333_ _10329_/X _10331_/X _10332_/X _10290_/A _10162_/X vssd1 vssd1 vccd1 vccd1
+ _10333_/X sky130_fd_sc_hd__o221a_1
XANTENNA__10572__A _10572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15143__A2 _15138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14044__A _14044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13154__A1 _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input54_A io_ibus_inst[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ _19888_/Q _13164_/B _13050_/X _13051_/X vssd1 vssd1 vccd1 vccd1 _13053_/B
+ sky130_fd_sc_hd__a211o_1
X_10264_ _09567_/A _10257_/X _10259_/X _10263_/X _09555_/A vssd1 vssd1 vccd1 vccd1
+ _10264_/X sky130_fd_sc_hd__a221o_2
XFILLER_121_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14979__A _14993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12003_ _12003_/A _12003_/B _12003_/C _09482_/B vssd1 vssd1 vccd1 vccd1 _12004_/D
+ sky130_fd_sc_hd__or4b_1
XANTENNA__17355__A _17411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17860_ _17860_/A vssd1 vssd1 vccd1 vccd1 _19804_/D sky130_fd_sc_hd__clkbuf_1
X_10195_ _19939_/Q _19553_/Q _20003_/Q _19122_/Q _10354_/S _10182_/X vssd1 vssd1 vccd1
+ vccd1 _10196_/B sky130_fd_sc_hd__mux4_1
XFILLER_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16811_ _16364_/X _19372_/Q _16819_/S vssd1 vssd1 vccd1 vccd1 _16812_/A sky130_fd_sc_hd__mux2_1
X_17791_ _17710_/X _19774_/Q _17793_/S vssd1 vssd1 vccd1 vccd1 _17792_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19530_ _19980_/CLK _19530_/D vssd1 vssd1 vccd1 vccd1 _19530_/Q sky130_fd_sc_hd__dfxtp_1
X_16742_ _16742_/A vssd1 vssd1 vccd1 vccd1 _19341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13954_ _14094_/A vssd1 vssd1 vccd1 vccd1 _13991_/A sky130_fd_sc_hd__buf_2
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12905_ _13092_/A _12904_/Y _19487_/Q _09342_/B vssd1 vssd1 vccd1 vccd1 _12906_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16673_ _16673_/A vssd1 vssd1 vccd1 vccd1 _19311_/D sky130_fd_sc_hd__clkbuf_1
X_19461_ _19855_/CLK _19461_/D vssd1 vssd1 vccd1 vccd1 _19461_/Q sky130_fd_sc_hd__dfxtp_1
X_13885_ _15769_/A vssd1 vssd1 vccd1 vccd1 _13885_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18412_ _17720_/X _20035_/Q _18418_/S vssd1 vssd1 vccd1 vccd1 _18413_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17090__A _17090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12836_ _12836_/A vssd1 vssd1 vccd1 vccd1 _12836_/X sky130_fd_sc_hd__clkbuf_2
X_15624_ _15624_/A vssd1 vssd1 vccd1 vccd1 _15901_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__12417__B1 _12416_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _19980_/CLK _19392_/D vssd1 vssd1 vccd1 vccd1 _19392_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18343_ _18343_/A vssd1 vssd1 vccd1 vccd1 _20004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15555_ _15552_/Y _15209_/X _15554_/X _15216_/X vssd1 vssd1 vccd1 vccd1 _15555_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12745_/A _12768_/C _18547_/Q vssd1 vssd1 vccd1 vccd1 _12769_/A sky130_fd_sc_hd__a21oi_1
XFILLER_43_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _18735_/Q _14503_/B _14505_/Y vssd1 vssd1 vccd1 vccd1 _18735_/D sky130_fd_sc_hd__o21a_1
X_18274_ _19974_/Q _17729_/A _18274_/S vssd1 vssd1 vccd1 vccd1 _18275_/A sky130_fd_sc_hd__mux2_1
X_11718_ _18824_/Q vssd1 vssd1 vccd1 vccd1 _13747_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15486_ _15077_/X _15483_/Y _15485_/X _14855_/A vssd1 vssd1 vccd1 vccd1 _15489_/B
+ sky130_fd_sc_hd__a211o_1
X_12698_ _18480_/Q _12556_/X _12557_/X vssd1 vssd1 vccd1 vccd1 _12698_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_174_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14437_ _18706_/Q _14439_/C _14436_/Y vssd1 vssd1 vccd1 vccd1 _18706_/D sky130_fd_sc_hd__o21a_1
X_17225_ _17225_/A vssd1 vssd1 vccd1 vccd1 _19532_/D sky130_fd_sc_hd__clkbuf_1
X_11649_ _11582_/X _11584_/Y _11636_/X _11639_/Y _11648_/X vssd1 vssd1 vccd1 vccd1
+ _11649_/X sky130_fd_sc_hd__a2111o_1
Xinput11 io_dbus_rdata[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_4
XANTENNA__14653__S _14667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput22 io_dbus_rdata[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12962__A _17001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15976__C _15976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput33 io_dbus_valid vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_6
XFILLER_156_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17156_ _17156_/A vssd1 vssd1 vccd1 vccd1 _19507_/D sky130_fd_sc_hd__clkbuf_1
Xinput44 io_ibus_inst[19] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10826__S0 _11467_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14368_ _14371_/B _14365_/C _14367_/Y vssd1 vssd1 vccd1 vccd1 _18686_/D sky130_fd_sc_hd__o21a_1
Xinput55 io_ibus_inst[29] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_4
Xinput66 io_ibus_valid vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_8
XFILLER_156_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16107_ _13161_/X _19076_/Q _16111_/S vssd1 vssd1 vccd1 vccd1 _16108_/A sky130_fd_sc_hd__mux2_1
X_13319_ _13319_/A vssd1 vssd1 vccd1 vccd1 _13319_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11943__A2 _12831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17087_ _17087_/A vssd1 vssd1 vccd1 vccd1 _17087_/X sky130_fd_sc_hd__clkbuf_2
X_14299_ _18665_/Q _14295_/B _14298_/Y vssd1 vssd1 vccd1 vccd1 _18665_/D sky130_fd_sc_hd__o21a_1
X_16038_ _13344_/X _19048_/Q _16042_/S vssd1 vssd1 vccd1 vccd1 _16039_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14889__A _14931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13696__A2 _11898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18084__A1 _11724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11251__S0 _10977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17989_ _18011_/A vssd1 vssd1 vccd1 vccd1 _17998_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_123_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19728_ _20018_/CLK _19728_/D vssd1 vssd1 vccd1 vccd1 _19728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10667__C1 _09686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17595__A0 _17144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19659_ _19755_/CLK _19659_/D vssd1 vssd1 vccd1 vccd1 _19659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09412_ _15779_/A _09411_/Y _18710_/Q vssd1 vssd1 vccd1 vccd1 _09412_/X sky130_fd_sc_hd__o21ba_1
XFILLER_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12856__B _12856_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09343_ _09305_/X _09339_/X _09342_/X vssd1 vssd1 vccd1 vccd1 _09442_/B sky130_fd_sc_hd__o21a_2
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09274_ _09274_/A _09502_/A _09316_/A vssd1 vssd1 vccd1 vccd1 _09274_/X sky130_fd_sc_hd__or3_1
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18035__S _18044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12872__A _19487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14581__A0 _18763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10198__A1 _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12591__B _15449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17874__S _17876_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10293__S1 _10329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__S0 _10797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13687__A2 _13517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14636__A1 _13685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09405__B _09405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10951_ _19664_/Q _19430_/Q _18495_/Q _19760_/Q _10907_/S _10624_/A vssd1 vssd1 vccd1
+ vccd1 _10952_/B sky130_fd_sc_hd__mux4_1
XFILLER_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13670_ _18474_/Q _13669_/X _13670_/S vssd1 vssd1 vccd1 vccd1 _13671_/A sky130_fd_sc_hd__mux2_1
X_10882_ _11473_/A _10882_/B vssd1 vssd1 vccd1 vccd1 _10882_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12621_ _12621_/A _12621_/B vssd1 vssd1 vccd1 vccd1 _12621_/X sky130_fd_sc_hd__xor2_4
XANTENNA__16953__S _16953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ _15399_/A _15340_/B _15340_/C vssd1 vssd1 vccd1 vccd1 _15340_/X sky130_fd_sc_hd__and3_1
X_12552_ _18538_/Q vssd1 vssd1 vccd1 vccd1 _12554_/A sky130_fd_sc_hd__buf_2
XFILLER_157_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11503_ _20022_/Q _19860_/Q _19269_/Q _19039_/Q _11488_/S _10856_/X vssd1 vssd1 vccd1
+ vccd1 _11503_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10830__C1 _09874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15271_ _15218_/X _15265_/Y _15270_/Y vssd1 vssd1 vccd1 vccd1 _15272_/C sky130_fd_sc_hd__a21oi_1
XFILLER_156_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12483_ _18774_/Q _18773_/Q _12483_/C vssd1 vssd1 vccd1 vccd1 _12532_/C sky130_fd_sc_hd__and3_2
XANTENNA__16561__A1 _13774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17010_ _17010_/A vssd1 vssd1 vccd1 vccd1 _17010_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14222_ _18946_/Q _18945_/Q _18944_/Q _14222_/D vssd1 vssd1 vccd1 vccd1 _14227_/C
+ sky130_fd_sc_hd__or4_1
X_11434_ _20009_/Q _19847_/Q _19256_/Q _19026_/Q _11154_/A _11107_/A vssd1 vssd1 vccd1
+ vccd1 _11435_/B sky130_fd_sc_hd__mux4_1
XFILLER_22_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11386__B1 _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153_ _18623_/Q _14153_/B _14153_/C vssd1 vssd1 vccd1 vccd1 _14154_/C sky130_fd_sc_hd__and3_1
XFILLER_164_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10284__S1 _10283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11365_ _19656_/Q _19422_/Q _18487_/Q _19752_/Q _11124_/A _11077_/A vssd1 vssd1 vccd1
+ vccd1 _11366_/B sky130_fd_sc_hd__mux4_1
XFILLER_113_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13104_ _18799_/Q _12880_/X _12984_/A _18766_/Q _13103_/X vssd1 vssd1 vccd1 vccd1
+ _13104_/X sky130_fd_sc_hd__a221o_2
X_10316_ _10054_/A _10313_/X _10315_/X vssd1 vssd1 vccd1 vccd1 _10316_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14084_ _14086_/B _14086_/C _14059_/X vssd1 vssd1 vccd1 vccd1 _14084_/Y sky130_fd_sc_hd__a21oi_1
X_18961_ _18967_/CLK _18961_/D vssd1 vssd1 vccd1 vccd1 _18961_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output160_A _12703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11296_ _11296_/A _11296_/B vssd1 vssd1 vccd1 vccd1 _11296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13678__A2 _13677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13817__S _13820_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17912_ _17912_/A vssd1 vssd1 vccd1 vccd1 _19827_/D sky130_fd_sc_hd__clkbuf_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _18556_/Q _13189_/A _13031_/X _13033_/X _13034_/X vssd1 vssd1 vccd1 vccd1
+ _13551_/B sky130_fd_sc_hd__a2111o_4
XFILLER_65_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10247_ _10106_/Y _11642_/B _11640_/B _11640_/A vssd1 vssd1 vccd1 vccd1 _10247_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__12721__S _12814_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12886__B1 _12879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18892_ _18926_/CLK _18892_/D vssd1 vssd1 vccd1 vccd1 _18892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_186_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17843_ _19797_/Q _17039_/X _17843_/S vssd1 vssd1 vccd1 vccd1 _17844_/A sky130_fd_sc_hd__mux2_1
X_10178_ _11640_/A vssd1 vssd1 vccd1 vccd1 _10179_/B sky130_fd_sc_hd__inv_2
XFILLER_121_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13118__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17774_ _17684_/X _19766_/Q _17782_/S vssd1 vssd1 vccd1 vccd1 _17775_/A sky130_fd_sc_hd__mux2_1
X_14986_ _15097_/A vssd1 vssd1 vccd1 vccd1 _14986_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19513_ _19868_/CLK _19513_/D vssd1 vssd1 vccd1 vccd1 _19513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16725_ _19334_/Q _13803_/X _16725_/S vssd1 vssd1 vccd1 vccd1 _16726_/A sky130_fd_sc_hd__mux2_1
X_13937_ _13946_/A _13937_/B _13937_/C vssd1 vssd1 vccd1 vccd1 _18553_/D sky130_fd_sc_hd__nor3_1
XFILLER_74_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17024__S _17024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19444_ _19936_/CLK _19444_/D vssd1 vssd1 vccd1 vccd1 _19444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16656_ _16656_/A vssd1 vssd1 vccd1 vccd1 _19303_/D sky130_fd_sc_hd__clkbuf_1
X_13868_ _12790_/X _12024_/Y _12027_/X _17203_/A vssd1 vssd1 vccd1 vccd1 _18520_/D
+ sky130_fd_sc_hd__a211o_1
X_15607_ _13664_/A _18917_/Q _15611_/S vssd1 vssd1 vccd1 vccd1 _15608_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17959__S _17965_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ _18788_/Q _12799_/A _12799_/B _12818_/Y _13650_/A vssd1 vssd1 vccd1 vccd1
+ _12820_/B sky130_fd_sc_hd__a311o_1
X_19375_ _20003_/CLK _19375_/D vssd1 vssd1 vccd1 vccd1 _19375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16587_ _19273_/Q _13813_/X _16591_/S vssd1 vssd1 vccd1 vccd1 _16588_/A sky130_fd_sc_hd__mux2_1
X_13799_ _13799_/A vssd1 vssd1 vccd1 vccd1 _18498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18326_ _18337_/A vssd1 vssd1 vccd1 vccd1 _18335_/S sky130_fd_sc_hd__buf_4
XFILLER_148_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11613__B2 _11462_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _15542_/A _15542_/B vssd1 vssd1 vccd1 vccd1 _15538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18257_ _19966_/Q _17704_/A _18263_/S vssd1 vssd1 vccd1 vccd1 _18258_/A sky130_fd_sc_hd__mux2_1
X_15469_ _18856_/Q _15457_/X _15468_/X vssd1 vssd1 vccd1 vccd1 _18856_/D sky130_fd_sc_hd__o21a_1
XANTENNA__16164__A _16221_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17208_ _17208_/A _17208_/B vssd1 vssd1 vccd1 vccd1 _17209_/A sky130_fd_sc_hd__and2_1
XFILLER_128_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18188_ _18188_/A vssd1 vssd1 vccd1 vccd1 _19935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17139_ _17138_/X _19502_/Q _17145_/S vssd1 vssd1 vccd1 vccd1 _17140_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11472__S0 _10776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09961_ _18861_/Q vssd1 vssd1 vccd1 vccd1 _09961_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18057__A1 _13572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11224__S0 _11171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__S1 _09612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16103__S _16111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09892_ _20038_/Q _19876_/Q _19285_/Q _19055_/Q _09733_/X _09768_/X vssd1 vssd1 vccd1
+ vccd1 _09892_/X sky130_fd_sc_hd__mux4_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12629__B1 _12170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15848__A2_N _15834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16339__A _17675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10387__A _10424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16773__S _16775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09326_ _18984_/Q _18983_/Q _18982_/Q _18981_/Q vssd1 vssd1 vccd1 vccd1 _12004_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_22_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09257_ _09502_/A _09501_/B _09499_/B _09248_/X vssd1 vssd1 vccd1 vccd1 _09265_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_166_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09188_ _09188_/A vssd1 vssd1 vccd1 vccd1 _09188_/Y sky130_fd_sc_hd__inv_6
XFILLER_153_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09216__B1_N input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11011__A _18841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ _19198_/Q _19789_/Q _19951_/Q _19166_/Q _09721_/A _10854_/A vssd1 vssd1 vccd1
+ vccd1 _11150_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10101_ _09946_/A _10098_/X _10100_/X vssd1 vssd1 vccd1 vccd1 _10101_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11215__S0 _11125_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ _11081_/A vssd1 vssd1 vccd1 vccd1 _11081_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10032_ _10007_/A _10031_/X _09780_/A vssd1 vssd1 vccd1 vccd1 _10032_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11540__B1 _09690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15806__B1 _15789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14840_ _14966_/A _15004_/A vssd1 vssd1 vccd1 vccd1 _14846_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09850__S _09855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14771_ _14771_/A _14771_/B vssd1 vssd1 vccd1 vccd1 _14778_/A sky130_fd_sc_hd__nor2_2
XFILLER_75_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input17_A io_dbus_rdata[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13293__B1 _11733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11983_ _18983_/Q _11982_/X _11983_/S vssd1 vssd1 vccd1 vccd1 _11983_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16249__A _16295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16510_ _16532_/A vssd1 vssd1 vccd1 vccd1 _16519_/S sky130_fd_sc_hd__buf_4
X_13722_ _18893_/Q _13723_/B vssd1 vssd1 vccd1 vccd1 _13737_/C sky130_fd_sc_hd__or2_1
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ _10934_/A _10934_/B vssd1 vssd1 vccd1 vccd1 _10934_/Y sky130_fd_sc_hd__nor2_1
X_17490_ _17189_/X _19651_/Q _17492_/S vssd1 vssd1 vccd1 vccd1 _17491_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16441_ _16441_/A vssd1 vssd1 vccd1 vccd1 _19208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13653_ _18884_/Q _13654_/B vssd1 vssd1 vccd1 vccd1 _13672_/C sky130_fd_sc_hd__or2_2
X_10865_ _11500_/A _10865_/B vssd1 vssd1 vccd1 vccd1 _10865_/X sky130_fd_sc_hd__or2_1
XANTENNA__16683__S _16685_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13596__A1 _13594_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12604_ _12338_/X _12602_/X _12603_/Y vssd1 vssd1 vccd1 vccd1 _12604_/Y sky130_fd_sc_hd__a21oi_1
X_16372_ _16371_/X _19182_/Q _16378_/S vssd1 vssd1 vccd1 vccd1 _16373_/A sky130_fd_sc_hd__mux2_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19160_ _19720_/CLK _19160_/D vssd1 vssd1 vccd1 vccd1 _19160_/Q sky130_fd_sc_hd__dfxtp_1
X_13584_ _13690_/A vssd1 vssd1 vccd1 vccd1 _13617_/S sky130_fd_sc_hd__buf_2
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _10954_/S vssd1 vssd1 vccd1 vccd1 _10953_/S sky130_fd_sc_hd__clkbuf_4
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18111_ _18857_/Q _11898_/X _18118_/S vssd1 vssd1 vccd1 vccd1 _18111_/X sky130_fd_sc_hd__mux2_1
X_15323_ _15323_/A _15323_/B _15323_/C vssd1 vssd1 vccd1 vccd1 _15323_/X sky130_fd_sc_hd__and3_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _15410_/A _12515_/B _12632_/A vssd1 vssd1 vccd1 vccd1 _12541_/A sky130_fd_sc_hd__o21a_1
X_19091_ _19942_/CLK _19091_/D vssd1 vssd1 vccd1 vccd1 _19091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18042_ _18042_/A vssd1 vssd1 vccd1 vccd1 _19884_/D sky130_fd_sc_hd__clkbuf_1
X_15254_ _15254_/A _15254_/B vssd1 vssd1 vccd1 vccd1 _15254_/Y sky130_fd_sc_hd__nor2_1
X_12466_ _12466_/A vssd1 vssd1 vccd1 vccd1 _12469_/A sky130_fd_sc_hd__clkinv_2
XFILLER_173_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14205_ _18640_/Q _14207_/C _14204_/Y vssd1 vssd1 vccd1 vccd1 _18640_/D sky130_fd_sc_hd__o21a_1
XFILLER_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ _11206_/A _11416_/X _09681_/A vssd1 vssd1 vccd1 vccd1 _11417_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15185_ _15348_/S _15244_/A _14835_/Y vssd1 vssd1 vccd1 vccd1 _15491_/B sky130_fd_sc_hd__a21o_1
XANTENNA__18403__S _18407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12397_ _18468_/Q _12012_/X _13648_/A vssd1 vssd1 vccd1 vccd1 _12397_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output85_A _12599_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14136_ _14144_/D vssd1 vssd1 vccd1 vccd1 _14142_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11348_ _19354_/Q _19689_/Q _11348_/S vssd1 vssd1 vccd1 vccd1 _11348_/X sky130_fd_sc_hd__mux2_1
X_19993_ _19993_/CLK _19993_/D vssd1 vssd1 vccd1 vccd1 _19993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14067_ _18597_/Q _14064_/B _14066_/Y vssd1 vssd1 vccd1 vccd1 _18597_/D sky130_fd_sc_hd__o21a_1
X_18944_ _18967_/CLK _18944_/D vssd1 vssd1 vccd1 vccd1 _18944_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10760__A _10760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ _19323_/Q _19594_/Q _19818_/Q _19562_/Q _11125_/S _11065_/X vssd1 vssd1 vccd1
+ vccd1 _11279_/X sky130_fd_sc_hd__mux4_1
X_13018_ _18867_/Q _12973_/B _13535_/A _13554_/A vssd1 vssd1 vccd1 vccd1 _13019_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_67_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18875_ _18878_/CLK _18875_/D vssd1 vssd1 vccd1 vccd1 _18875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17826_ _19789_/Q _17014_/X _17832_/S vssd1 vssd1 vccd1 vccd1 _17827_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17757_ _17757_/A vssd1 vssd1 vccd1 vccd1 _19758_/D sky130_fd_sc_hd__clkbuf_1
X_14969_ _15553_/B _14973_/A vssd1 vssd1 vccd1 vccd1 _14970_/D sky130_fd_sc_hd__nor2_1
XFILLER_63_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16708_ _19326_/Q _13778_/X _16714_/S vssd1 vssd1 vccd1 vccd1 _16709_/A sky130_fd_sc_hd__mux2_1
X_17688_ _17688_/A vssd1 vssd1 vccd1 vccd1 _17688_/X sky130_fd_sc_hd__buf_2
XFILLER_23_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17689__S _17698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19427_ _19757_/CLK _19427_/D vssd1 vssd1 vccd1 vccd1 _19427_/Q sky130_fd_sc_hd__dfxtp_1
X_16639_ _16326_/X _19296_/Q _16641_/S vssd1 vssd1 vccd1 vccd1 _16640_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19358_ _19758_/CLK _19358_/D vssd1 vssd1 vccd1 vccd1 _19358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09886__S0 _11553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18309_ _17675_/X _19989_/Q _18313_/S vssd1 vssd1 vccd1 vccd1 _18310_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19289_ _19389_/CLK _19289_/D vssd1 vssd1 vccd1 vccd1 _19289_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14407__A _14407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14536__A0 _14548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11445__S0 _11154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18313__S _18313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16289__A0 _13443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ _09946_/A _09943_/X _09809_/A vssd1 vssd1 vccd1 vccd1 _09944_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09875_ _09875_/A vssd1 vssd1 vccd1 vccd1 _09876_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A io_dbus_rdata[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10325__A1 _10194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_134_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ _18849_/Q _09843_/A _09883_/A _10649_/X vssd1 vssd1 vccd1 vccd1 _12847_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_16_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09309_ _09309_/A _09316_/A _09316_/B vssd1 vssd1 vccd1 vccd1 _14813_/B sky130_fd_sc_hd__nor3_2
XFILLER_70_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10581_ _10520_/A _10577_/X _10580_/X vssd1 vssd1 vccd1 vccd1 _10581_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_155_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12320_ _11904_/A _12841_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _12406_/A sky130_fd_sc_hd__a21oi_1
XFILLER_126_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12251_ _12479_/S _12249_/Y _12250_/X _12154_/X vssd1 vssd1 vccd1 vccd1 _12251_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10056__S _10254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11202_ _10983_/X _11200_/X _11425_/A vssd1 vssd1 vccd1 vccd1 _11202_/X sky130_fd_sc_hd__a21o_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _12182_/A _12182_/B vssd1 vssd1 vccd1 vccd1 _12215_/D sky130_fd_sc_hd__nor2_2
XFILLER_134_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11676__A _12060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _11133_/A _11133_/B _11133_/C vssd1 vssd1 vccd1 vccd1 _11133_/X sky130_fd_sc_hd__or3_1
X_16990_ _16399_/X _19452_/Q _16990_/S vssd1 vssd1 vccd1 vccd1 _16991_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11064_ _19523_/Q vssd1 vssd1 vccd1 vccd1 _11073_/A sky130_fd_sc_hd__buf_2
X_15941_ _19007_/Q _15921_/X _15940_/X vssd1 vssd1 vccd1 vccd1 _19007_/D sky130_fd_sc_hd__a21o_1
XFILLER_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10316__A1 _10054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_59_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10015_ _10294_/A _10014_/X _09799_/A vssd1 vssd1 vccd1 vccd1 _10015_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18660_ _18660_/CLK _18660_/D vssd1 vssd1 vccd1 vccd1 _18660_/Q sky130_fd_sc_hd__dfxtp_1
X_15872_ _09466_/A _15856_/X _15788_/X input50/X vssd1 vssd1 vccd1 vccd1 _16844_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17611_ _17167_/X _19708_/Q _17617_/S vssd1 vssd1 vccd1 vccd1 _17612_/A sky130_fd_sc_hd__mux2_1
X_14823_ _14956_/S _15004_/B vssd1 vssd1 vccd1 vccd1 _14973_/B sky130_fd_sc_hd__or2_2
X_18591_ _18724_/CLK _18591_/D vssd1 vssd1 vccd1 vccd1 _18591_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13266__B1 _18884_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output123_A _12854_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17542_ _19677_/Q vssd1 vssd1 vccd1 vccd1 _17543_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_45_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14754_ _09276_/X _09516_/B _14753_/X vssd1 vssd1 vccd1 vccd1 _14815_/C sky130_fd_sc_hd__o21ai_2
X_11966_ _12078_/B vssd1 vssd1 vccd1 vccd1 _14865_/A sky130_fd_sc_hd__buf_2
XFILLER_72_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ _15934_/B _12837_/B vssd1 vssd1 vccd1 vccd1 _10918_/B sky130_fd_sc_hd__and2_1
XFILLER_60_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13705_ _12422_/X _13704_/X _13514_/S vssd1 vssd1 vccd1 vccd1 _13705_/X sky130_fd_sc_hd__a21bo_1
X_17473_ _17163_/X _19643_/Q _17481_/S vssd1 vssd1 vccd1 vccd1 _17474_/A sky130_fd_sc_hd__mux2_1
X_14685_ _14742_/S vssd1 vssd1 vccd1 vccd1 _14694_/S sky130_fd_sc_hd__buf_2
X_11897_ _11897_/A _19018_/Q vssd1 vssd1 vccd1 vccd1 _11897_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13830__S _13836_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19212_ _19997_/CLK _19212_/D vssd1 vssd1 vccd1 vccd1 _19212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16424_ _19201_/Q _13787_/X _16424_/S vssd1 vssd1 vccd1 vccd1 _16425_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13636_ _18881_/Q _13637_/B vssd1 vssd1 vccd1 vccd1 _13646_/C sky130_fd_sc_hd__or2_2
X_10848_ _11493_/A _10848_/B vssd1 vssd1 vccd1 vccd1 _10848_/X sky130_fd_sc_hd__or2_1
XFILLER_60_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19143_ _19993_/CLK _19143_/D vssd1 vssd1 vccd1 vccd1 _19143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16355_ _17691_/A vssd1 vssd1 vccd1 vccd1 _16355_/X sky130_fd_sc_hd__clkbuf_2
X_13567_ _13700_/A _14548_/A _13566_/Y vssd1 vssd1 vccd1 vccd1 _13567_/X sky130_fd_sc_hd__a21o_1
X_10779_ _19204_/Q _19795_/Q _19957_/Q _19172_/Q _10704_/A _10048_/A vssd1 vssd1 vccd1
+ vccd1 _10780_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15306_ _15306_/A _15306_/B vssd1 vssd1 vccd1 vccd1 _15306_/Y sky130_fd_sc_hd__nor2_1
X_12518_ _12518_/A _14886_/A vssd1 vssd1 vccd1 vccd1 _12546_/A sky130_fd_sc_hd__xnor2_4
X_16286_ _16286_/A vssd1 vssd1 vccd1 vccd1 _19154_/D sky130_fd_sc_hd__clkbuf_1
X_19074_ _19664_/CLK _19074_/D vssd1 vssd1 vccd1 vccd1 _19074_/Q sky130_fd_sc_hd__dfxtp_1
X_13498_ _12960_/A _13485_/Y _13486_/X _13497_/Y _09532_/A vssd1 vssd1 vccd1 vccd1
+ _13498_/X sky130_fd_sc_hd__a311o_2
XFILLER_139_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18025_ _18025_/A vssd1 vssd1 vccd1 vccd1 _19878_/D sky130_fd_sc_hd__clkbuf_1
X_12449_ _18470_/Q _12343_/X _12344_/X vssd1 vssd1 vccd1 vccd1 _12449_/Y sky130_fd_sc_hd__o21ai_1
X_15237_ _15413_/A vssd1 vssd1 vccd1 vccd1 _15400_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15984__C _16846_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13741__A1 _19024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15168_ _15038_/X _15031_/X _15198_/S vssd1 vssd1 vccd1 vccd1 _15168_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10555__A1 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11752__B1 _12890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17972__S _17976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14119_ _18737_/Q _18736_/Q _18738_/Q _14504_/A vssd1 vssd1 vccd1 vccd1 _14513_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_125_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19976_ _19976_/CLK _19976_/D vssd1 vssd1 vccd1 vccd1 _19976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10490__A _15958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15099_ _15099_/A vssd1 vssd1 vccd1 vccd1 _15099_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18927_ _18928_/CLK _18927_/D vssd1 vssd1 vccd1 vccd1 _18927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09660_ _09660_/A _09660_/B vssd1 vssd1 vccd1 vccd1 _09660_/X sky130_fd_sc_hd__and2_1
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18858_ _18858_/CLK _18858_/D vssd1 vssd1 vccd1 vccd1 _18858_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17809_ _17809_/A vssd1 vssd1 vccd1 vccd1 _19782_/D sky130_fd_sc_hd__clkbuf_1
X_09591_ _10724_/S vssd1 vssd1 vccd1 vccd1 _10586_/S sky130_fd_sc_hd__buf_2
X_18789_ _18789_/CLK _18789_/D vssd1 vssd1 vccd1 vccd1 _18789_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11807__B2 _15738_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09859__S0 _09855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12864__B _12866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13041__A _17014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10546__B2 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09927_ _09568_/A _09922_/X _09924_/X _09926_/X _09862_/A vssd1 vssd1 vccd1 vccd1
+ _09927_/X sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_60_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09858_ _19349_/Q _19620_/Q _19844_/Q _19588_/Q _11532_/S _09614_/X vssd1 vssd1 vccd1
+ vccd1 _09858_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _09789_/A vssd1 vssd1 vccd1 vccd1 _11095_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _12881_/A vssd1 vssd1 vccd1 vccd1 _12944_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11728_/C _11748_/X _11750_/X vssd1 vssd1 vccd1 vccd1 _18748_/D sky130_fd_sc_hd__a21o_1
XFILLER_42_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ _10775_/A vssd1 vssd1 vccd1 vccd1 _10703_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10482__B1 _10162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14470_ _14495_/A _14470_/B _14470_/C vssd1 vssd1 vccd1 vccd1 _18722_/D sky130_fd_sc_hd__nor3_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11682_/A vssd1 vssd1 vccd1 vccd1 _13057_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13223_/X _13409_/Y _13420_/X vssd1 vssd1 vccd1 vccd1 _17081_/A sky130_fd_sc_hd__o21ai_2
X_10633_ _10695_/A _10633_/B vssd1 vssd1 vccd1 vccd1 _10633_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16140_ _13423_/X _19091_/Q _16144_/S vssd1 vssd1 vccd1 vccd1 _16141_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13352_ _12967_/X _13350_/X _13351_/X vssd1 vssd1 vccd1 vccd1 _17068_/A sky130_fd_sc_hd__o21a_4
XFILLER_154_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10564_ _18441_/Q _19470_/Q _19507_/Q _19081_/Q _10529_/S _10011_/A vssd1 vssd1 vccd1
+ vccd1 _10564_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10785__A1 _09848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__B2 _18845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _12340_/A _12303_/B vssd1 vssd1 vccd1 vccd1 _12312_/A sky130_fd_sc_hd__or2_1
XFILLER_10_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16071_ _16071_/A vssd1 vssd1 vccd1 vccd1 _19061_/D sky130_fd_sc_hd__clkbuf_1
X_13283_ _17697_/A vssd1 vssd1 vccd1 vccd1 _13283_/X sky130_fd_sc_hd__clkbuf_2
X_10495_ _19673_/Q _19439_/Q _18504_/Q _19769_/Q _09653_/A _10587_/A vssd1 vssd1 vccd1
+ vccd1 _10495_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15022_ _14934_/X _14936_/X _15023_/S vssd1 vssd1 vccd1 vccd1 _15022_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12234_ _12234_/A _12234_/B vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__and2_1
XFILLER_170_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18111__A0 _18857_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10537__A1 _09883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19830_ _20025_/CLK _19830_/D vssd1 vssd1 vccd1 vccd1 _19830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12165_ _12165_/A _16072_/A vssd1 vssd1 vccd1 vccd1 _12165_/X sky130_fd_sc_hd__or2_1
XANTENNA__10632__S1 _10010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11116_ _19327_/Q _19598_/Q _19822_/Q _19566_/Q _11186_/S _11022_/A vssd1 vssd1 vccd1
+ vccd1 _11116_/X sky130_fd_sc_hd__mux4_1
X_19761_ _20021_/CLK _19761_/D vssd1 vssd1 vccd1 vccd1 _19761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16973_ _16374_/X _19444_/Q _16975_/S vssd1 vssd1 vccd1 vccd1 _16974_/A sky130_fd_sc_hd__mux2_1
X_12096_ _18522_/Q _12128_/C vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__xor2_1
XFILLER_122_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17093__A _17093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18712_ _18762_/CLK _18712_/D vssd1 vssd1 vccd1 vccd1 _18712_/Q sky130_fd_sc_hd__dfxtp_1
X_15924_ _19000_/Q _15921_/X _15923_/X vssd1 vssd1 vccd1 vccd1 _19000_/D sky130_fd_sc_hd__a21o_1
X_11047_ _11257_/A _11047_/B vssd1 vssd1 vccd1 vccd1 _11047_/X sky130_fd_sc_hd__or2_1
XFILLER_65_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19692_ _19726_/CLK _19692_/D vssd1 vssd1 vccd1 vccd1 _19692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 io_dbus_rdata[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__13239__A0 _13238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18643_ _18655_/CLK _18643_/D vssd1 vssd1 vccd1 vccd1 _18643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15855_ _15855_/A vssd1 vssd1 vccd1 vccd1 _18979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14806_ _09282_/D _09520_/B _14756_/X _14758_/A vssd1 vssd1 vccd1 vccd1 _14807_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09323__B _17098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18574_ _19909_/CLK _18574_/D vssd1 vssd1 vccd1 vccd1 _18574_/Q sky130_fd_sc_hd__dfxtp_1
X_15786_ _18993_/Q _15786_/B _15690_/A input66/X vssd1 vssd1 vccd1 vccd1 _15787_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12998_ _13535_/A _13015_/C _13145_/A vssd1 vssd1 vccd1 vccd1 _12998_/X sky130_fd_sc_hd__a21o_1
XFILLER_73_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17525_ _17525_/A vssd1 vssd1 vccd1 vccd1 _19668_/D sky130_fd_sc_hd__clkbuf_1
X_14737_ _14737_/A vssd1 vssd1 vccd1 vccd1 _18818_/D sky130_fd_sc_hd__clkbuf_1
X_11949_ _14804_/C _11949_/B _14815_/A _14815_/B vssd1 vssd1 vccd1 vccd1 _11949_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14656__S _14667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17456_ _17456_/A vssd1 vssd1 vccd1 vccd1 _19635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14668_ _15813_/A _14668_/B vssd1 vssd1 vccd1 vccd1 _14669_/A sky130_fd_sc_hd__and2_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16407_ _19193_/Q _13762_/X _16413_/S vssd1 vssd1 vccd1 vccd1 _16408_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _19008_/Q _13619_/B vssd1 vssd1 vccd1 vccd1 _13619_/X sky130_fd_sc_hd__or2_1
X_17387_ _19605_/Q _17039_/X _17387_/S vssd1 vssd1 vccd1 vccd1 _17388_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14599_ _14612_/A _14599_/B vssd1 vssd1 vccd1 vccd1 _14600_/A sky130_fd_sc_hd__and2_1
X_19126_ _20007_/CLK _19126_/D vssd1 vssd1 vccd1 vccd1 _19126_/Q sky130_fd_sc_hd__dfxtp_1
X_16338_ _16338_/A vssd1 vssd1 vccd1 vccd1 _19171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19057_ _19856_/CLK _19057_/D vssd1 vssd1 vccd1 vccd1 _19057_/Q sky130_fd_sc_hd__dfxtp_1
X_16269_ _13283_/X _19147_/Q _16269_/S vssd1 vssd1 vccd1 vccd1 _16270_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18008_ _18008_/A vssd1 vssd1 vccd1 vccd1 _19870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12205__A _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19959_ _19959_/CLK _19959_/D vssd1 vssd1 vccd1 vccd1 _19959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09712_ _10172_/A vssd1 vssd1 vccd1 vccd1 _10434_/A sky130_fd_sc_hd__buf_2
XANTENNA__16111__S _16111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09643_ _18454_/Q _19483_/Q _19520_/Q _19094_/Q _09598_/X _09851_/A vssd1 vssd1 vccd1
+ vccd1 _09643_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10161__C1 _09807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__A1 _09883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13036__A _19488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _11473_/A vssd1 vssd1 vccd1 vccd1 _10723_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11456__A1_N _15925_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18038__S _18044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12594__B _12618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10311__S0 _09655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__A1 _10654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12814__S _12814_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13705__A1 _12422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14902__A0 _14996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10280_ _19678_/Q _19444_/Q _18509_/Q _19774_/Q _10279_/X _10329_/A vssd1 vssd1 vccd1
+ vccd1 _10280_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10650__A1_N _18849_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17906__A _17952_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11192__A1 _11340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19720_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13469__B1 _11843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17117__S _17129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13970_ _18564_/Q _13973_/C _13969_/X vssd1 vssd1 vccd1 vccd1 _13970_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14330__A _14413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _18352_/A _17098_/C vssd1 vssd1 vccd1 vccd1 _13386_/A sky130_fd_sc_hd__or2_4
XANTENNA__16956__S _16964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15640_ _18899_/Q _18520_/Q _15644_/S vssd1 vssd1 vccd1 vccd1 _15641_/A sky130_fd_sc_hd__mux2_1
X_12852_ _12863_/A vssd1 vssd1 vccd1 vccd1 _12857_/A sky130_fd_sc_hd__clkbuf_16
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _18750_/Q _17096_/B _11774_/X _11802_/Y vssd1 vssd1 vccd1 vccd1 _11803_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15571_ _15571_/A vssd1 vssd1 vccd1 vccd1 _18868_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12783_/A vssd1 vssd1 vccd1 vccd1 _15542_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17310_/A vssd1 vssd1 vccd1 vccd1 _19570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11734_ _11734_/A vssd1 vssd1 vccd1 vccd1 _11815_/A sky130_fd_sc_hd__clkbuf_4
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14522_ _14529_/A _14526_/C vssd1 vssd1 vccd1 vccd1 _14522_/Y sky130_fd_sc_hd__nor2_1
X_18290_ _18290_/A vssd1 vssd1 vccd1 vccd1 _19980_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17383__A1 _17033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17787__S _17793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17241_ _17141_/X _19540_/Q _17243_/S vssd1 vssd1 vccd1 vccd1 _17242_/A sky130_fd_sc_hd__mux2_1
X_11665_ _15738_/A _14761_/B _09522_/Y _15740_/A vssd1 vssd1 vccd1 vccd1 _11975_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14453_ _14453_/A vssd1 vssd1 vccd1 vccd1 _14459_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15933__A2 _15928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10616_ _15949_/B vssd1 vssd1 vccd1 vccd1 _10652_/A sky130_fd_sc_hd__inv_2
X_13404_ _13223_/X _13389_/Y _13403_/X vssd1 vssd1 vccd1 vccd1 _17078_/A sky130_fd_sc_hd__o21ai_4
XFILLER_174_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17172_ _17172_/A vssd1 vssd1 vccd1 vccd1 _19512_/D sky130_fd_sc_hd__clkbuf_1
X_14384_ _18691_/Q _18690_/Q _14384_/C vssd1 vssd1 vccd1 vccd1 _14390_/B sky130_fd_sc_hd__nand3_1
XFILLER_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11596_ _11599_/A _11595_/C _11595_/A vssd1 vssd1 vccd1 vccd1 _11596_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10302__S0 _09595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10758__A1 _09882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16123_ _16123_/A vssd1 vssd1 vccd1 vccd1 _19083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13335_ _18668_/Q _13335_/B vssd1 vssd1 vccd1 vccd1 _13335_/X sky130_fd_sc_hd__and2_1
X_10547_ _19337_/Q _19608_/Q _19832_/Q _19576_/Q _09653_/A _10587_/A vssd1 vssd1 vccd1
+ vccd1 _10547_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16054_ _16054_/A vssd1 vssd1 vccd1 vccd1 _19055_/D sky130_fd_sc_hd__clkbuf_1
X_13266_ _13256_/B _13267_/C _18884_/Q vssd1 vssd1 vccd1 vccd1 _13268_/B sky130_fd_sc_hd__a21oi_1
XFILLER_170_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10478_ _10382_/X _10468_/Y _10472_/Y _10477_/Y _09806_/A vssd1 vssd1 vccd1 vccd1
+ _10478_/X sky130_fd_sc_hd__o311a_1
XFILLER_170_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12217_ _12217_/A _14906_/A vssd1 vssd1 vccd1 vccd1 _12217_/Y sky130_fd_sc_hd__nand2_1
X_15005_ _15413_/A vssd1 vssd1 vccd1 vccd1 _15005_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10605__S1 _10654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13197_ _13473_/A _18847_/Q vssd1 vssd1 vccd1 vccd1 _13197_/X sky130_fd_sc_hd__or2_1
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19813_ _19975_/CLK _19813_/D vssd1 vssd1 vccd1 vccd1 _19813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12148_ _12183_/A _14909_/A vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__xnor2_4
XFILLER_150_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10930__A1 _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11864__A _15789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19744_ _19971_/CLK _19744_/D vssd1 vssd1 vccd1 vccd1 _19744_/Q sky130_fd_sc_hd__dfxtp_1
X_16956_ _16348_/X _19436_/Q _16964_/S vssd1 vssd1 vccd1 vccd1 _16957_/A sky130_fd_sc_hd__mux2_1
X_12079_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12080_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_96_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15907_ _11982_/X _11452_/A _15946_/A vssd1 vssd1 vccd1 vccd1 _15907_/X sky130_fd_sc_hd__mux2_1
X_19675_ _19996_/CLK _19675_/D vssd1 vssd1 vccd1 vccd1 _19675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16887_ _16887_/A vssd1 vssd1 vccd1 vccd1 _19405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18626_ _18660_/CLK _18626_/D vssd1 vssd1 vccd1 vccd1 _18626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15838_ _15871_/A _15838_/B vssd1 vssd1 vccd1 vccd1 _18974_/D sky130_fd_sc_hd__nor2_1
XFILLER_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18557_ _19883_/CLK _18557_/D vssd1 vssd1 vccd1 vccd1 _18557_/Q sky130_fd_sc_hd__dfxtp_1
X_15769_ _15769_/A vssd1 vssd1 vccd1 vccd1 _15769_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09300__A1 _16846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17508_ _19660_/Q vssd1 vssd1 vccd1 vccd1 _17509_/A sky130_fd_sc_hd__clkbuf_1
X_09290_ _09290_/A _09290_/B vssd1 vssd1 vccd1 vccd1 _09315_/B sky130_fd_sc_hd__or2_1
XANTENNA__12986__A2 _12984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18488_ _19485_/CLK _18488_/D vssd1 vssd1 vccd1 vccd1 _18488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17439_ _17496_/S vssd1 vssd1 vccd1 vccd1 _17448_/S sky130_fd_sc_hd__buf_2
XFILLER_165_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15924__A2 _15921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11097__S1 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19109_ _19636_/CLK _19109_/D vssd1 vssd1 vccd1 vccd1 _19109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_opt_2_0_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15688__A1 _18542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput110 _12838_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[10] sky130_fd_sc_hd__buf_2
XFILLER_115_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput121 _12851_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[20] sky130_fd_sc_hd__buf_2
Xoutput132 _12865_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[30] sky130_fd_sc_hd__buf_2
Xoutput143 _12288_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[10] sky130_fd_sc_hd__buf_2
Xoutput154 _12564_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[20] sky130_fd_sc_hd__buf_2
Xoutput165 _12801_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[30] sky130_fd_sc_hd__buf_2
XFILLER_142_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14150__A _14159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15860__A1 _09467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12589__B _12854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15860__B2 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17461__A _17483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ _09987_/A vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09557_ _09557_/A vssd1 vssd1 vccd1 vccd1 _11003_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13623__A0 _13621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12426__A1 _12422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09488_ _12960_/A _12393_/A _15127_/S vssd1 vssd1 vccd1 vccd1 _09489_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11014__A _11295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ _09701_/A _11438_/X _11449_/X _09841_/A _18833_/Q vssd1 vssd1 vccd1 vccd1
+ _11450_/X sky130_fd_sc_hd__a32o_1
XFILLER_149_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10401_ _19244_/Q _19739_/Q _10447_/S vssd1 vssd1 vccd1 vccd1 _10401_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11381_ _11425_/A _11381_/B vssd1 vssd1 vccd1 vccd1 _11381_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10835__S1 _10820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16016__S _16020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10853__A _11015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _13120_/A vssd1 vssd1 vccd1 vccd1 _13120_/X sky130_fd_sc_hd__buf_2
X_10332_ _19677_/Q _19443_/Q _18508_/Q _19773_/Q _10005_/A _10283_/X vssd1 vssd1 vccd1
+ vccd1 _10332_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13051_ _18755_/Q _11670_/A _11703_/A _18461_/Q _11791_/A vssd1 vssd1 vccd1 vccd1
+ _13051_/X sky130_fd_sc_hd__a221o_1
XFILLER_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13154__A2 _11857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10263_ _10064_/X _10262_/X _09980_/X vssd1 vssd1 vccd1 vccd1 _10263_/X sky130_fd_sc_hd__o21a_1
XANTENNA__17636__A _17717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12002_ _12279_/C vssd1 vssd1 vccd1 vccd1 _12393_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_79_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09853__S _11534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_A io_ibus_inst[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _10194_/A _10194_/B _10194_/C vssd1 vssd1 vccd1 vccd1 _10194_/X sky130_fd_sc_hd__or3_2
XFILLER_87_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16810_ _16821_/A vssd1 vssd1 vccd1 vccd1 _16819_/S sky130_fd_sc_hd__buf_6
XFILLER_120_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17790_ _17790_/A vssd1 vssd1 vccd1 vccd1 _19773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16741_ _19341_/Q _13826_/X _16747_/S vssd1 vssd1 vccd1 vccd1 _16742_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_163_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _18956_/CLK sky130_fd_sc_hd__clkbuf_16
X_13953_ _14745_/A vssd1 vssd1 vccd1 vccd1 _14094_/A sky130_fd_sc_hd__buf_2
XFILLER_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14995__A _15368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10676__B1 _09686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12904_ _14789_/A vssd1 vssd1 vccd1 vccd1 _12904_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19460_ _19950_/CLK _19460_/D vssd1 vssd1 vccd1 vccd1 _19460_/Q sky130_fd_sc_hd__dfxtp_1
X_16672_ _16374_/X _19311_/Q _16674_/S vssd1 vssd1 vccd1 vccd1 _16673_/A sky130_fd_sc_hd__mux2_1
X_13884_ _16836_/A vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18411_ _18411_/A vssd1 vssd1 vccd1 vccd1 _20034_/D sky130_fd_sc_hd__clkbuf_1
X_15623_ _15623_/A vssd1 vssd1 vccd1 vccd1 _18892_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _12833_/A _12835_/B vssd1 vssd1 vccd1 vccd1 _12836_/A sky130_fd_sc_hd__and2b_4
X_19391_ _19979_/CLK _19391_/D vssd1 vssd1 vccd1 vccd1 _19391_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12417__A1 _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _17723_/X _20004_/Q _18346_/S vssd1 vssd1 vccd1 vccd1 _18343_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_178_clock _18998_/CLK vssd1 vssd1 vccd1 vccd1 _19488_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15211_/X _12807_/B _15212_/X _15553_/X vssd1 vssd1 vccd1 vccd1 _15554_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12766_/A vssd1 vssd1 vccd1 vccd1 _12766_/Y sky130_fd_sc_hd__inv_6
XANTENNA__13090__A1 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14505_ _14514_/A _14510_/C vssd1 vssd1 vccd1 vccd1 _14505_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18273_ _18273_/A vssd1 vssd1 vccd1 vccd1 _19973_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_182_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ _11730_/A vssd1 vssd1 vccd1 vccd1 _11717_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12697_ _12693_/A _12696_/X _12697_/S vssd1 vssd1 vccd1 vccd1 _12697_/X sky130_fd_sc_hd__mux2_1
X_15485_ _15082_/A _15487_/B _15081_/X _15484_/X vssd1 vssd1 vccd1 vccd1 _15485_/X
+ sky130_fd_sc_hd__o211a_1
X_17224_ _17115_/X _19532_/Q _17232_/S vssd1 vssd1 vccd1 vccd1 _17225_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11648_ _11648_/A _11648_/B _11648_/C vssd1 vssd1 vccd1 vccd1 _11648_/X sky130_fd_sc_hd__or3_1
X_14436_ _18706_/Q _14439_/C _14427_/X vssd1 vssd1 vccd1 vccd1 _14436_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_101_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _20030_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput12 io_dbus_rdata[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_2
Xinput23 io_dbus_rdata[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_4
Xinput34 io_ibus_inst[0] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_2
Xinput45 io_ibus_inst[1] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17155_ _17154_/X _19507_/Q _17161_/S vssd1 vssd1 vccd1 vccd1 _17156_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10826__S1 _10820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10763__A _10824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11579_ _11655_/A _11657_/A _11530_/X _11529_/A vssd1 vssd1 vccd1 vccd1 _11579_/Y
+ sky130_fd_sc_hd__o211ai_1
X_14367_ _14371_/B _14365_/C _14366_/X vssd1 vssd1 vccd1 vccd1 _14367_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput56 io_ibus_inst[2] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_8
Xinput67 io_irq_motor_irq vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
X_16106_ _16106_/A vssd1 vssd1 vccd1 vccd1 _19075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13318_ _13340_/A vssd1 vssd1 vccd1 vccd1 _13318_/X sky130_fd_sc_hd__buf_2
XANTENNA__09329__A _18940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17086_ _17086_/A vssd1 vssd1 vccd1 vccd1 _19481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14298_ _14319_/A _14306_/D vssd1 vssd1 vccd1 vccd1 _14298_/Y sky130_fd_sc_hd__nor2_1
X_16037_ _16037_/A vssd1 vssd1 vccd1 vccd1 _19047_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_116_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _20005_/CLK sky130_fd_sc_hd__clkbuf_16
X_13249_ _17049_/A vssd1 vssd1 vccd1 vccd1 _17691_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18141__S _18147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11251__S1 _10983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17988_ _17988_/A vssd1 vssd1 vccd1 vccd1 _19861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19727_ _20015_/CLK _19727_/D vssd1 vssd1 vccd1 vccd1 _19727_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12656__A1 _18542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16939_ _16939_/A vssd1 vssd1 vccd1 vccd1 _19428_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16596__S _16602_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19658_ _19755_/CLK _19658_/D vssd1 vssd1 vccd1 vccd1 _19658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10762__S0 _10872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09411_ _18711_/Q vssd1 vssd1 vccd1 vccd1 _09411_/Y sky130_fd_sc_hd__inv_2
X_18609_ _19941_/CLK _18609_/D vssd1 vssd1 vccd1 vccd1 _18609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19589_ _20007_/CLK _19589_/D vssd1 vssd1 vccd1 vccd1 _19589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09342_ _18824_/Q _09342_/B _09341_/X vssd1 vssd1 vccd1 vccd1 _09342_/X sky130_fd_sc_hd__or3b_2
XFILLER_80_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09273_ _09273_/A _09276_/C vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__or2_2
XANTENNA__18316__S _18324_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13908__A1 _18547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14581__A1 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14333__A1 _14336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 _20036_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10658__B1 _10836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__A _19526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10950_ _10943_/X _10945_/X _10947_/X _10949_/X _09804_/A vssd1 vssd1 vccd1 vccd1
+ _10950_/X sky130_fd_sc_hd__a221o_1
XFILLER_44_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10753__S0 _09725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19836_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ _10492_/A vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09702__A _09702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10881_ _19923_/Q _19537_/Q _19987_/Q _19106_/Q _10704_/A _10710_/A vssd1 vssd1 vccd1
+ vccd1 _10882_/B sky130_fd_sc_hd__mux4_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12620_ _12598_/A _12598_/B _12619_/X vssd1 vssd1 vccd1 vccd1 _12621_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__10505__S0 _09653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12551_ _12551_/A vssd1 vssd1 vccd1 vccd1 _12551_/Y sky130_fd_sc_hd__inv_6
XFILLER_157_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12280__C1 _12722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18226__S _18230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ _11502_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11502_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12482_ _12452_/A _12483_/C _18774_/Q vssd1 vssd1 vccd1 vccd1 _12482_/Y sky130_fd_sc_hd__a21oi_1
X_15270_ _15270_/A _15270_/B vssd1 vssd1 vccd1 vccd1 _15270_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11433_ _11401_/A _11432_/X _11181_/A vssd1 vssd1 vccd1 vccd1 _11433_/X sky130_fd_sc_hd__o21a_1
X_14221_ _18934_/Q _18932_/Q _18931_/Q _14220_/X vssd1 vssd1 vccd1 vccd1 _14222_/D
+ sky130_fd_sc_hd__or4b_1
XANTENNA__13375__A2 _13269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10583__A _18850_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14055__A _14245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11386__B2 _12934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _20018_/CLK sky130_fd_sc_hd__clkbuf_16
X_14152_ _14153_/B _14153_/C _18623_/Q vssd1 vssd1 vccd1 vccd1 _14154_/B sky130_fd_sc_hd__a21oi_1
XFILLER_98_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11364_ _11292_/X _12826_/B _11452_/A _12825_/B vssd1 vssd1 vccd1 vccd1 _11608_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_153_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10315_ _10355_/A _10314_/X _10462_/A vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13103_ _18463_/Q _11740_/X _12881_/A _18687_/Q _13102_/X vssd1 vssd1 vccd1 vccd1
+ _13103_/X sky130_fd_sc_hd__a221o_1
XANTENNA__13127__A2 _13070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14083_ _18603_/Q _14080_/B _14082_/Y vssd1 vssd1 vccd1 vccd1 _18603_/D sky130_fd_sc_hd__o21a_1
X_18960_ _18960_/CLK _18960_/D vssd1 vssd1 vccd1 vccd1 _18960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11295_ _19355_/Q _19690_/Q _11295_/S vssd1 vssd1 vccd1 vccd1 _11296_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ _19827_/Q _17033_/X _17915_/S vssd1 vssd1 vccd1 vccd1 _17912_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _18588_/Q _11851_/A _11855_/B _18720_/Q vssd1 vssd1 vccd1 vccd1 _13034_/X
+ sky130_fd_sc_hd__a22o_1
X_10246_ _10246_/A _10246_/B vssd1 vssd1 vccd1 vccd1 _11640_/B sky130_fd_sc_hd__and2_1
X_18891_ _18923_/CLK _18891_/D vssd1 vssd1 vccd1 vccd1 _18891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output153_A _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_129_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _20023_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17274__A0 _17189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__B2 _18757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17842_ _17842_/A vssd1 vssd1 vccd1 vccd1 _19796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10177_ _15974_/B _12860_/C vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12303__A _12340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15824__A1 _18970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10992__S0 _11048_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15824__B2 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17773_ _17795_/A vssd1 vssd1 vccd1 vccd1 _17782_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14985_ _14923_/X _14982_/X _14984_/X vssd1 vssd1 vccd1 vccd1 _14985_/X sky130_fd_sc_hd__o21a_1
X_19512_ _19999_/CLK _19512_/D vssd1 vssd1 vccd1 vccd1 _19512_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13833__S _13836_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16724_ _16724_/A vssd1 vssd1 vccd1 vccd1 _19333_/D sky130_fd_sc_hd__clkbuf_1
X_13936_ _18553_/Q _13936_/B _13936_/C vssd1 vssd1 vccd1 vccd1 _13937_/C sky130_fd_sc_hd__and3_1
XFILLER_35_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10744__S0 _10750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19443_ _19644_/CLK _19443_/D vssd1 vssd1 vccd1 vccd1 _19443_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09612__A _09612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16655_ _16348_/X _19303_/Q _16663_/S vssd1 vssd1 vccd1 vccd1 _16656_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13867_ _15807_/A vssd1 vssd1 vccd1 vccd1 _17203_/A sky130_fd_sc_hd__buf_4
XFILLER_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15606_ _15606_/A vssd1 vssd1 vccd1 vccd1 _18884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19374_ _19644_/CLK _19374_/D vssd1 vssd1 vccd1 vccd1 _19374_/Q sky130_fd_sc_hd__dfxtp_1
X_12818_ _12799_/A _12799_/B _18788_/Q vssd1 vssd1 vccd1 vccd1 _12818_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13063__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16586_ _16586_/A vssd1 vssd1 vccd1 vccd1 _19272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13798_ _18498_/Q _13797_/X _13804_/S vssd1 vssd1 vccd1 vccd1 _13799_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13063__B2 _12874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18325_ _18325_/A vssd1 vssd1 vccd1 vccd1 _19996_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ _18862_/Q _15457_/X _15536_/X vssd1 vssd1 vccd1 vccd1 _18862_/D sky130_fd_sc_hd__o21a_1
XFILLER_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12750_/B _12750_/C _18785_/Q vssd1 vssd1 vccd1 vccd1 _12749_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17040__S _17040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18256_ _18256_/A vssd1 vssd1 vccd1 vccd1 _19965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15468_ _12621_/X _15458_/X _15467_/X _15454_/X vssd1 vssd1 vccd1 vccd1 _15468_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17207_ _17207_/A vssd1 vssd1 vccd1 vccd1 _19525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14419_ _18701_/Q _14422_/C _14419_/C vssd1 vssd1 vccd1 vccd1 _14420_/C sky130_fd_sc_hd__and3_1
X_18187_ _17707_/X _19935_/Q _18191_/S vssd1 vssd1 vccd1 vccd1 _18188_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15399_ _15399_/A _15399_/B _15399_/C vssd1 vssd1 vccd1 vccd1 _15399_/X sky130_fd_sc_hd__and3_1
XFILLER_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17138_ _17675_/A vssd1 vssd1 vccd1 vccd1 _17138_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11472__S1 _10596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17069_ _19476_/Q _17068_/X _17072_/S vssd1 vssd1 vccd1 vccd1 _17070_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09960_ _09953_/Y _09955_/Y _09957_/Y _09959_/Y _09807_/X vssd1 vssd1 vccd1 vccd1
+ _09960_/X sky130_fd_sc_hd__o221a_1
XFILLER_104_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12326__A0 _15938_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09891_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09891_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11224__S1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10888__B1 _10719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15276__C1 _15275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13743__S _16066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17215__S _17221_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09522__A _09522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10668__A _10668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09325_ _18984_/Q _12913_/A _09697_/B _09696_/B vssd1 vssd1 vccd1 vccd1 _09909_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12883__A _13164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11160__S0 _09721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__S _09668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09256_ _09256_/A _11920_/B _11920_/C vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__or3_2
XANTENNA__17885__S _17893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14554__A1 _13531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09187_ _11919_/A _09313_/A _09189_/A _14755_/A vssd1 vssd1 vccd1 vccd1 _09188_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_147_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15503__B1 _15502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10100_ _10007_/A _10099_/X _09798_/A vssd1 vssd1 vccd1 vccd1 _10100_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11080_ _11067_/Y _11072_/Y _11075_/Y _11079_/Y _09549_/A vssd1 vssd1 vccd1 vccd1
+ _11081_/A sky130_fd_sc_hd__o221a_1
XANTENNA__11215__S1 _11065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_130_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10031_ _18449_/Q _19478_/Q _19515_/Q _19089_/Q _10275_/A _09747_/A vssd1 vssd1 vccd1
+ vccd1 _10031_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14770_ _14771_/B vssd1 vssd1 vccd1 vccd1 _15747_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11982_ _18978_/Q vssd1 vssd1 vccd1 vccd1 _11982_/X sky130_fd_sc_hd__buf_4
XFILLER_57_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11681__B _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ _18481_/Q _13526_/A _13716_/Y _13720_/X vssd1 vssd1 vccd1 vccd1 _18481_/D
+ sky130_fd_sc_hd__o22a_1
X_10933_ _20018_/Q _19856_/Q _19265_/Q _19035_/Q _10776_/A _10709_/A vssd1 vssd1 vccd1
+ vccd1 _10934_/B sky130_fd_sc_hd__mux4_1
XFILLER_95_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16964__S _16964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16440_ _19208_/Q _13810_/X _16446_/S vssd1 vssd1 vccd1 vccd1 _16441_/A sky130_fd_sc_hd__mux2_1
X_10864_ _19139_/Q _19400_/Q _19299_/Q _19634_/Q _10953_/S _10793_/A vssd1 vssd1 vccd1
+ vccd1 _10865_/B sky130_fd_sc_hd__mux4_1
XFILLER_32_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13652_ _18472_/Q _13517_/X _13649_/Y _13651_/X vssd1 vssd1 vccd1 vccd1 _18472_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14992__B _14996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _18476_/Q _12556_/X _12557_/X vssd1 vssd1 vccd1 vccd1 _12603_/Y sky130_fd_sc_hd__o21ai_1
X_16371_ _17707_/A vssd1 vssd1 vccd1 vccd1 _16371_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _10858_/A _10795_/B vssd1 vssd1 vccd1 vccd1 _10795_/Y sky130_fd_sc_hd__nor2_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13583_ _13579_/X _13582_/Y _13583_/S vssd1 vssd1 vccd1 vccd1 _13583_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18110_ _18110_/A vssd1 vssd1 vccd1 vccd1 _19904_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_55_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15322_ _15305_/X _15316_/Y _15321_/Y vssd1 vssd1 vccd1 vccd1 _15323_/C sky130_fd_sc_hd__a21oi_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _19942_/CLK _19090_/D vssd1 vssd1 vccd1 vccd1 _19090_/Q sky130_fd_sc_hd__dfxtp_1
X_12534_ _18537_/Q _12415_/X _12528_/X _12533_/Y vssd1 vssd1 vccd1 vccd1 _12534_/X
+ sky130_fd_sc_hd__o22a_4
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18041_ hold8/X _19884_/Q _18044_/S vssd1 vssd1 vccd1 vccd1 _18042_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14545__A1 _18754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15253_ _15209_/X _15250_/Y _15252_/X _15216_/X vssd1 vssd1 vccd1 vccd1 _15256_/B
+ sky130_fd_sc_hd__a211o_1
X_12465_ _12465_/A _12495_/A vssd1 vssd1 vccd1 vccd1 _12466_/A sky130_fd_sc_hd__or2_1
X_14204_ _18640_/Q _14207_/C _14203_/X vssd1 vssd1 vccd1 vccd1 _14204_/Y sky130_fd_sc_hd__a21oi_1
X_11416_ _19320_/Q _19591_/Q _19815_/Q _19559_/Q _10980_/A _10972_/A vssd1 vssd1 vccd1
+ vccd1 _11416_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12396_ _16066_/S vssd1 vssd1 vccd1 vccd1 _13648_/A sky130_fd_sc_hd__clkbuf_4
X_15184_ _15100_/A _15043_/X _14984_/A vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__o21ai_1
XFILLER_153_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17096__A _17203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11347_ _11340_/Y _11342_/Y _11344_/Y _11346_/Y _09816_/A vssd1 vssd1 vccd1 vccd1
+ _11347_/X sky130_fd_sc_hd__o221a_2
X_14135_ _18618_/Q _18617_/Q _18616_/Q _14135_/D vssd1 vssd1 vccd1 vccd1 _14144_/D
+ sky130_fd_sc_hd__and4_1
X_19992_ _19993_/CLK _19992_/D vssd1 vssd1 vccd1 vccd1 _19992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16204__S _16206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09607__A _09607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14066_ _14090_/A _14070_/C vssd1 vssd1 vccd1 vccd1 _14066_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_output78_A _12443_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18943_ _18974_/CLK _18943_/D vssd1 vssd1 vccd1 vccd1 _18943_/Q sky130_fd_sc_hd__dfxtp_1
X_11278_ _11278_/A _11278_/B vssd1 vssd1 vccd1 vccd1 _11278_/X sky130_fd_sc_hd__or2_1
XANTENNA__10760__B _12843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11348__S _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10229_ _09798_/A _10221_/X _10225_/Y _10228_/Y _09807_/A vssd1 vssd1 vccd1 vccd1
+ _10229_/X sky130_fd_sc_hd__o221a_1
X_13017_ _18870_/Q vssd1 vssd1 vccd1 vccd1 _13554_/A sky130_fd_sc_hd__clkbuf_2
X_18874_ _18911_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 _18874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17825_ _17825_/A vssd1 vssd1 vccd1 vccd1 _19788_/D sky130_fd_sc_hd__clkbuf_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__14659__S _14667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17756_ _17659_/X _19758_/Q _17760_/S vssd1 vssd1 vccd1 vccd1 _17757_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14968_ _15553_/B _14973_/A vssd1 vssd1 vccd1 vccd1 _14970_/C sky130_fd_sc_hd__and2_1
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16707_ _16707_/A vssd1 vssd1 vccd1 vccd1 _19325_/D sky130_fd_sc_hd__clkbuf_1
X_13919_ _18605_/Q _18604_/Q _18606_/Q _14081_/A vssd1 vssd1 vccd1 vccd1 _14089_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17687_ _17687_/A vssd1 vssd1 vccd1 vccd1 _19734_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10488__A _18852_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14899_ _15078_/B _12760_/A _14915_/S vssd1 vssd1 vccd1 vccd1 _14899_/X sky130_fd_sc_hd__mux2_1
X_19426_ _19758_/CLK _19426_/D vssd1 vssd1 vccd1 vccd1 _19426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16638_ _16638_/A vssd1 vssd1 vccd1 vccd1 _19295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19357_ _19758_/CLK _19357_/D vssd1 vssd1 vccd1 vccd1 _19357_/Q sky130_fd_sc_hd__dfxtp_1
X_16569_ _19265_/Q _13787_/X _16569_/S vssd1 vssd1 vccd1 vccd1 _16570_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15981__B1 _15928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16175__A _16221_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18308_ _18308_/A vssd1 vssd1 vccd1 vccd1 _19988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09488__S _15127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19288_ _19389_/CLK _19288_/D vssd1 vssd1 vccd1 vccd1 _19288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18239_ _19958_/Q _17678_/A _18241_/S vssd1 vssd1 vccd1 vccd1 _18240_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12011__A2 _11994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11445__S1 _11107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09517__A _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09943_ _20037_/Q _19875_/Q _19284_/Q _19054_/Q _09939_/X _09940_/A vssd1 vssd1 vccd1
+ vccd1 _09943_/X sky130_fd_sc_hd__mux4_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11258__S _11258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _09874_/A vssd1 vssd1 vccd1 vccd1 _09875_/A sky130_fd_sc_hd__buf_4
XFILLER_135_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09951__S _10094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16069__B _16069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16784__S _16786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09402__D _09402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11038__B1 _09774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14775__A1 _12866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10941__A1_N _18842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09308_ _12290_/B _12831_/A vssd1 vssd1 vccd1 vccd1 _14821_/A sky130_fd_sc_hd__nand2_2
XFILLER_70_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10580_ _10149_/A _10578_/X _10579_/X vssd1 vssd1 vccd1 vccd1 _10580_/X sky130_fd_sc_hd__o21a_1
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_clock clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__14317__B _18670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09239_ _18992_/Q _18967_/Q _18966_/Q _18965_/Q vssd1 vssd1 vccd1 vccd1 _09247_/C
+ sky130_fd_sc_hd__or4bb_1
XANTENNA__11022__A _11022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10326__A1_N _18855_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ _12279_/A _12393_/B _12393_/C _12246_/X vssd1 vssd1 vccd1 vccd1 _12250_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_108_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11201_ _11335_/A vssd1 vssd1 vccd1 vccd1 _11425_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_123_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11210__B1 _11058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12181_ _12217_/A _14906_/A vssd1 vssd1 vccd1 vccd1 _12182_/B sky130_fd_sc_hd__nor2_1
XFILLER_150_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11132_ _11137_/A _11129_/X _11131_/X _11058_/X vssd1 vssd1 vccd1 vccd1 _11133_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11063_ _11410_/S vssd1 vssd1 vccd1 vccd1 _11063_/X sky130_fd_sc_hd__buf_4
X_15940_ _15940_/A _15955_/A _15940_/C vssd1 vssd1 vccd1 vccd1 _15940_/X sky130_fd_sc_hd__and3_1
XFILLER_135_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10014_ _20034_/Q _19872_/Q _19281_/Q _19051_/Q _10275_/A _10082_/A vssd1 vssd1 vccd1
+ vccd1 _10014_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15871_ _15871_/A _16843_/B vssd1 vssd1 vccd1 vccd1 _18984_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17610_ _17610_/A vssd1 vssd1 vccd1 vccd1 _19707_/D sky130_fd_sc_hd__clkbuf_1
X_14822_ _15368_/A _14822_/B _14822_/C _14822_/D vssd1 vssd1 vccd1 vccd1 _15004_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_64_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18590_ _18724_/CLK _18590_/D vssd1 vssd1 vccd1 vccd1 _18590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17541_ _17541_/A vssd1 vssd1 vccd1 vccd1 _19676_/D sky130_fd_sc_hd__clkbuf_1
X_14753_ _09280_/Y _11663_/A _11975_/A _12859_/A vssd1 vssd1 vccd1 vccd1 _14753_/X
+ sky130_fd_sc_hd__a211o_1
X_11965_ _11945_/A _11943_/X _11945_/Y vssd1 vssd1 vccd1 vccd1 _12078_/B sky130_fd_sc_hd__o21a_1
XANTENNA_output116_A _12847_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__S0 _10980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13704_ _11813_/X _13702_/X _13703_/Y _11831_/X _19019_/Q vssd1 vssd1 vccd1 vccd1
+ _13704_/X sky130_fd_sc_hd__a32o_2
X_17472_ _17483_/A vssd1 vssd1 vccd1 vccd1 _17481_/S sky130_fd_sc_hd__buf_4
X_10916_ _15934_/B _12837_/B vssd1 vssd1 vccd1 vccd1 _10918_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14684_ _14684_/A vssd1 vssd1 vccd1 vccd1 _18794_/D sky130_fd_sc_hd__clkbuf_1
X_11896_ _19018_/Q _11896_/B vssd1 vssd1 vccd1 vccd1 _11896_/X sky130_fd_sc_hd__or2_1
X_19211_ _19771_/CLK _19211_/D vssd1 vssd1 vccd1 vccd1 _19211_/Q sky130_fd_sc_hd__dfxtp_1
X_16423_ _16423_/A vssd1 vssd1 vccd1 vccd1 _19200_/D sky130_fd_sc_hd__clkbuf_1
X_13635_ _13635_/A vssd1 vssd1 vccd1 vccd1 _18469_/D sky130_fd_sc_hd__clkbuf_1
X_10847_ _19203_/Q _19794_/Q _19956_/Q _19171_/Q _10953_/S _10793_/A vssd1 vssd1 vccd1
+ vccd1 _10848_/B sky130_fd_sc_hd__mux4_1
X_19142_ _19637_/CLK _19142_/D vssd1 vssd1 vccd1 vccd1 _19142_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12777__B1 _12864_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16354_ _16354_/A vssd1 vssd1 vccd1 vccd1 _19176_/D sky130_fd_sc_hd__clkbuf_1
X_13566_ _13580_/C _13565_/Y _12557_/A vssd1 vssd1 vccd1 vccd1 _13566_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10778_ _10886_/A _10777_/X _10712_/A vssd1 vssd1 vccd1 vccd1 _10778_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14227__B _14227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15305_ _15305_/A vssd1 vssd1 vccd1 vccd1 _15305_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19073_ _19824_/CLK _19073_/D vssd1 vssd1 vccd1 vccd1 _19073_/Q sky130_fd_sc_hd__dfxtp_1
X_12517_ _15958_/C _18916_/Q _12517_/S vssd1 vssd1 vccd1 vccd1 _14886_/A sky130_fd_sc_hd__mux2_4
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16285_ _13406_/X _19154_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _16286_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18414__S _18418_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13497_ _12875_/X _13495_/X _13496_/X vssd1 vssd1 vccd1 vccd1 _13497_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_145_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18024_ _19878_/Q _17093_/X _18024_/S vssd1 vssd1 vccd1 vccd1 _18025_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15236_ _15236_/A _15236_/B _15236_/C vssd1 vssd1 vccd1 vccd1 _15236_/X sky130_fd_sc_hd__and3_1
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12448_ _12443_/A _12447_/X _12448_/S vssd1 vssd1 vccd1 vccd1 _12448_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15167_ _15165_/X _15166_/X _15190_/S vssd1 vssd1 vccd1 vccd1 _15167_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13741__A2 _13472_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12379_ _12537_/A _12843_/A _12318_/B vssd1 vssd1 vccd1 vccd1 _12379_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14118_ _18733_/Q _18735_/Q _18734_/Q _14496_/A vssd1 vssd1 vccd1 vccd1 _14504_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_141_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19975_ _19975_/CLK _19975_/D vssd1 vssd1 vccd1 vccd1 _19975_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10490__B _12850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15098_ _14978_/X _15096_/X _15097_/X vssd1 vssd1 vccd1 vccd1 _15098_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14049_ _14051_/B _14051_/C _14048_/Y vssd1 vssd1 vccd1 vccd1 _18592_/D sky130_fd_sc_hd__o21a_1
X_18926_ _18926_/CLK _18926_/D vssd1 vssd1 vccd1 vccd1 _18926_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11504__A1 _10858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12701__B1 _12170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18857_ _19025_/CLK _18857_/D vssd1 vssd1 vccd1 vccd1 _18857_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_95_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09590_ _11468_/S vssd1 vssd1 vccd1 vccd1 _10724_/S sky130_fd_sc_hd__clkbuf_4
X_17808_ _17735_/X _19782_/Q _17808_/S vssd1 vssd1 vccd1 vccd1 _17809_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18788_ _18789_/CLK _18788_/D vssd1 vssd1 vccd1 vccd1 _18788_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17739_ _17795_/A vssd1 vssd1 vccd1 vccd1 _17808_/S sky130_fd_sc_hd__buf_6
XANTENNA__11268__B1 _09546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11107__A _11107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10011__A _10011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13009__B2 _12165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19409_ _19965_/CLK _19409_/D vssd1 vssd1 vccd1 vccd1 _19409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16109__S _16111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13322__A _17062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__S1 _09642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12864__C _12864_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15706__B1 _14529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18324__S _18324_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17459__A0 _17144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13193__B1 _11852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11777__A _15760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15485__A2 _15487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09926_ _09933_/A _09925_/X _09690_/A vssd1 vssd1 vccd1 vccd1 _09926_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09857_ _09851_/X _09854_/X _09856_/X _11547_/A _09568_/X vssd1 vssd1 vccd1 vccd1
+ _09862_/B sky130_fd_sc_hd__o221a_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _09788_/A vssd1 vssd1 vccd1 vccd1 _09789_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17403__S _17409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11017__A _11017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _18748_/Q _13910_/A _14670_/S vssd1 vssd1 vccd1 vccd1 _11750_/X sky130_fd_sc_hd__and3_1
XFILLER_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10482__A1 _10001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ _15947_/C _12844_/A vssd1 vssd1 vccd1 vccd1 _11599_/A sky130_fd_sc_hd__or2_1
XFILLER_14_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11869_/A _11688_/A vssd1 vssd1 vccd1 vccd1 _11682_/A sky130_fd_sc_hd__nor2_2
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14328__A _14479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12759__A0 _15978_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13420_ _13307_/X _13411_/Y _13412_/Y _13419_/Y _09532_/A vssd1 vssd1 vccd1 vccd1
+ _13420_/X sky130_fd_sc_hd__a221o_2
X_10632_ _19929_/Q _19543_/Q _19993_/Q _19112_/Q _10637_/S _10010_/A vssd1 vssd1 vccd1
+ vccd1 _10633_/B sky130_fd_sc_hd__mux4_1
XFILLER_22_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ _10572_/A _10563_/B vssd1 vssd1 vccd1 vccd1 _10563_/Y sky130_fd_sc_hd__nor2_1
X_13351_ input16/X _13340_/X _13319_/X vssd1 vssd1 vccd1 vccd1 _13351_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _18529_/Q vssd1 vssd1 vccd1 vccd1 _12340_/A sky130_fd_sc_hd__buf_2
X_16070_ _19061_/Q _16069_/Y _16073_/S vssd1 vssd1 vccd1 vccd1 _16071_/A sky130_fd_sc_hd__mux2_1
X_10494_ _10448_/A _10493_/X _09987_/A vssd1 vssd1 vccd1 vccd1 _10494_/X sky130_fd_sc_hd__a21o_1
X_13282_ _17055_/A vssd1 vssd1 vccd1 vccd1 _17697_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15173__B2 _12124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09927__A1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15021_ _15018_/X _15019_/X _15114_/S vssd1 vssd1 vccd1 vccd1 _15021_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12233_ _12228_/X _12229_/Y _12231_/X _12232_/Y vssd1 vssd1 vccd1 vccd1 _12233_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_136_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18111__A1 _11898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12164_ _18762_/Q _16072_/A vssd1 vssd1 vccd1 vccd1 _12164_/X sky130_fd_sc_hd__and2_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16689__S _16689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11115_ _11145_/A _11115_/B vssd1 vssd1 vccd1 vccd1 _11115_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16972_ _16972_/A vssd1 vssd1 vccd1 vccd1 _19443_/D sky130_fd_sc_hd__clkbuf_1
X_19760_ _20018_/CLK _19760_/D vssd1 vssd1 vccd1 vccd1 _19760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12095_ _18522_/Q _12583_/A vssd1 vssd1 vccd1 vccd1 _12113_/A sky130_fd_sc_hd__or2_1
XFILLER_150_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18711_ _18993_/CLK _18711_/D vssd1 vssd1 vccd1 vccd1 _18711_/Q sky130_fd_sc_hd__dfxtp_2
X_15923_ _15940_/A _15955_/A _15923_/C vssd1 vssd1 vccd1 vccd1 _15923_/X sky130_fd_sc_hd__and3_1
X_11046_ _19662_/Q _19428_/Q _18493_/Q _19758_/Q _10977_/S _11045_/X vssd1 vssd1 vccd1
+ vccd1 _11047_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09786__S0 _11553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19691_ _19755_/CLK _19691_/D vssd1 vssd1 vccd1 vccd1 _19691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18642_ _18655_/CLK _18642_/D vssd1 vssd1 vccd1 vccd1 _18642_/Q sky130_fd_sc_hd__dfxtp_1
X_15854_ _15861_/A _17206_/B vssd1 vssd1 vccd1 vccd1 _15855_/A sky130_fd_sc_hd__and2_1
XFILLER_49_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14805_ _14805_/A _14812_/B vssd1 vssd1 vccd1 vccd1 _14807_/C sky130_fd_sc_hd__nor2_1
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18573_ _20005_/CLK _18573_/D vssd1 vssd1 vccd1 vccd1 _18573_/Q sky130_fd_sc_hd__dfxtp_1
X_15785_ input34/X vssd1 vssd1 vccd1 vccd1 _15785_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12030__B _14865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ _12997_/A vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__buf_2
XFILLER_80_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11345__S0 _11230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16189__A0 _13238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17524_ _19668_/Q vssd1 vssd1 vccd1 vccd1 _17525_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__17313__S _17315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12998__B1 _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14736_ _18818_/Q _13727_/X _14738_/S vssd1 vssd1 vccd1 vccd1 _14737_/A sky130_fd_sc_hd__mux2_1
X_11948_ _11948_/A _11948_/B vssd1 vssd1 vccd1 vccd1 _14815_/B sky130_fd_sc_hd__or2_1
XFILLER_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _17138_/X _19635_/Q _17459_/S vssd1 vssd1 vccd1 vccd1 _17456_/A sky130_fd_sc_hd__mux2_1
X_14667_ _18788_/Q _13750_/B _14667_/S vssd1 vssd1 vccd1 vccd1 _14668_/B sky130_fd_sc_hd__mux2_1
X_11879_ _11731_/X _11877_/X _11878_/Y _11723_/X _19017_/Q vssd1 vssd1 vccd1 vccd1
+ _11879_/X sky130_fd_sc_hd__a32o_4
X_16406_ _16406_/A vssd1 vssd1 vccd1 vccd1 _19192_/D sky130_fd_sc_hd__clkbuf_1
X_13618_ _13618_/A vssd1 vssd1 vccd1 vccd1 _18467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17386_ _17386_/A vssd1 vssd1 vccd1 vccd1 _19604_/D sky130_fd_sc_hd__clkbuf_1
X_14598_ _18768_/Q _11833_/D _14598_/S vssd1 vssd1 vccd1 vccd1 _14599_/B sky130_fd_sc_hd__mux2_1
XANTENNA__17689__A0 _17688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19125_ _20038_/CLK _19125_/D vssd1 vssd1 vccd1 vccd1 _19125_/Q sky130_fd_sc_hd__dfxtp_1
X_16337_ _16336_/X _19171_/Q _16346_/S vssd1 vssd1 vccd1 vccd1 _16338_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13549_ _18459_/Q _13548_/X _13575_/S vssd1 vssd1 vccd1 vccd1 _13550_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19056_ _19975_/CLK _19056_/D vssd1 vssd1 vccd1 vccd1 _19056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16268_ _16268_/A vssd1 vssd1 vccd1 vccd1 _19146_/D sky130_fd_sc_hd__clkbuf_1
X_18007_ _19870_/Q _17068_/X _18009_/S vssd1 vssd1 vccd1 vccd1 _18008_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17983__S _17987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15219_ _15219_/A _15219_/B vssd1 vssd1 vccd1 vccd1 _15219_/Y sky130_fd_sc_hd__nor2_1
X_16199_ _16199_/A vssd1 vssd1 vccd1 vccd1 _19116_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17284__A _17352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19958_ _19989_/CLK _19958_/D vssd1 vssd1 vccd1 vccd1 _19958_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13478__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_177_clock_A _18998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ _10572_/A vssd1 vssd1 vccd1 vccd1 _10172_/A sky130_fd_sc_hd__clkbuf_2
X_18909_ _18911_/CLK _18909_/D vssd1 vssd1 vccd1 vccd1 _18909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19889_ _19896_/CLK _19889_/D vssd1 vssd1 vccd1 vccd1 _19889_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16416__A1 _13774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09642_ _09642_/A vssd1 vssd1 vccd1 vccd1 _09851_/A sky130_fd_sc_hd__buf_2
XFILLER_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09573_ _10934_/A vssd1 vssd1 vccd1 vccd1 _11473_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09303__C1 _18827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12989__B1 _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09854__B1 _09933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10464__A1 _10411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11661__B1 _11657_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10311__S1 _10260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17893__S _17893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14902__A1 _12783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14314__C _14314_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16302__S _16314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09909_ _09909_/A _09909_/B _09909_/C vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__nand3_1
XANTENNA__09705__A _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12141__B2 _09261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20029_ _20031_/CLK _20029_/D vssd1 vssd1 vccd1 vccd1 _20029_/Q sky130_fd_sc_hd__dfxtp_1
X_12920_ _16993_/A _18352_/B vssd1 vssd1 vccd1 vccd1 _17098_/C sky130_fd_sc_hd__or2_1
XANTENNA__13227__A _13227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _12851_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12851_/Y sky130_fd_sc_hd__nor2_4
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15091__B1 _15457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17133__S _17145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _11860_/B _13519_/B _17096_/B vssd1 vssd1 vccd1 vccd1 _11802_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _12973_/B _18900_/Q _15578_/S vssd1 vssd1 vccd1 vccd1 _15571_/A sky130_fd_sc_hd__mux2_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11247__A3 _19165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12782_ _12781_/Y _18927_/Q _12782_/S vssd1 vssd1 vccd1 vccd1 _12783_/A sky130_fd_sc_hd__mux2_4
XANTENNA__17907__A1 _17026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11101__C1 _09817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14521_ _14521_/A vssd1 vssd1 vccd1 vccd1 _14526_/C sky130_fd_sc_hd__clkbuf_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _11824_/A vssd1 vssd1 vccd1 vccd1 _11733_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _17240_/A vssd1 vssd1 vccd1 vccd1 _19539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14452_/A _14452_/B _14452_/C vssd1 vssd1 vccd1 vccd1 _18716_/D sky130_fd_sc_hd__nor3_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11664_/A vssd1 vssd1 vccd1 vccd1 _15740_/A sky130_fd_sc_hd__buf_2
XFILLER_30_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15933__A3 _12239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13403_ _13307_/X _13393_/X _13394_/Y _13402_/Y _13460_/A vssd1 vssd1 vccd1 vccd1
+ _13403_/X sky130_fd_sc_hd__a221o_1
X_17171_ _17170_/X _19512_/Q _17177_/S vssd1 vssd1 vccd1 vccd1 _17172_/A sky130_fd_sc_hd__mux2_1
X_10615_ _18849_/Q _09538_/A _09547_/A _10614_/X vssd1 vssd1 vccd1 vccd1 _15949_/B
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__13897__A _14385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14383_ _18691_/Q _14391_/D vssd1 vssd1 vccd1 vccd1 _14385_/B sky130_fd_sc_hd__or2_1
XFILLER_155_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11595_ _11595_/A _11599_/A _11595_/C vssd1 vssd1 vccd1 vccd1 _11595_/X sky130_fd_sc_hd__and3_1
XANTENNA__10302__S1 _10260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16122_ _13283_/X _19083_/Q _16122_/S vssd1 vssd1 vccd1 vccd1 _16123_/A sky130_fd_sc_hd__mux2_1
X_13334_ _18604_/Q vssd1 vssd1 vccd1 vccd1 _14086_/B sky130_fd_sc_hd__clkbuf_2
X_10546_ _10542_/X _10544_/X _10545_/X _10553_/A _09563_/A vssd1 vssd1 vccd1 vccd1
+ _10551_/B sky130_fd_sc_hd__o221a_1
XFILLER_116_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_4_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_127_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16053_ _13463_/X _19055_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16054_/A sky130_fd_sc_hd__mux2_1
X_13265_ _13265_/A vssd1 vssd1 vccd1 vccd1 _18442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10477_ _10380_/A _10474_/X _10476_/X vssd1 vssd1 vccd1 vccd1 _10477_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15004_ _15004_/A _15004_/B _14955_/S vssd1 vssd1 vccd1 vccd1 _15413_/A sky130_fd_sc_hd__nor3b_1
XFILLER_108_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12216_ _12092_/A _12120_/X _12122_/B _12150_/A _12215_/D vssd1 vssd1 vccd1 vccd1
+ _12216_/X sky130_fd_sc_hd__o2111a_1
XFILLER_123_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13196_ _18564_/Q _13189_/X _13192_/X _13193_/X _13195_/X vssd1 vssd1 vccd1 vccd1
+ _13619_/B sky130_fd_sc_hd__a2111o_2
XANTENNA__13836__S _13836_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__A1 _09522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19812_ _19876_/CLK _19812_/D vssd1 vssd1 vccd1 vccd1 _19812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ _15923_/C _18903_/Q _12358_/S vssd1 vssd1 vccd1 vccd1 _14909_/A sky130_fd_sc_hd__mux2_2
XFILLER_2_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19743_ _20032_/CLK _19743_/D vssd1 vssd1 vccd1 vccd1 _19743_/Q sky130_fd_sc_hd__dfxtp_1
X_16955_ _16977_/A vssd1 vssd1 vccd1 vccd1 _16964_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12078_ _12078_/A _12078_/B _12078_/C _12078_/D vssd1 vssd1 vccd1 vccd1 _12209_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13137__A _17668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15906_ _15906_/A vssd1 vssd1 vccd1 vccd1 _18995_/D sky130_fd_sc_hd__clkbuf_1
X_11029_ _11032_/A _11028_/X _09791_/A vssd1 vssd1 vccd1 vccd1 _11029_/Y sky130_fd_sc_hd__o21ai_1
X_19674_ _19996_/CLK _19674_/D vssd1 vssd1 vccd1 vccd1 _19674_/Q sky130_fd_sc_hd__dfxtp_1
X_16886_ _16352_/X _19405_/Q _16892_/S vssd1 vssd1 vccd1 vccd1 _16887_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15837_ input38/X _15834_/X _15789_/X _15740_/A vssd1 vssd1 vccd1 vccd1 _15838_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_18625_ _18660_/CLK _18625_/D vssd1 vssd1 vccd1 vccd1 _18625_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14667__S _14667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18139__S _18147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15768_ _18953_/Q _15775_/B vssd1 vssd1 vccd1 vccd1 _15768_/X sky130_fd_sc_hd__or2_1
X_18556_ _19883_/CLK _18556_/D vssd1 vssd1 vccd1 vccd1 _18556_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14719_ _18810_/Q _13667_/X _14727_/S vssd1 vssd1 vccd1 vccd1 _14720_/A sky130_fd_sc_hd__mux2_1
X_17507_ _17507_/A vssd1 vssd1 vccd1 vccd1 _19659_/D sky130_fd_sc_hd__clkbuf_1
X_18487_ _19946_/CLK _18487_/D vssd1 vssd1 vccd1 vccd1 _18487_/Q sky130_fd_sc_hd__dfxtp_1
X_15699_ _18926_/Q _18547_/Q _15699_/S vssd1 vssd1 vccd1 vccd1 _15700_/A sky130_fd_sc_hd__mux2_1
X_17438_ _17438_/A vssd1 vssd1 vccd1 vccd1 _19627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13396__B1 _12944_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17369_ _17369_/A vssd1 vssd1 vccd1 vccd1 _19596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19108_ _19636_/CLK _19108_/D vssd1 vssd1 vccd1 vccd1 _19108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039_ _19636_/CLK _19039_/D vssd1 vssd1 vccd1 vccd1 _19039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput100 _12186_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[7] sky130_fd_sc_hd__buf_2
XANTENNA__09509__B _14766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput111 _12840_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[11] sky130_fd_sc_hd__buf_2
Xoutput122 _12853_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[21] sky130_fd_sc_hd__buf_2
Xoutput133 _12867_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[31] sky130_fd_sc_hd__buf_2
XFILLER_133_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput144 _12313_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[11] sky130_fd_sc_hd__buf_2
XFILLER_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput155 _12585_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[21] sky130_fd_sc_hd__buf_2
Xoutput166 _12821_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[31] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_opt_6_0_clock_A _18998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11557__S0 _11553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15860__A2 _15856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09625_ _10674_/A vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__buf_2
XFILLER_44_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ _19525_/Q vssd1 vssd1 vccd1 vccd1 _09557_/A sky130_fd_sc_hd__inv_2
XFILLER_102_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13623__A1 _13622_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09487_ _15945_/A vssd1 vssd1 vccd1 vccd1 _15127_/S sky130_fd_sc_hd__buf_4
XFILLER_62_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13387__A0 _13385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10400_ _10400_/A _10400_/B vssd1 vssd1 vccd1 vccd1 _10400_/X sky130_fd_sc_hd__and2_1
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11380_ _19193_/Q _19784_/Q _19946_/Q _19161_/Q _09586_/A _11208_/A vssd1 vssd1 vccd1
+ vccd1 _11381_/B sky130_fd_sc_hd__mux4_1
XFILLER_109_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ _10210_/A _10330_/X _10335_/A vssd1 vssd1 vccd1 vccd1 _10331_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10262_ _19343_/Q _19614_/Q _19838_/Q _19582_/Q _10059_/S _10261_/X vssd1 vssd1 vccd1
+ vccd1 _10262_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13050_ _18685_/Q _11819_/A _11671_/A _18750_/Q vssd1 vssd1 vccd1 vccd1 _13050_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12898__C1 _12897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ _12001_/A vssd1 vssd1 vccd1 vccd1 _12279_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10193_ _10369_/A _10189_/X _10191_/X _10192_/X vssd1 vssd1 vccd1 vccd1 _10194_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16967__S _16975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11548__S0 _11534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16740_ _16740_/A vssd1 vssd1 vccd1 vccd1 _19340_/D sky130_fd_sc_hd__clkbuf_1
X_13952_ _13956_/B _13956_/C _13951_/Y vssd1 vssd1 vccd1 vccd1 _18558_/D sky130_fd_sc_hd__o21a_1
XFILLER_143_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12903_ _18830_/Q vssd1 vssd1 vccd1 vccd1 _13092_/A sky130_fd_sc_hd__inv_2
X_16671_ _16671_/A vssd1 vssd1 vccd1 vccd1 _19310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11873__B1 _09405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13883_ _13900_/A vssd1 vssd1 vccd1 vccd1 _13883_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18410_ _17716_/X _20034_/Q _18418_/S vssd1 vssd1 vccd1 vccd1 _18411_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15622_ _13714_/B _18924_/Q _15622_/S vssd1 vssd1 vccd1 vccd1 _15623_/A sky130_fd_sc_hd__mux2_1
X_12834_ _12834_/A _12844_/B vssd1 vssd1 vccd1 vccd1 _12834_/Y sky130_fd_sc_hd__nor2_4
X_19390_ _19979_/CLK _19390_/D vssd1 vssd1 vccd1 vccd1 _19390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12417__A2 _12416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17798__S _17804_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18341_ _18341_/A vssd1 vssd1 vccd1 vccd1 _20003_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15553_/A _15553_/B vssd1 vssd1 vccd1 vccd1 _15553_/X sky130_fd_sc_hd__or2_1
X_12765_ _12765_/A _12765_/B vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__xnor2_4
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14504_/A vssd1 vssd1 vccd1 vccd1 _14510_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_125_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18272_ _19973_/Q _17726_/A _18274_/S vssd1 vssd1 vccd1 vccd1 _18273_/A sky130_fd_sc_hd__mux2_1
X_11716_ _11716_/A _18825_/Q vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__and2_2
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15553_/A _15487_/A vssd1 vssd1 vccd1 vccd1 _15484_/X sky130_fd_sc_hd__or2_1
X_12696_ _12696_/A _12719_/B vssd1 vssd1 vccd1 vccd1 _12696_/X sky130_fd_sc_hd__or2_1
XFILLER_159_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17223_ _17280_/S vssd1 vssd1 vccd1 vccd1 _17232_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_174_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17099__A _17180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14435_ _18705_/Q _14432_/C _14434_/Y vssd1 vssd1 vccd1 vccd1 _18705_/D sky130_fd_sc_hd__o21a_1
X_11647_ _11647_/A _11647_/B vssd1 vssd1 vccd1 vccd1 _11648_/C sky130_fd_sc_hd__xnor2_1
Xinput13 io_dbus_rdata[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_4
XFILLER_128_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11928__A1 hold2/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput24 io_dbus_rdata[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_4
XFILLER_174_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17154_ _17691_/A vssd1 vssd1 vccd1 vccd1 _17154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput35 io_ibus_inst[10] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_4
X_14366_ _14427_/A vssd1 vssd1 vccd1 vccd1 _14366_/X sky130_fd_sc_hd__buf_2
X_11578_ _11529_/A _11530_/X _11657_/A _11655_/A vssd1 vssd1 vccd1 vccd1 _11578_/X
+ sky130_fd_sc_hd__a211o_1
Xinput46 io_ibus_inst[20] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput57 io_ibus_inst[30] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16105_ _13150_/X _19075_/Q _16111_/S vssd1 vssd1 vccd1 vccd1 _16106_/A sky130_fd_sc_hd__mux2_1
Xinput68 io_irq_spi_irq vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_4
X_13317_ _13068_/X _13316_/X _13460_/A vssd1 vssd1 vccd1 vccd1 _13317_/Y sky130_fd_sc_hd__a21oi_2
X_10529_ _19242_/Q _19737_/Q _10529_/S vssd1 vssd1 vccd1 vccd1 _10529_/X sky130_fd_sc_hd__mux2_1
X_17085_ _19481_/Q _17084_/X _17088_/S vssd1 vssd1 vccd1 vccd1 _17086_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18422__S _18422_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14297_ _18665_/Q _18664_/Q _18663_/Q _14297_/D vssd1 vssd1 vccd1 vccd1 _14306_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_143_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16036_ _13323_/X _19047_/Q _16042_/S vssd1 vssd1 vccd1 vccd1 _16037_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09349__A2 _12895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13248_ _13248_/A _13248_/B vssd1 vssd1 vccd1 vccd1 _17049_/A sky130_fd_sc_hd__nor2_4
XFILLER_124_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13179_ _17036_/A vssd1 vssd1 vccd1 vccd1 _17678_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17987_ _19861_/Q _17039_/X _17987_/S vssd1 vssd1 vccd1 vccd1 _17988_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16877__S _16881_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11539__S0 _09635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19726_ _19726_/CLK _19726_/D vssd1 vssd1 vccd1 vccd1 _19726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16938_ _16323_/X _19428_/Q _16942_/S vssd1 vssd1 vccd1 vccd1 _16939_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10667__A1 _10674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19657_ _19947_/CLK _19657_/D vssd1 vssd1 vccd1 vccd1 _19657_/Q sky130_fd_sc_hd__dfxtp_1
X_16869_ _16869_/A vssd1 vssd1 vccd1 vccd1 _19397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10762__S1 _10664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ _09410_/A _09410_/B _09410_/C _09410_/D vssd1 vssd1 vccd1 vccd1 _09410_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18608_ _18734_/CLK _18608_/D vssd1 vssd1 vccd1 vccd1 _18608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19588_ _19974_/CLK _19588_/D vssd1 vssd1 vccd1 vccd1 _19588_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09904__S0 _11566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ _09418_/B vssd1 vssd1 vccd1 vccd1 _09341_/X sky130_fd_sc_hd__clkbuf_4
X_18539_ _18548_/CLK _18539_/D vssd1 vssd1 vccd1 vccd1 _18539_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__15810__A _15813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ _09272_/A _09306_/C _09272_/C vssd1 vssd1 vccd1 vccd1 _09275_/C sky130_fd_sc_hd__and3_1
XFILLER_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13369__B1 _13368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17472__A _17483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10658__A1 _10822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10753__S1 _10638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ _10497_/A vssd1 vssd1 vccd1 vccd1 _10492_/A sky130_fd_sc_hd__buf_2
XFILLER_16_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13505__A _18996_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10880_ _09685_/A _10871_/Y _10875_/Y _10879_/Y _09874_/A vssd1 vssd1 vccd1 vccd1
+ _10880_/X sky130_fd_sc_hd__o311a_1
XFILLER_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ _09539_/A vssd1 vssd1 vccd1 vccd1 _09540_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10505__S1 _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _12550_/A _12550_/B vssd1 vssd1 vccd1 vccd1 _12551_/A sky130_fd_sc_hd__xnor2_4
XFILLER_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11501_ _19205_/Q _19796_/Q _19958_/Q _19173_/Q _10787_/X _10788_/X vssd1 vssd1 vccd1
+ vccd1 _11502_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10830__A1 _09686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12481_ _18471_/Q _12343_/X _12522_/A _12479_/X _12480_/X vssd1 vssd1 vccd1 vccd1
+ _12481_/X sky130_fd_sc_hd__o221a_1
XANTENNA__16027__S _16031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14336__A _18676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14220_ _18935_/Q _18933_/Q _18930_/Q _18929_/Q vssd1 vssd1 vccd1 vccd1 _14220_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11432_ _18424_/Q _19453_/Q _19490_/Q _19064_/Q _11154_/A _11107_/A vssd1 vssd1 vccd1
+ vccd1 _11432_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14151_ _14407_/A vssd1 vssd1 vccd1 vccd1 _14189_/A sky130_fd_sc_hd__buf_2
X_11363_ _09880_/A _11347_/X _11361_/Y _09910_/A _12956_/B vssd1 vssd1 vccd1 vccd1
+ _12825_/B sky130_fd_sc_hd__o32a_2
XFILLER_153_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13102_ _19890_/Q _13209_/B vssd1 vssd1 vccd1 vccd1 _13102_/X sky130_fd_sc_hd__and2_1
X_10314_ _19246_/Q _19741_/Q _10314_/S vssd1 vssd1 vccd1 vccd1 _10314_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14082_ _14090_/A _14086_/C vssd1 vssd1 vccd1 vccd1 _14082_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11269__A2_N _11223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11294_ _11186_/S _11272_/Y _11293_/Y _11015_/A vssd1 vssd1 vccd1 vccd1 _11294_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_112_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17910_ _17910_/A vssd1 vssd1 vccd1 vccd1 _19826_/D sky130_fd_sc_hd__clkbuf_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _14278_/B _12889_/A _11794_/X _18620_/Q vssd1 vssd1 vccd1 vccd1 _13033_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10245_ _10245_/A vssd1 vssd1 vccd1 vccd1 _11642_/B sky130_fd_sc_hd__inv_2
XANTENNA__10346__B1 _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18890_ _18923_/CLK _18890_/D vssd1 vssd1 vccd1 vccd1 _18890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17841_ _19796_/Q _17036_/X _17843_/S vssd1 vssd1 vccd1 vccd1 _17842_/A sky130_fd_sc_hd__mux2_1
X_10176_ _15974_/B _12860_/C vssd1 vssd1 vccd1 vccd1 _10246_/A sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_51_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16697__S _16703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17772_ _17772_/A vssd1 vssd1 vccd1 vccd1 _19765_/D sky130_fd_sc_hd__clkbuf_1
X_14984_ _14984_/A vssd1 vssd1 vccd1 vccd1 _14984_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19511_ _19966_/CLK _19511_/D vssd1 vssd1 vccd1 vccd1 _19511_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10649__A1 _09820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16723_ _19333_/Q _13800_/X _16725_/S vssd1 vssd1 vccd1 vccd1 _16724_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13935_ _13936_/B _13936_/C _18553_/Q vssd1 vssd1 vccd1 vccd1 _13937_/B sky130_fd_sc_hd__a21oi_1
XFILLER_19_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10744__S1 _10626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19442_ _19966_/CLK _19442_/D vssd1 vssd1 vccd1 vccd1 _19442_/Q sky130_fd_sc_hd__dfxtp_1
X_16654_ _16676_/A vssd1 vssd1 vccd1 vccd1 _16663_/S sky130_fd_sc_hd__clkbuf_8
X_13866_ _13879_/A vssd1 vssd1 vccd1 vccd1 _15807_/A sky130_fd_sc_hd__buf_6
X_15605_ _18884_/Q _18916_/Q _15611_/S vssd1 vssd1 vccd1 vccd1 _15606_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12817_ _13900_/A vssd1 vssd1 vccd1 vccd1 _12820_/A sky130_fd_sc_hd__clkbuf_2
X_19373_ _19644_/CLK _19373_/D vssd1 vssd1 vccd1 vccd1 _19373_/Q sky130_fd_sc_hd__dfxtp_1
X_16585_ _19272_/Q _13810_/X _16591_/S vssd1 vssd1 vccd1 vccd1 _16586_/A sky130_fd_sc_hd__mux2_1
X_13797_ _17033_/A vssd1 vssd1 vccd1 vccd1 _13797_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13063__A2 _12906_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18324_ _17697_/X _19996_/Q _18324_/S vssd1 vssd1 vccd1 vccd1 _18325_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15536_ _12766_/Y _15458_/X _15535_/X _15954_/A vssd1 vssd1 vccd1 vccd1 _15536_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12338_/A _12746_/X _12747_/Y vssd1 vssd1 vccd1 vccd1 _12748_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18255_ _19965_/Q _17700_/A _18263_/S vssd1 vssd1 vccd1 vccd1 _18256_/A sky130_fd_sc_hd__mux2_1
X_15467_ _15419_/X _15229_/X _15466_/X _15428_/X vssd1 vssd1 vccd1 vccd1 _15467_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10774__A _10824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ _18782_/Q _12679_/B _12679_/C vssd1 vssd1 vccd1 vccd1 _12700_/B sky130_fd_sc_hd__and3_1
XFILLER_31_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17206_ _17208_/A _17206_/B vssd1 vssd1 vccd1 vccd1 _17207_/A sky130_fd_sc_hd__and2_1
X_14418_ _14422_/C _14419_/C _18701_/Q vssd1 vssd1 vccd1 vccd1 _14420_/B sky130_fd_sc_hd__a21oi_1
X_18186_ _18186_/A vssd1 vssd1 vccd1 vccd1 _19934_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12023__B1 _13650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15398_ _15384_/X _15392_/Y _15397_/Y vssd1 vssd1 vccd1 vccd1 _15399_/C sky130_fd_sc_hd__a21oi_1
XFILLER_129_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17137_ _17137_/A vssd1 vssd1 vccd1 vccd1 _19501_/D sky130_fd_sc_hd__clkbuf_1
X_14349_ _14350_/B _14350_/C _18681_/Q vssd1 vssd1 vccd1 vccd1 _14351_/B sky130_fd_sc_hd__a21oi_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18152__S _18158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17068_ _17068_/A vssd1 vssd1 vccd1 vccd1 _17068_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16019_ _16019_/A vssd1 vssd1 vccd1 vccd1 _19039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09890_ _19221_/Q _19812_/Q _19974_/Q _19189_/Q _11553_/A _09826_/A vssd1 vssd1 vccd1
+ vccd1 _09891_/B sky130_fd_sc_hd__mux4_1
XFILLER_98_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10888__A1 _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16400__S _16400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19709_ _19935_/CLK _19709_/D vssd1 vssd1 vccd1 vccd1 _19709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09803__A _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__B1 _15789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18327__S _18335_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _18937_/Q _09468_/A vssd1 vssd1 vccd1 vccd1 _09696_/B sky130_fd_sc_hd__or2b_1
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10273__C1 _09876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10812__A1 _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11160__S1 _11015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09255_ _18988_/Q _18987_/Q _18986_/Q vssd1 vssd1 vccd1 vccd1 _11920_/C sky130_fd_sc_hd__or3_2
XFILLER_138_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09186_ _09230_/A _09283_/A vssd1 vssd1 vccd1 vccd1 _14755_/A sky130_fd_sc_hd__nand2_2
XANTENNA__15751__A1 _11982_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_162_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _18993_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_119_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15503__A1 _12693_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13514__A0 _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_177_clock _18998_/CLK vssd1 vssd1 vccd1 vccd1 _18858_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10030_ _10093_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10030_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10879__A1 _10824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_clock clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 _18998_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_100_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19998_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09713__A _10434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11981_ _09882_/A _11347_/X _11361_/Y _09911_/A _12956_/B vssd1 vssd1 vccd1 vccd1
+ _11981_/Y sky130_fd_sc_hd__o32ai_4
XANTENNA__13293__A2 _11683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13720_ _12422_/X _13719_/X _13514_/S vssd1 vssd1 vccd1 vccd1 _13720_/X sky130_fd_sc_hd__a21bo_1
X_10932_ _11006_/A _10932_/B vssd1 vssd1 vccd1 vccd1 _10932_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13651_ _13650_/X _11764_/X _13517_/A vssd1 vssd1 vccd1 vccd1 _13651_/X sky130_fd_sc_hd__a21bo_1
X_10863_ _19331_/Q _19602_/Q _19826_/Q _19570_/Q _10787_/X _10788_/X vssd1 vssd1 vccd1
+ vccd1 _10863_/X sky130_fd_sc_hd__mux4_1
XANTENNA__18237__S _18241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_115_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19941_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ _12599_/A _12601_/Y _12697_/S vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__mux2_1
X_16370_ _16370_/A vssd1 vssd1 vccd1 vccd1 _19181_/D sky130_fd_sc_hd__clkbuf_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13593_/B _13582_/B vssd1 vssd1 vccd1 vccd1 _13582_/Y sky130_fd_sc_hd__nand2_2
X_10794_ _20021_/Q _19859_/Q _19268_/Q _19038_/Q _10787_/X _10793_/X vssd1 vssd1 vccd1
+ vccd1 _10795_/B sky130_fd_sc_hd__mux4_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10264__C1 _09555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15321_ _15321_/A _15321_/B vssd1 vssd1 vccd1 vccd1 _15321_/Y sky130_fd_sc_hd__nor2_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _12530_/X _12531_/Y _12582_/C _12425_/X vssd1 vssd1 vccd1 vccd1 _12533_/Y
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__10594__A _10824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16980__S _16986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18040_ _18836_/Q _12347_/A _16072_/B vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__a21o_1
XFILLER_8_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15252_ _15211_/X _15254_/B _15212_/X _15251_/X vssd1 vssd1 vccd1 vccd1 _15252_/X
+ sky130_fd_sc_hd__o211a_1
X_12464_ _12464_/A _14880_/A vssd1 vssd1 vccd1 vccd1 _12495_/A sky130_fd_sc_hd__nor2_1
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14203_ _14427_/A vssd1 vssd1 vccd1 vccd1 _14203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11415_ _19128_/Q _19389_/Q _19288_/Q _19623_/Q _09586_/A _11208_/A vssd1 vssd1 vccd1
+ vccd1 _11415_/X sky130_fd_sc_hd__mux4_2
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15183_ _15183_/A vssd1 vssd1 vccd1 vccd1 _15348_/S sky130_fd_sc_hd__clkinv_2
XFILLER_125_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12395_ _14744_/B vssd1 vssd1 vccd1 vccd1 _16066_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_165_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14134_ _14143_/A _14134_/B _14134_/C vssd1 vssd1 vccd1 vccd1 _18617_/D sky130_fd_sc_hd__nor3_1
XFILLER_125_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11346_ _11311_/A _11345_/X _11181_/X vssd1 vssd1 vccd1 vccd1 _11346_/Y sky130_fd_sc_hd__o21ai_1
X_19991_ _20020_/CLK _19991_/D vssd1 vssd1 vccd1 vccd1 _19991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14065_ _14065_/A vssd1 vssd1 vccd1 vccd1 _14070_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18942_ _18975_/CLK _18942_/D vssd1 vssd1 vccd1 vccd1 _18942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11277_ _19131_/Q _19392_/Q _19291_/Q _19626_/Q _11121_/S _11077_/X vssd1 vssd1 vccd1
+ vccd1 _11278_/B sky130_fd_sc_hd__mux4_1
XFILLER_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13016_ _19486_/Q vssd1 vssd1 vccd1 vccd1 _13359_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__10414__S0 _10314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ _10438_/A _10227_/X _10159_/X vssd1 vssd1 vccd1 vccd1 _10228_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18873_ _18911_/CLK _18873_/D vssd1 vssd1 vccd1 vccd1 _18873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17824_ _19788_/Q _17010_/X _17832_/S vssd1 vssd1 vccd1 vccd1 _17825_/A sky130_fd_sc_hd__mux2_1
X_10159_ _10382_/A vssd1 vssd1 vccd1 vccd1 _10159_/X sky130_fd_sc_hd__buf_2
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14967_ _14830_/X _14856_/X _14965_/Y _15007_/B vssd1 vssd1 vccd1 vccd1 _14972_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__09488__A1 _12393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17755_ _17755_/A vssd1 vssd1 vccd1 vccd1 _19757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13145__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16706_ _19325_/Q _13774_/X _16714_/S vssd1 vssd1 vccd1 vccd1 _16707_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13918_ _18601_/Q _18603_/Q _18602_/Q _14073_/A vssd1 vssd1 vccd1 vccd1 _14081_/A
+ sky130_fd_sc_hd__and4_1
X_17686_ _17684_/X _19734_/Q _17698_/S vssd1 vssd1 vccd1 vccd1 _17687_/A sky130_fd_sc_hd__mux2_1
X_14898_ _14898_/A vssd1 vssd1 vccd1 vccd1 _15078_/B sky130_fd_sc_hd__buf_2
XFILLER_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19425_ _20016_/CLK _19425_/D vssd1 vssd1 vccd1 vccd1 _19425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13849_ _18514_/Q _13848_/X _13852_/S vssd1 vssd1 vccd1 vccd1 _13850_/A sky130_fd_sc_hd__mux2_1
X_16637_ _16323_/X _19295_/Q _16641_/S vssd1 vssd1 vccd1 vccd1 _16638_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18147__S _18147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15430__B1 _15429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19356_ _19981_/CLK _19356_/D vssd1 vssd1 vccd1 vccd1 _19356_/Q sky130_fd_sc_hd__dfxtp_1
X_16568_ _16568_/A vssd1 vssd1 vccd1 vccd1 _19264_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15981__A1 _19024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12795__A1 _18484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18307_ _17672_/X _19988_/Q _18313_/S vssd1 vssd1 vccd1 vccd1 _18308_/A sky130_fd_sc_hd__mux2_1
X_15519_ _14991_/X _15516_/Y _15518_/X _14998_/X vssd1 vssd1 vccd1 vccd1 _15522_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__16890__S _16892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19287_ _20040_/CLK _19287_/D vssd1 vssd1 vccd1 vccd1 _19287_/Q sky130_fd_sc_hd__dfxtp_1
X_16499_ _16545_/S vssd1 vssd1 vccd1 vccd1 _16508_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18238_ _18238_/A vssd1 vssd1 vccd1 vccd1 _19957_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15733__A1 _18971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13744__A0 _18484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18169_ _17681_/X _19927_/Q _18169_/S vssd1 vssd1 vccd1 vccd1 _18170_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_94_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _20003_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09942_ _09942_/A _09942_/B vssd1 vssd1 vccd1 vccd1 _09942_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12224__A _12234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10405__S0 _09995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ _09873_/A vssd1 vssd1 vccd1 vccd1 _09874_/A sky130_fd_sc_hd__buf_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17226__S _17232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15254__B _15254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19986_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12894__A _13215_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14775__A2 _09279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09307_ _09492_/A _09491_/A vssd1 vssd1 vccd1 vccd1 _12831_/A sky130_fd_sc_hd__and2_4
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17896__S _17904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19861_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14317__C _18669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09238_ _18973_/Q vssd1 vssd1 vccd1 vccd1 _09284_/A sky130_fd_sc_hd__inv_2
XFILLER_103_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13735__A0 _18483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ _18967_/Q vssd1 vssd1 vccd1 vccd1 _09283_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_119_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16305__S _16314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14614__A _14648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _19356_/Q _19691_/Q _11270_/S vssd1 vssd1 vccd1 vccd1 _11200_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10644__S0 _09726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ _12217_/A _14906_/A vssd1 vssd1 vccd1 vccd1 _12182_/A sky130_fd_sc_hd__and2_1
XFILLER_150_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11131_ _11131_/A _11131_/B vssd1 vssd1 vccd1 vccd1 _11131_/X sky130_fd_sc_hd__or2_1
XFILLER_162_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11062_ _11421_/A vssd1 vssd1 vccd1 vccd1 _11283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17136__S _17145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ _10013_/A vssd1 vssd1 vccd1 vccd1 _10082_/A sky130_fd_sc_hd__buf_4
XFILLER_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15445__A _15449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15870_ input49/X _15834_/X _15789_/X _09328_/Y vssd1 vssd1 vccd1 vccd1 _16843_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16040__S _16042_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input22_A io_dbus_rdata[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ _14821_/A _14821_/B vssd1 vssd1 vccd1 vccd1 _14822_/D sky130_fd_sc_hd__nor2_1
XFILLER_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16975__S _16975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17540_ _19676_/Q vssd1 vssd1 vccd1 vccd1 _17541_/A sky130_fd_sc_hd__clkbuf_1
X_14752_ _12055_/B _12055_/C _14750_/X _14808_/A _09508_/A vssd1 vssd1 vccd1 vccd1
+ _14752_/X sky130_fd_sc_hd__o311a_1
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11964_ _11964_/A _14901_/A vssd1 vssd1 vccd1 vccd1 _11971_/A sky130_fd_sc_hd__xnor2_4
XFILLER_45_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13703_ _13732_/A _19019_/Q vssd1 vssd1 vccd1 vccd1 _13703_/Y sky130_fd_sc_hd__nand2_1
X_17471_ _17471_/A vssd1 vssd1 vccd1 vccd1 _19642_/D sky130_fd_sc_hd__clkbuf_1
X_10915_ _09702_/A _10903_/X _10914_/X _09842_/A _18843_/Q vssd1 vssd1 vccd1 vccd1
+ _12837_/B sky130_fd_sc_hd__a32o_4
XANTENNA__11372__S1 _10972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14683_ _18794_/Q hold7/X _14683_/S vssd1 vssd1 vccd1 vccd1 _14684_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11895_ _18670_/Q _11889_/X _11892_/X _11893_/X _11894_/X vssd1 vssd1 vccd1 vccd1
+ _11896_/B sky130_fd_sc_hd__a2111o_2
XANTENNA_output109_A _12822_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19210_ _20027_/CLK _19210_/D vssd1 vssd1 vccd1 vccd1 _19210_/Q sky130_fd_sc_hd__dfxtp_1
X_16422_ _19200_/Q _13784_/X _16424_/S vssd1 vssd1 vccd1 vccd1 _16423_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13634_ _18469_/Q _13633_/X _13670_/S vssd1 vssd1 vccd1 vccd1 _13635_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10846_ _20020_/Q _19858_/Q _19267_/Q _19037_/Q _10797_/X _10793_/X vssd1 vssd1 vccd1
+ vccd1 _10846_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12777__A1 _12260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19141_ _19636_/CLK _19141_/D vssd1 vssd1 vccd1 vccd1 _19141_/Q sky130_fd_sc_hd__dfxtp_1
X_16353_ _16352_/X _19176_/Q _16362_/S vssd1 vssd1 vccd1 vccd1 _16354_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12777__B2 _11945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13565_ _18872_/Q _13565_/B vssd1 vssd1 vccd1 vccd1 _13565_/Y sky130_fd_sc_hd__nand2_1
X_10777_ _18436_/Q _19465_/Q _19502_/Q _19076_/Q _10776_/X _10710_/A vssd1 vssd1 vccd1
+ vccd1 _10777_/X sky130_fd_sc_hd__mux4_2
XFILLER_157_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15304_ _15284_/X _15301_/Y _15303_/X _15268_/X vssd1 vssd1 vccd1 vccd1 _15308_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19072_ _19567_/CLK _19072_/D vssd1 vssd1 vccd1 vccd1 _19072_/Q sky130_fd_sc_hd__dfxtp_1
X_12516_ _15410_/A _12516_/B vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__xnor2_4
X_16284_ _16284_/A vssd1 vssd1 vccd1 vccd1 _19153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10883__S0 _10919_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13496_ _13188_/A _18864_/Q _12957_/A vssd1 vssd1 vccd1 vccd1 _13496_/X sky130_fd_sc_hd__a21o_1
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18023_ _18023_/A vssd1 vssd1 vccd1 vccd1 _19877_/D sky130_fd_sc_hd__clkbuf_1
X_15235_ _15218_/X _15230_/Y _15234_/Y vssd1 vssd1 vccd1 vccd1 _15236_/C sky130_fd_sc_hd__a21oi_1
XFILLER_8_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12447_ _12447_/A _12501_/C vssd1 vssd1 vccd1 vccd1 _12447_/X sky130_fd_sc_hd__or2_1
XANTENNA__16215__S _16217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output90_A _12717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15166_ _15021_/X _15034_/X _15189_/S vssd1 vssd1 vccd1 vccd1 _15166_/X sky130_fd_sc_hd__mux2_1
X_12378_ _12378_/A vssd1 vssd1 vccd1 vccd1 _12378_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_126_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14117_ _18731_/Q _18730_/Q _18732_/Q _14488_/A vssd1 vssd1 vccd1 vccd1 _14496_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__11752__A2 _13081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _19915_/Q _19529_/Q _19979_/Q _19098_/Q _11328_/X _11322_/X vssd1 vssd1 vccd1
+ vccd1 _11330_/B sky130_fd_sc_hd__mux4_1
X_19974_ _19974_/CLK _19974_/D vssd1 vssd1 vccd1 vccd1 _19974_/Q sky130_fd_sc_hd__dfxtp_1
X_15097_ _15097_/A vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14048_ _14051_/B _14051_/C _14019_/X vssd1 vssd1 vccd1 vccd1 _14048_/Y sky130_fd_sc_hd__a21oi_1
X_18925_ _18926_/CLK _18925_/D vssd1 vssd1 vccd1 vccd1 _18925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11883__A _14159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18856_ _19025_/CLK _18856_/D vssd1 vssd1 vccd1 vccd1 _18856_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17807_ _17807_/A vssd1 vssd1 vccd1 vccd1 _19781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18787_ _19912_/CLK _18787_/D vssd1 vssd1 vccd1 vccd1 _18787_/Q sky130_fd_sc_hd__dfxtp_1
X_15999_ _15999_/A vssd1 vssd1 vccd1 vccd1 _19030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17738_ _17738_/A _17738_/B vssd1 vssd1 vccd1 vccd1 _17795_/A sky130_fd_sc_hd__or2_4
XFILLER_36_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17669_ _17736_/S vssd1 vssd1 vccd1 vccd1 _17682_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_36_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16186__A _16208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15403__B1 _15402_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19408_ _19996_/CLK _19408_/D vssd1 vssd1 vccd1 vccd1 _19408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19339_ _20028_/CLK _19339_/D vssd1 vssd1 vccd1 vccd1 _19339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_173_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10962__A _11023_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15182__A2 _15177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16125__S _16133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14434__A _14472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18340__S _18346_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09925_ _19348_/Q _19619_/Q _19843_/Q _19587_/Q _09659_/S _09614_/A vssd1 vssd1 vccd1
+ vccd1 _09925_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12889__A _12889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13496__A2 _18864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09856_ _19684_/Q _19450_/Q _18515_/Q _19780_/Q _11532_/S _09660_/A vssd1 vssd1 vccd1
+ vccd1 _09856_/X sky130_fd_sc_hd__mux4_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_98_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09263__A _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16795__S _16797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09787_ _19387_/Q vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15642__A0 _18900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12456__B1 _12455_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15712__B _15740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _09883_/A _10687_/X _10698_/X _09912_/A _10699_/Y vssd1 vssd1 vccd1 vccd1
+ _12844_/A sky130_fd_sc_hd__o32a_4
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13513__A _13520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11697_/A _11680_/B _11697_/C vssd1 vssd1 vccd1 vccd1 _11688_/A sky130_fd_sc_hd__or3_4
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10631_ _10749_/S vssd1 vssd1 vccd1 vccd1 _10637_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13350_ _13348_/X _13349_/X _13350_/S vssd1 vssd1 vccd1 vccd1 _13350_/X sky130_fd_sc_hd__mux2_1
X_10562_ _19930_/Q _19544_/Q _19994_/Q _19113_/Q _10521_/X _10522_/X vssd1 vssd1 vccd1
+ vccd1 _10563_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12301_ _12301_/A _12301_/B vssd1 vssd1 vccd1 vccd1 _12301_/X sky130_fd_sc_hd__xor2_4
XFILLER_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13281_ _13268_/X _13279_/Y _13280_/Y vssd1 vssd1 vccd1 vccd1 _17055_/A sky130_fd_sc_hd__a21oi_4
X_10493_ _19242_/Q _19737_/Q _10493_/S vssd1 vssd1 vccd1 vccd1 _10493_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15020_ _15020_/A vssd1 vssd1 vccd1 vccd1 _15114_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_136_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12232_ _12231_/A _12255_/C _13700_/A vssd1 vssd1 vccd1 vccd1 _12232_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12163_ _16075_/A _12163_/B _12163_/C vssd1 vssd1 vccd1 vccd1 _16072_/A sky130_fd_sc_hd__nor3_2
XANTENNA__18250__S _18252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11114_ _19135_/Q _19396_/Q _19295_/Q _19630_/Q _09721_/A _10854_/A vssd1 vssd1 vccd1
+ vccd1 _11115_/B sky130_fd_sc_hd__mux4_1
X_16971_ _16371_/X _19443_/Q _16975_/S vssd1 vssd1 vccd1 vccd1 _16972_/A sky130_fd_sc_hd__mux2_1
X_12094_ _12215_/A _12215_/B vssd1 vssd1 vccd1 vccd1 _12094_/X sky130_fd_sc_hd__xor2_4
XFILLER_110_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13487__A2 _13290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18710_ _18993_/CLK _18710_/D vssd1 vssd1 vccd1 vccd1 _18710_/Q sky130_fd_sc_hd__dfxtp_1
X_11045_ _11320_/A vssd1 vssd1 vccd1 vccd1 _11045_/X sky130_fd_sc_hd__clkbuf_4
X_15922_ _15946_/A vssd1 vssd1 vccd1 vccd1 _15955_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09786__S1 _09768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19690_ _20012_/CLK _19690_/D vssd1 vssd1 vccd1 vccd1 _19690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18641_ _18688_/CLK _18641_/D vssd1 vssd1 vccd1 vccd1 _18641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15853_ _12032_/X _15842_/X _15843_/X input43/X vssd1 vssd1 vccd1 vccd1 _17206_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_0_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_14804_ _14804_/A _14804_/B _14804_/C _14804_/D vssd1 vssd1 vccd1 vccd1 _14822_/C
+ sky130_fd_sc_hd__nor4_1
XANTENNA__11208__A _11208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18572_ _19023_/CLK _18572_/D vssd1 vssd1 vccd1 vccd1 _18572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15784_ _12316_/A _11867_/X _15783_/X _13885_/X vssd1 vssd1 vccd1 vccd1 _18960_/D
+ sky130_fd_sc_hd__o211a_1
X_12996_ _13535_/A _13015_/C vssd1 vssd1 vccd1 vccd1 _12996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12030__C _15094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17523_ _17523_/A vssd1 vssd1 vccd1 vccd1 _19667_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11345__S1 _11108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11947_ _12845_/A _14819_/B _11947_/C vssd1 vssd1 vccd1 vccd1 _14815_/A sky130_fd_sc_hd__nand3_1
X_14735_ _14735_/A vssd1 vssd1 vccd1 vccd1 _18817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17454_ _17454_/A vssd1 vssd1 vccd1 vccd1 _19634_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _15883_/A vssd1 vssd1 vccd1 vccd1 _15813_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11878_ _11897_/A _19017_/Q vssd1 vssd1 vccd1 vccd1 _11878_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14238__B _14242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16405_ _19192_/Q _13754_/X _16413_/S vssd1 vssd1 vccd1 vccd1 _16406_/A sky130_fd_sc_hd__mux2_1
X_13617_ _18467_/Q _13616_/X _13617_/S vssd1 vssd1 vccd1 vccd1 _13618_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10829_ _09624_/A _10828_/X _10719_/X vssd1 vssd1 vccd1 vccd1 _10829_/Y sky130_fd_sc_hd__o21ai_1
X_17385_ _19604_/Q _17036_/X _17387_/S vssd1 vssd1 vccd1 vccd1 _17386_/A sky130_fd_sc_hd__mux2_1
X_14597_ _14648_/A vssd1 vssd1 vccd1 vccd1 _14612_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19124_ _19747_/CLK _19124_/D vssd1 vssd1 vccd1 vccd1 _19124_/Q sky130_fd_sc_hd__dfxtp_1
X_16336_ _17672_/A vssd1 vssd1 vccd1 vccd1 _16336_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13548_ _13546_/X _13547_/Y _13583_/S vssd1 vssd1 vccd1 vccd1 _13548_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16267_ _13263_/X _19146_/Q _16269_/S vssd1 vssd1 vccd1 vccd1 _16268_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19055_ _19055_/CLK _19055_/D vssd1 vssd1 vccd1 vccd1 _19055_/Q sky130_fd_sc_hd__dfxtp_1
X_13479_ _13474_/X _13477_/X _13478_/X vssd1 vssd1 vccd1 vccd1 _17090_/A sky130_fd_sc_hd__o21a_2
XFILLER_69_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18006_ _18006_/A vssd1 vssd1 vccd1 vccd1 _19869_/D sky130_fd_sc_hd__clkbuf_1
X_15218_ _15305_/A vssd1 vssd1 vccd1 vccd1 _15218_/X sky130_fd_sc_hd__clkbuf_2
X_16198_ _13302_/X _19116_/Q _16206_/S vssd1 vssd1 vccd1 vccd1 _16199_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15149_ _12094_/X _15146_/X _15951_/A vssd1 vssd1 vccd1 vccd1 _15149_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19957_ _19957_/CLK _19957_/D vssd1 vssd1 vccd1 vccd1 _19957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14675__A1 _14554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09710_ _10643_/A vssd1 vssd1 vccd1 vccd1 _10572_/A sky130_fd_sc_hd__buf_2
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15872__B1 _15788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11489__A1 _09830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18908_ _18911_/CLK _18908_/D vssd1 vssd1 vccd1 vccd1 _18908_/Q sky130_fd_sc_hd__dfxtp_1
X_19888_ _19888_/CLK _19888_/D vssd1 vssd1 vccd1 vccd1 _19888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09641_ _11538_/A _09641_/B vssd1 vssd1 vccd1 vccd1 _09641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18839_ _19950_/CLK _18839_/D vssd1 vssd1 vccd1 vccd1 _18839_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15813__A _15813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ _11001_/A vssd1 vssd1 vccd1 vccd1 _10934_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10022__A _10529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09854__A1 _11533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18335__S _18335_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10847__S0 _10953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09908_ _11574_/A _09908_/B _09908_/C vssd1 vssd1 vccd1 vccd1 _09908_/Y sky130_fd_sc_hd__nor3_1
XFILLER_76_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13874__C1 _17203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20028_ _20028_/CLK _20028_/D vssd1 vssd1 vccd1 vccd1 _20028_/Q sky130_fd_sc_hd__dfxtp_1
X_09839_ _09809_/X _09812_/X _09814_/X _11574_/A _09838_/X vssd1 vssd1 vccd1 vccd1
+ _09839_/X sky130_fd_sc_hd__a311o_1
XFILLER_59_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17414__S _17420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ _12851_/A _12850_/B vssd1 vssd1 vccd1 vccd1 _12850_/Y sky130_fd_sc_hd__nor2_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15091__A1 _11994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09721__A _09721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11801_ _11801_/A vssd1 vssd1 vccd1 vccd1 _13519_/B sky130_fd_sc_hd__inv_2
XFILLER_61_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _15980_/B vssd1 vssd1 vccd1 vccd1 _12781_/Y sky130_fd_sc_hd__inv_2
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14528_/A _14520_/B _14520_/C vssd1 vssd1 vccd1 vccd1 _18740_/D sky130_fd_sc_hd__nor3_1
XFILLER_92_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11732_ _13057_/A vssd1 vssd1 vccd1 vccd1 _11732_/X sky130_fd_sc_hd__buf_2
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14451_ _14450_/A _14450_/B _18716_/Q vssd1 vssd1 vccd1 vccd1 _14452_/C sky130_fd_sc_hd__a21oi_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11663_/A vssd1 vssd1 vccd1 vccd1 _15738_/A sky130_fd_sc_hd__buf_2
XFILLER_14_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13439_/A _13708_/B vssd1 vssd1 vccd1 vccd1 _13402_/Y sky130_fd_sc_hd__nand2_1
X_17170_ _17707_/A vssd1 vssd1 vccd1 vccd1 _17170_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10614_ _10592_/X _10604_/X _10613_/X _10668_/A vssd1 vssd1 vccd1 vccd1 _10614_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14382_ _14399_/A _14382_/B _14391_/D vssd1 vssd1 vccd1 vccd1 _18690_/D sky130_fd_sc_hd__nor3_1
X_11594_ _11594_/A _11594_/B vssd1 vssd1 vccd1 vccd1 _11628_/A sky130_fd_sc_hd__nor2_1
X_16121_ _16121_/A vssd1 vssd1 vccd1 vccd1 _19082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13333_ _18572_/Q _13054_/B _13330_/X _13332_/X vssd1 vssd1 vccd1 vccd1 _13333_/X
+ sky130_fd_sc_hd__o22a_1
X_10545_ _19672_/Q _19438_/Q _18503_/Q _19768_/Q _10493_/S _10587_/A vssd1 vssd1 vccd1
+ vccd1 _10545_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10806__S _11486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16052_ _16052_/A vssd1 vssd1 vccd1 vccd1 _19054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13264_ _13263_/X _18442_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__mux2_1
X_10476_ _10376_/A _10475_/X _10382_/A vssd1 vssd1 vccd1 vccd1 _10476_/X sky130_fd_sc_hd__o21a_1
XFILLER_142_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11168__B1 _09911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15003_ _15055_/S _14996_/B _15438_/A _14999_/X _15002_/Y vssd1 vssd1 vccd1 vccd1
+ _15003_/X sky130_fd_sc_hd__o2111a_1
XFILLER_124_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12215_ _12215_/A _12215_/B _12215_/C _12215_/D vssd1 vssd1 vccd1 vccd1 _12215_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__10107__A _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11263__S0 _11367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13195_ _18596_/Q _13120_/X _13194_/X _18728_/Q vssd1 vssd1 vccd1 vccd1 _13195_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10915__B1 _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14802__A _15147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19811_ _20037_/CLK _19811_/D vssd1 vssd1 vccd1 vccd1 _19811_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17843__A1 _17039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09781__B1 _09837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ _12179_/S vssd1 vssd1 vccd1 vccd1 _12358_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_121_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19742_ _20032_/CLK _19742_/D vssd1 vssd1 vccd1 vccd1 _19742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16954_ _16954_/A vssd1 vssd1 vccd1 vccd1 _19435_/D sky130_fd_sc_hd__clkbuf_1
X_12077_ _12077_/A vssd1 vssd1 vccd1 vccd1 _12077_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15905_ _18995_/Q _15904_/X _15914_/S vssd1 vssd1 vccd1 vccd1 _15906_/A sky130_fd_sc_hd__mux2_1
X_11028_ _19328_/Q _19599_/Q _19823_/Q _19567_/Q _10892_/A _11157_/A vssd1 vssd1 vccd1
+ vccd1 _11028_/X sky130_fd_sc_hd__mux4_1
X_19673_ _19995_/CLK _19673_/D vssd1 vssd1 vccd1 vccd1 _19673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16885_ _16885_/A vssd1 vssd1 vccd1 vccd1 _19404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14948__S _14948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17324__S _17326_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13852__S _13852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18624_ _18655_/CLK _18624_/D vssd1 vssd1 vccd1 vccd1 _18624_/Q sky130_fd_sc_hd__dfxtp_1
X_15836_ _15871_/A _15836_/B vssd1 vssd1 vccd1 vccd1 _18973_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10139__A2_N _09539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09631__A _10073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18555_ _19883_/CLK _18555_/D vssd1 vssd1 vccd1 vccd1 _18555_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _14749_/A _15765_/X _15766_/X _15756_/X vssd1 vssd1 vccd1 vccd1 _18952_/D
+ sky130_fd_sc_hd__o211a_1
X_12979_ _12978_/X _18427_/Q _13003_/S vssd1 vssd1 vccd1 vccd1 _12980_/A sky130_fd_sc_hd__mux2_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17506_ _19659_/Q vssd1 vssd1 vccd1 vccd1 _17507_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14718_ _14729_/A vssd1 vssd1 vccd1 vccd1 _14727_/S sky130_fd_sc_hd__clkbuf_2
X_18486_ _19946_/CLK _18486_/D vssd1 vssd1 vccd1 vccd1 _18486_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15698_ _15698_/A vssd1 vssd1 vccd1 vccd1 _18925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17437_ _17112_/X _19627_/Q _17437_/S vssd1 vssd1 vccd1 vccd1 _17438_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14649_ _18783_/Q _13710_/X _14649_/S vssd1 vssd1 vccd1 vccd1 _14650_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_46_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17368_ _19596_/Q _17010_/X _17376_/S vssd1 vssd1 vccd1 vccd1 _17369_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19107_ _19637_/CLK _19107_/D vssd1 vssd1 vccd1 vccd1 _19107_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17994__S _17998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16319_ _16319_/A vssd1 vssd1 vccd1 vccd1 _19165_/D sky130_fd_sc_hd__clkbuf_1
X_17299_ _17299_/A vssd1 vssd1 vccd1 vccd1 _19565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19038_ _19633_/CLK _19038_/D vssd1 vssd1 vccd1 vccd1 _19038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput101 _12221_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[8] sky130_fd_sc_hd__buf_2
XANTENNA__11159__B1 _11227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput112 _12841_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[12] sky130_fd_sc_hd__buf_2
XANTENNA__17295__A _17352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput123 _12854_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[22] sky130_fd_sc_hd__buf_2
XFILLER_99_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput134 _12826_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[3] sky130_fd_sc_hd__buf_2
XANTENNA__10017__A _10380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput145 _12352_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[12] sky130_fd_sc_hd__buf_2
Xoutput156 _12608_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[22] sky130_fd_sc_hd__buf_2
XFILLER_88_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09806__A _09806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput167 _12077_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13320__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17598__A0 _17147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09624_ _09624_/A vssd1 vssd1 vccd1 vccd1 _10674_/A sky130_fd_sc_hd__buf_2
XFILLER_110_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11882__A1 _12060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09555_ _09555_/A vssd1 vssd1 vccd1 vccd1 _09862_/A sky130_fd_sc_hd__buf_2
XFILLER_102_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11790__B _11790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13084__B1 _13077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14159__A _14159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14820__A1 _09522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _15624_/A vssd1 vssd1 vccd1 vccd1 _15945_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12407__A _12459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10330_ _19246_/Q _19741_/Q _10330_/S vssd1 vssd1 vccd1 vccd1 _10330_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14887__A1 _15410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17409__S _17409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ _10261_/A vssd1 vssd1 vccd1 vccd1 _10261_/X sky130_fd_sc_hd__buf_2
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12000_ _12279_/B vssd1 vssd1 vccd1 vccd1 _12393_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09716__A _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10192_ _10192_/A vssd1 vssd1 vccd1 vccd1 _10192_/X sky130_fd_sc_hd__buf_2
XFILLER_79_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14639__A1 _11879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__B2 _18854_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11548__S1 _09660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17589__A0 _17135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13951_ _13956_/B _13956_/C _11884_/X vssd1 vssd1 vccd1 vccd1 _13951_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16549__A _16617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12902_ _12936_/A _18865_/Q vssd1 vssd1 vccd1 vccd1 _12902_/X sky130_fd_sc_hd__or2_1
XFILLER_47_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16670_ _16371_/X _19310_/Q _16674_/S vssd1 vssd1 vccd1 vccd1 _16671_/A sky130_fd_sc_hd__mux2_1
X_13882_ _12312_/A _12312_/B _14447_/B vssd1 vssd1 vccd1 vccd1 _18529_/D sky130_fd_sc_hd__a21o_1
XANTENNA__11873__A1 _12060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16261__A0 _13219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12833_ _12833_/A vssd1 vssd1 vccd1 vccd1 _12844_/B sky130_fd_sc_hd__buf_6
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ _15621_/A vssd1 vssd1 vccd1 vccd1 _18891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _17720_/X _20003_/Q _18346_/S vssd1 vssd1 vccd1 vccd1 _18341_/A sky130_fd_sc_hd__mux2_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15552_/A vssd1 vssd1 vccd1 vccd1 _15552_/Y sky130_fd_sc_hd__inv_2
X_12764_ _12742_/A _12742_/B _12741_/A vssd1 vssd1 vccd1 vccd1 _12765_/B sky130_fd_sc_hd__a21o_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _19010_/Q _13227_/A _11714_/Y vssd1 vssd1 vccd1 vccd1 _11715_/X sky130_fd_sc_hd__or3b_1
X_14503_ _14528_/A _14503_/B _14503_/C vssd1 vssd1 vccd1 vccd1 _18734_/D sky130_fd_sc_hd__nor3_1
X_18271_ _18271_/A vssd1 vssd1 vccd1 vccd1 _19972_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _15487_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _15483_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _18543_/Q _18544_/Q _12695_/C vssd1 vssd1 vccd1 vccd1 _12719_/B sky130_fd_sc_hd__and3_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17222_ _17222_/A vssd1 vssd1 vccd1 vccd1 _19531_/D sky130_fd_sc_hd__clkbuf_1
X_11646_ _11645_/A _11645_/B _11645_/C vssd1 vssd1 vccd1 vccd1 _11648_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14434_ _14472_/A _14439_/C vssd1 vssd1 vccd1 vccd1 _14434_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09677__S0 _09855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 io_dbus_rdata[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
Xinput25 io_dbus_rdata[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_4
X_17153_ _17153_/A vssd1 vssd1 vccd1 vccd1 _19506_/D sky130_fd_sc_hd__clkbuf_1
X_14365_ _14399_/A _14365_/B _14365_/C vssd1 vssd1 vccd1 vccd1 _18685_/D sky130_fd_sc_hd__nor3_1
XFILLER_156_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11577_ _15982_/B _12866_/C vssd1 vssd1 vccd1 vccd1 _11655_/A sky130_fd_sc_hd__and2_2
Xinput36 io_ibus_inst[11] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_2
Xinput47 io_ibus_inst[21] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_6
X_16104_ _16104_/A vssd1 vssd1 vccd1 vccd1 _19074_/D sky130_fd_sc_hd__clkbuf_1
Xinput58 io_ibus_inst[31] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13316_ _18854_/Q _13675_/B _13458_/A vssd1 vssd1 vccd1 vccd1 _13316_/X sky130_fd_sc_hd__mux2_1
X_10528_ _19370_/Q _19705_/Q _10573_/S vssd1 vssd1 vccd1 vccd1 _10528_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput69 io_irq_uart_irq vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_8
XFILLER_128_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17084_ _17084_/A vssd1 vssd1 vccd1 vccd1 _17084_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14296_ _18664_/Q _14300_/D _14295_/Y vssd1 vssd1 vccd1 vccd1 _18664_/D sky130_fd_sc_hd__o21a_1
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16035_ _16035_/A vssd1 vssd1 vccd1 vccd1 _19046_/D sky130_fd_sc_hd__clkbuf_1
X_13247_ _13267_/C _13244_/Y _13246_/Y _12960_/A _13223_/A vssd1 vssd1 vccd1 vccd1
+ _13248_/B sky130_fd_sc_hd__o221a_1
X_10459_ _18443_/Q _19472_/Q _19509_/Q _19083_/Q _09995_/A _10400_/A vssd1 vssd1 vccd1
+ vccd1 _10459_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11010__C1 _11133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ _12967_/X _13176_/X _13177_/X vssd1 vssd1 vccd1 vccd1 _17036_/A sky130_fd_sc_hd__o21a_4
XFILLER_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11367__S _11367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _12129_/A _12477_/C vssd1 vssd1 vccd1 vccd1 _12130_/D sky130_fd_sc_hd__nor2_1
X_17986_ _17986_/A vssd1 vssd1 vccd1 vccd1 _19860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11539__S1 _09639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19725_ _19757_/CLK _19725_/D vssd1 vssd1 vccd1 vccd1 _19725_/Q sky130_fd_sc_hd__dfxtp_1
X_16937_ _16937_/A vssd1 vssd1 vccd1 vccd1 _19427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18241__A1 _17681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15363__A _15457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19656_ _19656_/CLK _19656_/D vssd1 vssd1 vccd1 vccd1 _19656_/Q sky130_fd_sc_hd__dfxtp_1
X_16868_ _16326_/X _19397_/Q _16870_/S vssd1 vssd1 vccd1 vccd1 _16869_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18607_ _19941_/CLK _18607_/D vssd1 vssd1 vccd1 vccd1 _18607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15819_ _15819_/A vssd1 vssd1 vccd1 vccd1 _18968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19587_ _19587_/CLK _19587_/D vssd1 vssd1 vccd1 vccd1 _19587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16799_ _16821_/A vssd1 vssd1 vccd1 vccd1 _16808_/S sky130_fd_sc_hd__buf_4
XFILLER_46_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09340_ _18826_/Q _18825_/Q vssd1 vssd1 vccd1 vccd1 _09418_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18538_ _18911_/CLK _18538_/D vssd1 vssd1 vccd1 vccd1 _18538_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10300__A _15966_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09271_ _09313_/A _11951_/B vssd1 vssd1 vccd1 vccd1 _09272_/C sky130_fd_sc_hd__nor2_2
XFILLER_34_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18469_ _18773_/CLK _18469_/D vssd1 vssd1 vccd1 vccd1 _18469_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13369__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13330__B _14555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12227__A _12393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16922__A _16990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11131__A _11131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16133__S _16133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11785__B _11790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09607_ _09607_/A vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13505__B _13505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ _09538_/A vssd1 vssd1 vccd1 vccd1 _09539_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10210__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12280__A1 _12814_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ _18989_/Q vssd1 vssd1 vccd1 vccd1 _09471_/C sky130_fd_sc_hd__buf_4
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16308__S _16314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _11500_/A _11500_/B vssd1 vssd1 vccd1 vccd1 _11500_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14557__A0 _18757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12480_ _12557_/A vssd1 vssd1 vccd1 vccd1 _12480_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14336__B _14336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _11440_/A _11431_/B vssd1 vssd1 vccd1 vccd1 _11431_/X sky130_fd_sc_hd__or2_1
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10356__S _10356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14150_ _14159_/A vssd1 vssd1 vccd1 vccd1 _14407_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11362_ _18835_/Q vssd1 vssd1 vccd1 vccd1 _12956_/B sky130_fd_sc_hd__clkinv_4
XFILLER_152_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13101_ input32/X _13091_/A _13094_/A vssd1 vssd1 vccd1 vccd1 _13113_/A sky130_fd_sc_hd__a21o_1
X_10313_ _19374_/Q _19709_/Q _10313_/S vssd1 vssd1 vccd1 vccd1 _10313_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17139__S _17145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14081_ _14081_/A vssd1 vssd1 vccd1 vccd1 _14086_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_11293_ _11293_/A _19227_/Q vssd1 vssd1 vccd1 vccd1 _11293_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13032_ _18652_/Q vssd1 vssd1 vccd1 vccd1 _14278_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input52_A io_ibus_inst[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10244_ _11639_/A _11647_/A vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__or2_1
XANTENNA__10346__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16978__S _16986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15809__B1 _15798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11187__S _11295_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17840_ _17840_/A vssd1 vssd1 vccd1 vccd1 _19795_/D sky130_fd_sc_hd__clkbuf_1
X_10175_ _09702_/X _10161_/X _10174_/X _09843_/X _18860_/Q vssd1 vssd1 vccd1 vccd1
+ _12860_/C sky130_fd_sc_hd__a32o_4
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13296__A0 _18853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17771_ _17681_/X _19765_/Q _17771_/S vssd1 vssd1 vccd1 vccd1 _17772_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14983_ _15103_/B _14983_/B vssd1 vssd1 vccd1 vccd1 _14984_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10104__B _12856_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19510_ _19997_/CLK _19510_/D vssd1 vssd1 vccd1 vccd1 _19510_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output139_A _12834_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16722_ _16722_/A vssd1 vssd1 vccd1 vccd1 _19332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15183__A _15183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13934_ _13936_/B _13936_/C _13933_/Y vssd1 vssd1 vccd1 vccd1 _18552_/D sky130_fd_sc_hd__o21a_1
XFILLER_75_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19441_ _19996_/CLK _19441_/D vssd1 vssd1 vccd1 vccd1 _19441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ _16653_/A vssd1 vssd1 vccd1 vccd1 _19302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13865_ _13865_/A vssd1 vssd1 vccd1 vccd1 _18519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17602__S _17606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11059__C1 _11058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15604_ _15604_/A vssd1 vssd1 vccd1 vccd1 _18883_/D sky130_fd_sc_hd__clkbuf_1
X_19372_ _19965_/CLK _19372_/D vssd1 vssd1 vccd1 vccd1 _19372_/Q sky130_fd_sc_hd__dfxtp_1
X_12816_ _12522_/X _12814_/X _12815_/X vssd1 vssd1 vccd1 vccd1 _12816_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13021__A1_N _13005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16584_ _16584_/A vssd1 vssd1 vccd1 vccd1 _19271_/D sky130_fd_sc_hd__clkbuf_1
X_13796_ _13796_/A vssd1 vssd1 vccd1 vccd1 _18497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14260__A2 _14264_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18323_ _18323_/A vssd1 vssd1 vccd1 vccd1 _19995_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15535_ _15243_/A _15075_/X _15534_/X _15093_/X vssd1 vssd1 vccd1 vccd1 _15535_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _18482_/Q _12556_/X _12557_/X vssd1 vssd1 vccd1 vccd1 _12747_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12746__S _12770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _18265_/A vssd1 vssd1 vccd1 vccd1 _18263_/S sky130_fd_sc_hd__buf_6
XFILLER_31_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12678_ _12679_/B _12679_/C _18782_/Q vssd1 vssd1 vccd1 vccd1 _12678_/Y sky130_fd_sc_hd__a21oi_1
X_15466_ _15365_/X _15228_/X _15465_/X _15400_/X vssd1 vssd1 vccd1 vccd1 _15466_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14246__B _14279_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17205_ _17205_/A vssd1 vssd1 vccd1 vccd1 _19524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11629_ _11629_/A vssd1 vssd1 vccd1 vccd1 _11629_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12023__A1 _12020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14417_ _14422_/C _14419_/C _14416_/Y vssd1 vssd1 vccd1 vccd1 _18700_/D sky130_fd_sc_hd__o21a_1
X_18185_ _17704_/X _19934_/Q _18191_/S vssd1 vssd1 vccd1 vccd1 _18186_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10034__A0 _19680_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15397_ _15397_/A _15397_/B vssd1 vssd1 vccd1 vccd1 _15397_/Y sky130_fd_sc_hd__nor2_1
X_17136_ _17135_/X _19501_/Q _17145_/S vssd1 vssd1 vccd1 vccd1 _17137_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14348_ _14350_/B _14350_/C _14347_/Y vssd1 vssd1 vccd1 vccd1 _18680_/D sky130_fd_sc_hd__o21a_1
XFILLER_7_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11886__A _14665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11209__S0 _11273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17067_ _17067_/A vssd1 vssd1 vccd1 vccd1 _19475_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10790__A _10843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14279_ _18655_/Q _14279_/B _14279_/C _14279_/D vssd1 vssd1 vccd1 vccd1 _14280_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__14262__A _14265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16018_ _13180_/X _19039_/Q _16020_/S vssd1 vssd1 vccd1 vccd1 _16019_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16888__S _16892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15276__A1 _12273_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _17969_/A vssd1 vssd1 vccd1 vccd1 _19852_/D sky130_fd_sc_hd__clkbuf_1
X_19708_ _19935_/CLK _19708_/D vssd1 vssd1 vccd1 vccd1 _19708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19639_ _19828_/CLK _19639_/D vssd1 vssd1 vccd1 vccd1 _19639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09323_ _09468_/A _17098_/A vssd1 vssd1 vccd1 vccd1 _09697_/B sky130_fd_sc_hd__or2_1
XFILLER_40_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09254_ _18990_/Q _18989_/Q _18991_/Q vssd1 vssd1 vccd1 vccd1 _11920_/B sky130_fd_sc_hd__or3b_1
XFILLER_21_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12014__A1 _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ _09283_/B _18966_/Q _09283_/D vssd1 vssd1 vccd1 vccd1 _09189_/A sky130_fd_sc_hd__or3_1
XFILLER_147_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14554__A3 _09341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10576__A1 _10223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11796__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09813__S0 _09898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17483__A _17483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10205__A _10208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_168_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13278__A0 _18852_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15715__B _15715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13516__A _13520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11980_ _14765_/A _14822_/B _14819_/A _11980_/D vssd1 vssd1 vccd1 vccd1 _12174_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10931_ _19201_/Q _19792_/Q _19954_/Q _19169_/Q _10776_/A _10662_/A vssd1 vssd1 vccd1
+ vccd1 _10932_/B sky130_fd_sc_hd__mux4_1
XFILLER_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17422__S _17424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10862_ _10009_/A _10859_/X _10861_/X vssd1 vssd1 vccd1 vccd1 _10862_/X sky130_fd_sc_hd__a21o_1
X_13650_ _13650_/A vssd1 vssd1 vccd1 vccd1 _13650_/X sky130_fd_sc_hd__clkbuf_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12601_ _12601_/A _12623_/C vssd1 vssd1 vccd1 vccd1 _12601_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _13580_/A _13580_/C _13110_/A vssd1 vssd1 vccd1 vccd1 _13582_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__16038__S _16042_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10793_ _10793_/A vssd1 vssd1 vccd1 vccd1 _10793_/X sky130_fd_sc_hd__buf_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12532_ _18776_/Q _18775_/Q _12532_/C vssd1 vssd1 vccd1 vccd1 _12582_/C sky130_fd_sc_hd__and3_2
X_15320_ _15284_/X _15316_/Y _15319_/X _15268_/X vssd1 vssd1 vccd1 vccd1 _15323_/B
+ sky130_fd_sc_hd__a211o_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12463_ _12464_/A _14880_/A vssd1 vssd1 vccd1 vccd1 _12465_/A sky130_fd_sc_hd__and2_1
XANTENNA__11439__S0 _11356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15251_ _15302_/A _15254_/A vssd1 vssd1 vccd1 vccd1 _15251_/X sky130_fd_sc_hd__or2_1
XFILLER_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ _11414_/A _11414_/B vssd1 vssd1 vccd1 vccd1 _11414_/Y sky130_fd_sc_hd__nor2_1
X_14202_ _18639_/Q _14200_/B _14201_/Y vssd1 vssd1 vccd1 vccd1 _18639_/D sky130_fd_sc_hd__o21a_1
X_15182_ _15178_/B _15177_/B _15180_/X _15181_/Y vssd1 vssd1 vccd1 vccd1 _15182_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12394_ _12448_/S _12390_/A _12393_/X _12012_/X vssd1 vssd1 vccd1 vccd1 _12394_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11764__B1 _13660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ _18617_/Q _14133_/B _14133_/C vssd1 vssd1 vccd1 vccd1 _14134_/C sky130_fd_sc_hd__and3_1
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ _18426_/Q _19455_/Q _19492_/Q _19066_/Q _11230_/X _11108_/A vssd1 vssd1 vccd1
+ vccd1 _11345_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19990_ _19990_/CLK _19990_/D vssd1 vssd1 vccd1 vccd1 _19990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14064_ _14088_/A _14064_/B _14064_/C vssd1 vssd1 vccd1 vccd1 _18596_/D sky130_fd_sc_hd__nor3_1
X_18941_ _18975_/CLK _18941_/D vssd1 vssd1 vccd1 vccd1 _18941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11276_ _11271_/Y _11274_/X _11275_/X _11278_/A vssd1 vssd1 vccd1 vccd1 _11276_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12314__B _12587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13015_ _18869_/Q _18870_/Q _13015_/C vssd1 vssd1 vccd1 vccd1 _13046_/C sky130_fd_sc_hd__and3_1
X_10227_ _19346_/Q _19617_/Q _19841_/Q _19585_/Q _10330_/S _10013_/A vssd1 vssd1 vccd1
+ vccd1 _10227_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18872_ _19001_/CLK _18872_/D vssd1 vssd1 vccd1 vccd1 _18872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17823_ _17880_/S vssd1 vssd1 vccd1 vccd1 _17832_/S sky130_fd_sc_hd__buf_2
X_10158_ _19219_/Q _19810_/Q _19972_/Q _19187_/Q _10328_/S _10027_/A vssd1 vssd1 vccd1
+ vccd1 _10158_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17754_ _17656_/X _19757_/Q _17760_/S vssd1 vssd1 vccd1 vccd1 _17755_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10089_ _19216_/Q _19807_/Q _19969_/Q _19184_/Q _10095_/S _10028_/X vssd1 vssd1 vccd1
+ vccd1 _10089_/X sky130_fd_sc_hd__mux4_1
X_14966_ _14966_/A _14990_/C vssd1 vssd1 vccd1 vccd1 _15007_/B sky130_fd_sc_hd__nor2_1
XFILLER_94_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16705_ _16762_/S vssd1 vssd1 vccd1 vccd1 _16714_/S sky130_fd_sc_hd__buf_2
XFILLER_48_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13917_ _18599_/Q _18598_/Q _18600_/Q _14065_/A vssd1 vssd1 vccd1 vccd1 _14073_/A
+ sky130_fd_sc_hd__and4_1
X_17685_ _17717_/A vssd1 vssd1 vccd1 vccd1 _17698_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_75_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14897_ _15100_/B _12738_/A _14933_/S vssd1 vssd1 vccd1 vccd1 _14897_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19424_ _20013_/CLK _19424_/D vssd1 vssd1 vccd1 vccd1 _19424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16636_ _16636_/A vssd1 vssd1 vccd1 vccd1 _19294_/D sky130_fd_sc_hd__clkbuf_1
X_13848_ _17084_/A vssd1 vssd1 vccd1 vccd1 _13848_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15430__A1 _12551_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19355_ _19981_/CLK _19355_/D vssd1 vssd1 vccd1 vccd1 _19355_/Q sky130_fd_sc_hd__dfxtp_1
X_16567_ _19264_/Q _13784_/X _16569_/S vssd1 vssd1 vccd1 vccd1 _16568_/A sky130_fd_sc_hd__mux2_1
X_13779_ _18492_/Q _13778_/X _13788_/S vssd1 vssd1 vccd1 vccd1 _13780_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13161__A _17675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18306_ _18306_/A vssd1 vssd1 vccd1 vccd1 _19987_/D sky130_fd_sc_hd__clkbuf_1
X_15518_ _15101_/X _15520_/B _14994_/X _15517_/X vssd1 vssd1 vccd1 vccd1 _15518_/X
+ sky130_fd_sc_hd__o211a_1
X_19286_ _19877_/CLK _19286_/D vssd1 vssd1 vccd1 vccd1 _19286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16498_ _16498_/A vssd1 vssd1 vccd1 vccd1 _19233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18237_ _19957_/Q _17675_/A _18241_/S vssd1 vssd1 vccd1 vccd1 _18238_/A sky130_fd_sc_hd__mux2_1
X_15449_ _15449_/A _15449_/B vssd1 vssd1 vccd1 vccd1 _15449_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18163__S _18169_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09948__B1 _09837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18168_ _18168_/A vssd1 vssd1 vccd1 vccd1 _19926_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17119_ _17656_/A vssd1 vssd1 vccd1 vccd1 _17119_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10724__S _10724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18099_ _18097_/X _19901_/Q _18112_/S vssd1 vssd1 vccd1 vccd1 _18100_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09941_ _19220_/Q _19811_/Q _19973_/Q _19188_/Q _09939_/X _09940_/X vssd1 vssd1 vccd1
+ vccd1 _09942_/B sky130_fd_sc_hd__mux4_1
XFILLER_132_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11507__B1 _09882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15816__A _15875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10405__S1 _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__A _10037_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _09872_/A vssd1 vssd1 vccd1 vccd1 _09873_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16411__S _16413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09814__A _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18338__S _18346_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11268__A2_N _09537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15270__B _15270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13432__B1 _12944_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _09306_/A _09480_/A _09306_/C vssd1 vssd1 vccd1 vccd1 _12290_/B sky130_fd_sc_hd__or3_2
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10341__S0 _10166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _09311_/A _09514_/A _09276_/C vssd1 vssd1 vccd1 vccd1 _09499_/B sky130_fd_sc_hd__or3_2
XANTENNA__14317__D _14317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_94_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _09306_/A vssd1 vssd1 vccd1 vccd1 _11961_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10644__S1 _10626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11130_ _19134_/Q _19395_/Q _19294_/Q _19629_/Q _11270_/S _10996_/A vssd1 vssd1 vccd1
+ vccd1 _11131_/B sky130_fd_sc_hd__mux4_1
XFILLER_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12134__B _12134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15726__A _17098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _11325_/A vssd1 vssd1 vccd1 vccd1 _11421_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16321__S _16330_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10012_ _10153_/A vssd1 vssd1 vccd1 vccd1 _10013_/A sky130_fd_sc_hd__buf_2
XFILLER_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09724__A _10859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15445__B _15449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14820_ _09522_/A _12859_/A _09272_/C _14782_/C _14819_/Y vssd1 vssd1 vccd1 vccd1
+ _14821_/B sky130_fd_sc_hd__a311o_1
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15660__A1 _12340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input15_A io_dbus_rdata[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14751_ _09516_/A _09516_/B _12833_/A _11931_/C vssd1 vssd1 vccd1 vccd1 _14808_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11963_ _11960_/Y _18898_/Q _12039_/A vssd1 vssd1 vccd1 vccd1 _14901_/A sky130_fd_sc_hd__mux2_2
XFILLER_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18248__S _18252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17152__S _17161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13702_ _19019_/Q _13702_/B vssd1 vssd1 vccd1 vccd1 _13702_/X sky130_fd_sc_hd__or2_1
X_17470_ _17160_/X _19642_/Q _17470_/S vssd1 vssd1 vccd1 vccd1 _17471_/A sky130_fd_sc_hd__mux2_1
X_10914_ _09775_/A _10905_/X _10909_/X _10913_/X _09819_/A vssd1 vssd1 vccd1 vccd1
+ _10914_/X sky130_fd_sc_hd__a311o_1
XFILLER_60_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14682_ _14682_/A vssd1 vssd1 vccd1 vccd1 _18793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11894_ _18574_/Q _13189_/A _11776_/X _18738_/Q vssd1 vssd1 vccd1 vccd1 _11894_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16421_ _16421_/A vssd1 vssd1 vccd1 vccd1 _19199_/D sky130_fd_sc_hd__clkbuf_1
X_10845_ _10211_/A _10844_/X _09775_/A vssd1 vssd1 vccd1 vccd1 _10845_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13633_ _13629_/X _13632_/Y _13689_/S vssd1 vssd1 vccd1 vccd1 _13633_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15963__A2 _15951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10237__B1 _09798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19140_ _19636_/CLK _19140_/D vssd1 vssd1 vccd1 vccd1 _19140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16352_ _17688_/A vssd1 vssd1 vccd1 vccd1 _16352_/X sky130_fd_sc_hd__clkbuf_2
X_10776_ _10776_/A vssd1 vssd1 vccd1 vccd1 _10776_/X sky130_fd_sc_hd__clkbuf_4
X_13564_ _18872_/Q _13565_/B vssd1 vssd1 vccd1 vccd1 _13580_/C sky130_fd_sc_hd__or2_4
XANTENNA__10332__S0 _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15303_ _15286_/X _15306_/B _15287_/X _15302_/X vssd1 vssd1 vccd1 vccd1 _15303_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19071_ _19693_/CLK _19071_/D vssd1 vssd1 vccd1 vccd1 _19071_/Q sky130_fd_sc_hd__dfxtp_1
X_12515_ _12515_/A _12515_/B vssd1 vssd1 vccd1 vccd1 _12516_/B sky130_fd_sc_hd__nand2_2
X_16283_ _13385_/X _19153_/Q _16291_/S vssd1 vssd1 vccd1 vccd1 _16284_/A sky130_fd_sc_hd__mux2_1
X_13495_ _18581_/Q _12877_/X _13490_/X _13492_/X _13494_/X vssd1 vssd1 vccd1 vccd1
+ _13495_/X sky130_fd_sc_hd__a2111o_4
XANTENNA__10883__S1 _10596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18022_ _19877_/Q _17090_/X _18024_/S vssd1 vssd1 vccd1 vccd1 _18023_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15234_ _15234_/A _15234_/B vssd1 vssd1 vccd1 vccd1 _15234_/Y sky130_fd_sc_hd__nor2_1
X_12446_ _12446_/A _12446_/B vssd1 vssd1 vccd1 vccd1 _12501_/C sky130_fd_sc_hd__and2_1
XANTENNA__18114__A0 _18858_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11737__B1 _11733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15165_ _15012_/X _15024_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _15165_/X sky130_fd_sc_hd__mux2_1
X_12377_ _12377_/A _12377_/B vssd1 vssd1 vccd1 vccd1 _12378_/A sky130_fd_sc_hd__and2_4
XANTENNA__15479__B2 _12645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output83_A _12551_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _11328_/A vssd1 vssd1 vccd1 vccd1 _11328_/X sky130_fd_sc_hd__clkbuf_4
X_14116_ _18727_/Q _18729_/Q _18728_/Q _14480_/A vssd1 vssd1 vccd1 vccd1 _14488_/A
+ sky130_fd_sc_hd__and4_1
X_19973_ _19973_/CLK _19973_/D vssd1 vssd1 vccd1 vccd1 _19973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15096_ _14922_/S _15095_/X _14984_/X vssd1 vssd1 vccd1 vccd1 _15096_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13855__S _13858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18924_ _18924_/CLK _18924_/D vssd1 vssd1 vccd1 vccd1 _18924_/Q sky130_fd_sc_hd__dfxtp_1
X_14047_ _18591_/Q _14044_/B _14046_/Y vssd1 vssd1 vccd1 vccd1 _18591_/D sky130_fd_sc_hd__o21a_1
X_11259_ _19357_/Q _19692_/Q _11270_/S vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18855_ _19010_/CLK _18855_/D vssd1 vssd1 vccd1 vccd1 _18855_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17806_ _17732_/X _19781_/Q _17808_/S vssd1 vssd1 vccd1 vccd1 _17807_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12060__A _12060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18786_ _18819_/CLK _18786_/D vssd1 vssd1 vccd1 vccd1 _18786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15998_ _13002_/X _19030_/Q _15998_/S vssd1 vssd1 vccd1 vccd1 _15999_/A sky130_fd_sc_hd__mux2_1
X_17737_ _17737_/A vssd1 vssd1 vccd1 vccd1 _19750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_161_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _18762_/CLK sky130_fd_sc_hd__clkbuf_16
X_14949_ _14947_/X _14948_/X _15014_/S vssd1 vssd1 vccd1 vccd1 _14949_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18158__S _18158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10476__B1 _10382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17668_ _17668_/A vssd1 vssd1 vccd1 vccd1 _17668_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15403__A1 _12498_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19407_ _19995_/CLK _19407_/D vssd1 vssd1 vccd1 vccd1 _19407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16619_ _18208_/A _17426_/B vssd1 vssd1 vccd1 vccd1 _16676_/A sky130_fd_sc_hd__or2_2
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13414__B1 _12944_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17599_ _17599_/A vssd1 vssd1 vccd1 vccd1 _19702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19338_ _19865_/CLK _19338_/D vssd1 vssd1 vccd1 vccd1 _19338_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_116_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_176_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19025_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19269_ _20022_/CLK _19269_/D vssd1 vssd1 vccd1 vccd1 _19269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09809__A _09809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18105__A0 _18855_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13193__A2 _12889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11777__C _11777_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17237__S _17243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09924_ _09929_/A _09924_/B vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_114_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _18734_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15890__A1 _14750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15890__B2 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input7_A io_dbus_rdata[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _09855_/A vssd1 vssd1 vccd1 vccd1 _11532_/S sky130_fd_sc_hd__clkbuf_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15265__B _15270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _20039_/Q _19877_/Q _19286_/Q _19056_/Q _11553_/A _09768_/X vssd1 vssd1 vccd1
+ vccd1 _09786_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_129_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18928_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12456__A1 _11904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__C1 _09568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10630_ _10630_/A _10630_/B vssd1 vssd1 vccd1 vccd1 _10630_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10561_ _09849_/A _10551_/X _10560_/X _09539_/A _18850_/Q vssd1 vssd1 vccd1 vccd1
+ _15952_/C sky130_fd_sc_hd__a32o_4
X_12300_ _12272_/A _12272_/B _12299_/Y vssd1 vssd1 vccd1 vccd1 _12301_/B sky130_fd_sc_hd__a21bo_1
XFILLER_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17001__A _17001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13280_ input11/X _13231_/X _13234_/X vssd1 vssd1 vccd1 vccd1 _13280_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10492_ _10492_/A _10492_/B vssd1 vssd1 vccd1 vccd1 _10492_/X sky130_fd_sc_hd__and2_1
XFILLER_155_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ _12231_/A _12255_/C vssd1 vssd1 vccd1 vccd1 _12231_/X sky130_fd_sc_hd__or2_1
XFILLER_108_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12162_ _12162_/A _12162_/B vssd1 vssd1 vccd1 vccd1 _12167_/A sky130_fd_sc_hd__nor2_1
XFILLER_122_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11113_ _11164_/A _11103_/X _11109_/X _11112_/Y vssd1 vssd1 vccd1 vccd1 _11113_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_16970_ _16970_/A vssd1 vssd1 vccd1 vccd1 _19442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16051__S _16053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12093_ _12043_/B _12046_/B _12043_/A vssd1 vssd1 vccd1 vccd1 _12215_/B sky130_fd_sc_hd__o21bai_4
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09454__A _14749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ _11322_/A vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__clkbuf_4
X_15921_ _15982_/A vssd1 vssd1 vccd1 vccd1 _15921_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16986__S _16986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18640_ _18677_/CLK _18640_/D vssd1 vssd1 vccd1 vccd1 _18640_/Q sky130_fd_sc_hd__dfxtp_1
X_15852_ _15852_/A vssd1 vssd1 vccd1 vccd1 _18978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14803_ _15954_/A vssd1 vssd1 vccd1 vccd1 _14803_/X sky130_fd_sc_hd__buf_8
XFILLER_18_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13644__A0 _18471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18571_ _20005_/CLK _18571_/D vssd1 vssd1 vccd1 vccd1 _18571_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output121_A _12851_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15783_ _18960_/Q _15783_/B vssd1 vssd1 vccd1 vccd1 _15783_/X sky130_fd_sc_hd__or2_1
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12995_ _18869_/Q vssd1 vssd1 vccd1 vccd1 _13535_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17522_ _19667_/Q vssd1 vssd1 vccd1 vccd1 _17523_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14734_ _18817_/Q _13719_/X _14738_/S vssd1 vssd1 vccd1 vccd1 _14735_/A sky130_fd_sc_hd__mux2_1
X_11946_ _09282_/D _09198_/A _09190_/X vssd1 vssd1 vccd1 vccd1 _11947_/C sky130_fd_sc_hd__a21o_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_93_clock clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 _19939_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _17135_/X _19634_/Q _17459_/S vssd1 vssd1 vccd1 vccd1 _17454_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _14665_/A vssd1 vssd1 vccd1 vccd1 _15883_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _19017_/Q _11877_/B vssd1 vssd1 vccd1 vccd1 _11877_/X sky130_fd_sc_hd__or2_1
XFILLER_32_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16404_ _16472_/S vssd1 vssd1 vccd1 vccd1 _16413_/S sky130_fd_sc_hd__buf_2
XFILLER_60_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13616_ _13612_/X _13615_/Y _13623_/S vssd1 vssd1 vccd1 vccd1 _13616_/X sky130_fd_sc_hd__mux2_1
X_10828_ _19331_/Q _19602_/Q _19826_/Q _19570_/Q _10764_/S _09606_/A vssd1 vssd1 vccd1
+ vccd1 _10828_/X sky130_fd_sc_hd__mux4_1
X_17384_ _17384_/A vssd1 vssd1 vccd1 vccd1 _19603_/D sky130_fd_sc_hd__clkbuf_1
X_14596_ _14596_/A vssd1 vssd1 vccd1 vccd1 _18767_/D sky130_fd_sc_hd__clkbuf_1
X_19123_ _20006_/CLK _19123_/D vssd1 vssd1 vccd1 vccd1 _19123_/Q sky130_fd_sc_hd__dfxtp_1
X_16335_ _16335_/A vssd1 vssd1 vccd1 vccd1 _19170_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15149__B1 _15951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13547_ _13554_/A _13554_/C vssd1 vssd1 vccd1 vccd1 _13547_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ _10760_/A _12843_/A vssd1 vssd1 vccd1 vccd1 _10759_/X sky130_fd_sc_hd__and2_1
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09629__A _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19054_ _19587_/CLK _19054_/D vssd1 vssd1 vccd1 vccd1 _19054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16266_ _16266_/A vssd1 vssd1 vccd1 vccd1 _19145_/D sky130_fd_sc_hd__clkbuf_1
X_13478_ input24/X _13340_/X _13319_/X vssd1 vssd1 vccd1 vccd1 _13478_/X sky130_fd_sc_hd__a21o_1
X_18005_ _19869_/Q _17065_/X _18009_/S vssd1 vssd1 vccd1 vccd1 _18006_/A sky130_fd_sc_hd__mux2_1
X_15217_ _15209_/X _15210_/Y _15215_/X _15216_/X vssd1 vssd1 vccd1 vccd1 _15221_/B
+ sky130_fd_sc_hd__a211o_1
X_12429_ _12537_/A _12847_/B _12318_/B vssd1 vssd1 vccd1 vccd1 _12429_/Y sky130_fd_sc_hd__o21ai_1
X_16197_ _16208_/A vssd1 vssd1 vccd1 vccd1 _16206_/S sky130_fd_sc_hd__buf_6
XFILLER_127_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12383__A0 _10760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19985_/CLK sky130_fd_sc_hd__clkbuf_16
X_15148_ _15920_/A vssd1 vssd1 vccd1 vccd1 _15951_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19956_ _20020_/CLK _19956_/D vssd1 vssd1 vccd1 vccd1 _19956_/Q sky130_fd_sc_hd__dfxtp_1
X_15079_ _15286_/A vssd1 vssd1 vccd1 vccd1 _15082_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15872__A1 _09466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15872__B2 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18907_ _18911_/CLK _18907_/D vssd1 vssd1 vccd1 vccd1 _18907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _20020_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_42_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19887_ _19887_/CLK _19887_/D vssd1 vssd1 vccd1 vccd1 _19887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09640_ _19943_/Q _19557_/Q _20007_/Q _19126_/Q _09635_/X _09639_/X vssd1 vssd1 vccd1
+ vccd1 _09641_/B sky130_fd_sc_hd__mux4_1
XFILLER_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10303__A _10411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18838_ _19324_/CLK _18838_/D vssd1 vssd1 vccd1 vccd1 _18838_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09571_ _11278_/A vssd1 vssd1 vccd1 vccd1 _11001_/A sky130_fd_sc_hd__clkbuf_2
X_18769_ _18994_/CLK _18769_/D vssd1 vssd1 vccd1 vccd1 _18769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16197__A _16208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12989__A2 _11686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10449__S _10449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16136__S _16144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10973__A _10973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09539__A _09539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15312__B1 _15311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ _11558_/A _09904_/X _09906_/X _09809_/X vssd1 vssd1 vccd1 vccd1 _09908_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13508__B _13508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12677__A1 _12338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20027_ _20027_/CLK _20027_/D vssd1 vssd1 vccd1 vccd1 _20027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09838_ _09826_/X _09835_/X _09836_/X _09750_/A _09837_/X vssd1 vssd1 vccd1 vccd1
+ _09838_/X sky130_fd_sc_hd__o221a_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09769_ _18454_/Q _19483_/Q _19520_/Q _19094_/Q _09733_/X _09768_/X vssd1 vssd1 vccd1
+ vccd1 _09769_/X sky130_fd_sc_hd__mux4_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15091__A2 _15482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _18997_/Q _11798_/Y _11799_/Y _11831_/A vssd1 vssd1 vccd1 vccd1 _11801_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _15542_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _12784_/A sky130_fd_sc_hd__xnor2_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11731_ _13656_/A vssd1 vssd1 vccd1 vccd1 _11731_/X sky130_fd_sc_hd__buf_2
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _14450_/A _14450_/B _18716_/Q vssd1 vssd1 vccd1 vccd1 _14452_/B sky130_fd_sc_hd__and3_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11650_/X _14758_/B _11653_/X _11661_/X vssd1 vssd1 vccd1 vccd1 _12153_/B
+ sky130_fd_sc_hd__o211a_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _18576_/Q _13189_/X _13397_/X _13399_/X _13400_/X vssd1 vssd1 vccd1 vccd1
+ _13708_/B sky130_fd_sc_hd__a2111o_1
X_10613_ _09562_/A _10606_/Y _10608_/Y _10610_/Y _10612_/Y vssd1 vssd1 vccd1 vccd1
+ _10613_/X sky130_fd_sc_hd__o32a_1
X_11593_ _11624_/A _11592_/C _11592_/A vssd1 vssd1 vccd1 vccd1 _11594_/B sky130_fd_sc_hd__a21oi_1
X_14381_ _18690_/Q _18689_/Q _18688_/Q _14381_/D vssd1 vssd1 vccd1 vccd1 _14391_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16120_ _13263_/X _19082_/Q _16122_/S vssd1 vssd1 vccd1 vccd1 _16121_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10544_ _10822_/A _10543_/X _09987_/A vssd1 vssd1 vccd1 vccd1 _10544_/X sky130_fd_sc_hd__a21o_1
X_13332_ _18476_/Q _13511_/A _14672_/A _18812_/Q _13331_/X vssd1 vssd1 vccd1 vccd1
+ _13332_/X sky130_fd_sc_hd__a221o_2
XFILLER_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11698__B _11712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10094__S _10094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16051_ _13443_/X _19054_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16052_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14354__A1 _14355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13263_ _17694_/A vssd1 vssd1 vccd1 vccd1 _13263_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10475_ _19339_/Q _19610_/Q _19834_/Q _19578_/Q _10208_/A _10473_/A vssd1 vssd1 vccd1
+ vccd1 _10475_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18261__S _18263_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__A1 _09881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15002_ _15181_/A _15002_/B vssd1 vssd1 vccd1 vccd1 _15002_/Y sky130_fd_sc_hd__nand2_1
X_12214_ _12214_/A vssd1 vssd1 vccd1 vccd1 _12220_/A sky130_fd_sc_hd__clkinv_2
XFILLER_68_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13194_ _13194_/A vssd1 vssd1 vccd1 vccd1 _13194_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10915__A1 _09702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10915__B2 _18843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output169_A _12140_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19810_ _19810_/CLK _19810_/D vssd1 vssd1 vccd1 vccd1 _19810_/Q sky130_fd_sc_hd__dfxtp_1
X_12145_ _15178_/B _12145_/B vssd1 vssd1 vccd1 vccd1 _12183_/A sky130_fd_sc_hd__xor2_4
XFILLER_123_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16953_ _16345_/X _19435_/Q _16953_/S vssd1 vssd1 vccd1 vccd1 _16954_/A sky130_fd_sc_hd__mux2_1
X_19741_ _20031_/CLK _19741_/D vssd1 vssd1 vccd1 vccd1 _19741_/Q sky130_fd_sc_hd__dfxtp_1
X_12076_ _12076_/A _12076_/B vssd1 vssd1 vccd1 vccd1 _12077_/A sky130_fd_sc_hd__and2_2
XFILLER_104_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15904_ _15847_/A _11960_/Y _15946_/A vssd1 vssd1 vccd1 vccd1 _15904_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09533__A1 _14782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11027_ _11149_/A _11027_/B vssd1 vssd1 vccd1 vccd1 _11027_/Y sky130_fd_sc_hd__nor2_1
X_19672_ _19994_/CLK _19672_/D vssd1 vssd1 vccd1 vccd1 _19672_/Q sky130_fd_sc_hd__dfxtp_1
X_16884_ _16348_/X _19404_/Q _16892_/S vssd1 vssd1 vccd1 vccd1 _16885_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10123__A _10657_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18623_ _18655_/CLK _18623_/D vssd1 vssd1 vccd1 vccd1 _18623_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09912__A _09912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15835_ input37/X _15834_/X _11865_/A _15738_/A vssd1 vssd1 vccd1 vccd1 _15836_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11891__A2 _11845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18554_ _18693_/CLK _18554_/D vssd1 vssd1 vccd1 vccd1 _18554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _18952_/Q _15775_/B vssd1 vssd1 vccd1 vccd1 _15766_/X sky130_fd_sc_hd__or2_1
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12978_ _17646_/A vssd1 vssd1 vccd1 vccd1 _12978_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17505_/A vssd1 vssd1 vccd1 vccd1 _19658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14717_ _14717_/A vssd1 vssd1 vccd1 vccd1 _18809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13153__B _18845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11929_ _11903_/A _12823_/B _11928_/X vssd1 vssd1 vccd1 vccd1 _12078_/A sky130_fd_sc_hd__a21o_1
X_18485_ _18773_/CLK _18485_/D vssd1 vssd1 vccd1 vccd1 _18485_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15697_ _18925_/Q _12745_/A _15699_/S vssd1 vssd1 vccd1 vccd1 _15698_/A sky130_fd_sc_hd__mux2_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17340__S _17348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17436_ _17436_/A vssd1 vssd1 vccd1 vccd1 _19626_/D sky130_fd_sc_hd__clkbuf_1
X_14648_ _14648_/A vssd1 vssd1 vccd1 vccd1 _14663_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11889__A _12889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13396__A2 _12943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17367_ _17424_/S vssd1 vssd1 vccd1 vccd1 _17376_/S sky130_fd_sc_hd__buf_2
X_14579_ _14665_/A vssd1 vssd1 vccd1 vccd1 _14648_/A sky130_fd_sc_hd__buf_2
XFILLER_20_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15790__B1 _15789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14265__A _14265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19106_ _19633_/CLK _19106_/D vssd1 vssd1 vccd1 vccd1 _19106_/Q sky130_fd_sc_hd__dfxtp_1
X_16318_ _16316_/X _19165_/Q _16330_/S vssd1 vssd1 vccd1 vccd1 _16319_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17298_ _17119_/X _19565_/Q _17304_/S vssd1 vssd1 vccd1 vccd1 _17299_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19037_ _19637_/CLK _19037_/D vssd1 vssd1 vccd1 vccd1 _19037_/Q sky130_fd_sc_hd__dfxtp_1
X_16249_ _16295_/S vssd1 vssd1 vccd1 vccd1 _16258_/S sky130_fd_sc_hd__buf_2
XFILLER_146_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11159__A1 _11237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput102 _12246_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[9] sky130_fd_sc_hd__buf_2
XANTENNA__12356__B1 _12459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 _12842_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[13] sky130_fd_sc_hd__buf_2
Xoutput124 _12855_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[23] sky130_fd_sc_hd__buf_2
XFILLER_161_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput135 _12827_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[4] sky130_fd_sc_hd__buf_2
XFILLER_115_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput146 _12378_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[13] sky130_fd_sc_hd__buf_2
Xoutput157 _12631_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[23] sky130_fd_sc_hd__buf_2
XFILLER_115_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput168 _12114_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[4] sky130_fd_sc_hd__buf_2
XANTENNA__13609__A _19007_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19939_ _19939_/CLK _19939_/D vssd1 vssd1 vccd1 vccd1 _19939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13328__B _13359_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ _10886_/A vssd1 vssd1 vccd1 vccd1 _09624_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11882__A2 _14528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09554_ _10194_/A vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10517__S0 _10529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09485_ _12193_/A vssd1 vssd1 vccd1 vccd1 _12393_/A sky130_fd_sc_hd__buf_2
XANTENNA__18346__S _18346_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17250__S _17254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__S0 _11156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10907__S _10907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10208__A _10208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _10260_/A vssd1 vssd1 vccd1 vccd1 _10261_/A sky130_fd_sc_hd__buf_2
XFILLER_11_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12898__A1 _12875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13519__A _13689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _10191_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10191_/X sky130_fd_sc_hd__or2_1
XFILLER_132_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13311__A2 _11755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13950_ _18557_/Q _13946_/C _13949_/Y vssd1 vssd1 vccd1 vccd1 _18557_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09732__A _10094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ _13175_/A vssd1 vssd1 vccd1 vccd1 _12936_/A sky130_fd_sc_hd__clkbuf_2
X_13881_ _12287_/A _12287_/B _14447_/B vssd1 vssd1 vccd1 vccd1 _18528_/D sky130_fd_sc_hd__a21o_1
XANTENNA__11873__A2 _11772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ _13714_/A _18923_/Q _15622_/S vssd1 vssd1 vccd1 vccd1 _15621_/A sky130_fd_sc_hd__mux2_1
X_12832_ _15738_/A _09492_/A _12845_/A vssd1 vssd1 vccd1 vccd1 _12833_/A sky130_fd_sc_hd__o21a_4
XFILLER_36_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15551_/A vssd1 vssd1 vccd1 vccd1 _18863_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12786_/A _12763_/B vssd1 vssd1 vccd1 vccd1 _12765_/A sky130_fd_sc_hd__nor2_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14501_/A _14501_/C _18734_/Q vssd1 vssd1 vccd1 vccd1 _14503_/C sky130_fd_sc_hd__a21oi_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _19972_/Q _17723_/A _18274_/S vssd1 vssd1 vccd1 vccd1 _18271_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _18566_/Q _13054_/B _11713_/X vssd1 vssd1 vccd1 vccd1 _11714_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _15482_/A _15482_/B vssd1 vssd1 vccd1 vccd1 _15482_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12674_/A _12695_/C _18544_/Q vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__a21oi_1
XFILLER_14_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _17112_/X _19531_/Q _17221_/S vssd1 vssd1 vccd1 vccd1 _17222_/A sky130_fd_sc_hd__mux2_1
X_14433_ _18705_/Q _18704_/Q _14433_/C _14433_/D vssd1 vssd1 vccd1 vccd1 _14439_/C
+ sky130_fd_sc_hd__and4_1
X_11645_ _11645_/A _11645_/B _11645_/C vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__and3_1
XFILLER_30_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09677__S1 _09642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17152_ _17151_/X _19506_/Q _17161_/S vssd1 vssd1 vccd1 vccd1 _17153_/A sky130_fd_sc_hd__mux2_1
Xinput15 io_dbus_rdata[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_4
X_14364_ _14364_/A _14373_/D vssd1 vssd1 vccd1 vccd1 _14365_/C sky130_fd_sc_hd__and2_1
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11576_ _15982_/B _12866_/C vssd1 vssd1 vccd1 vccd1 _11657_/A sky130_fd_sc_hd__nor2_2
Xinput26 io_dbus_rdata[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_2
Xinput37 io_ibus_inst[12] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_8
XFILLER_167_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16103_ _13137_/X _19074_/Q _16111_/S vssd1 vssd1 vccd1 vccd1 _16104_/A sky130_fd_sc_hd__mux2_1
Xinput48 io_ibus_inst[22] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_4
Xinput59 io_ibus_inst[3] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_1
X_13315_ _18603_/Q _13120_/X _13312_/X _13313_/X _13314_/X vssd1 vssd1 vccd1 vccd1
+ _13675_/B sky130_fd_sc_hd__a2111o_1
X_10527_ _10572_/A _10527_/B vssd1 vssd1 vccd1 vccd1 _10527_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17083_ _17083_/A vssd1 vssd1 vccd1 vccd1 _19480_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16504__S _16508_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14295_ _14319_/A _14295_/B vssd1 vssd1 vccd1 vccd1 _14295_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14813__A _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16034_ _13302_/X _19046_/Q _16042_/S vssd1 vssd1 vccd1 vccd1 _16035_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10458_ _10458_/A _10458_/B vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__or2_1
XFILLER_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13246_ _12875_/X _18850_/Q _13245_/X vssd1 vssd1 vccd1 vccd1 _13246_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10389_ _10013_/A _10388_/X _10001_/A vssd1 vssd1 vccd1 vccd1 _10389_/X sky130_fd_sc_hd__a21o_1
XFILLER_123_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13177_ input5/X _13091_/X _13094_/X vssd1 vssd1 vccd1 vccd1 _13177_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15827__A1 _18971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15827__B2 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12128_ _18522_/Q _18523_/Q _12128_/C vssd1 vssd1 vccd1 vccd1 _12477_/C sky130_fd_sc_hd__and3_2
X_17985_ _19860_/Q _17036_/X _17987_/S vssd1 vssd1 vccd1 vccd1 _17986_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17335__S _17337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12059_ _12059_/A vssd1 vssd1 vccd1 vccd1 _12059_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19724_ _19982_/CLK _19724_/D vssd1 vssd1 vccd1 vccd1 _19724_/Q sky130_fd_sc_hd__dfxtp_1
X_16936_ _16320_/X _19427_/Q _16942_/S vssd1 vssd1 vccd1 vccd1 _16937_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11313__A1 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10747__S0 _09725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09642__A _09642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19655_ _19656_/CLK _19655_/D vssd1 vssd1 vccd1 vccd1 _19655_/Q sky130_fd_sc_hd__dfxtp_1
X_16867_ _16867_/A vssd1 vssd1 vccd1 vccd1 _19396_/D sky130_fd_sc_hd__clkbuf_1
X_18606_ _19941_/CLK _18606_/D vssd1 vssd1 vccd1 vccd1 _18606_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15818_ _15831_/A _15818_/B vssd1 vssd1 vccd1 vccd1 _15819_/A sky130_fd_sc_hd__and2_1
X_19586_ _19972_/CLK _19586_/D vssd1 vssd1 vccd1 vccd1 _19586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16798_ _16798_/A vssd1 vssd1 vccd1 vccd1 _19366_/D sky130_fd_sc_hd__clkbuf_1
X_18537_ _18548_/CLK _18537_/D vssd1 vssd1 vccd1 vccd1 _18537_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15749_ _15847_/A _15734_/X _15748_/X _15743_/X vssd1 vssd1 vccd1 vccd1 _18945_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10300__B _12855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09270_ _11663_/A _14755_/A _09520_/B vssd1 vssd1 vccd1 vccd1 _11948_/B sky130_fd_sc_hd__nor3_2
X_18468_ _18994_/CLK _18468_/D vssd1 vssd1 vccd1 vccd1 _18468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17419_ _17419_/A vssd1 vssd1 vccd1 vccd1 _19619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13611__B _19007_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18399_ _17700_/X _20029_/Q _18407_/S vssd1 vssd1 vccd1 vccd1 _18400_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12508__A _12508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10028__A _10329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09817__A _09817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17268__A0 _17179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16491__A1 _13778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10738__S0 _09725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09552__A _10668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17440__A0 _17115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09606_ _09606_/A vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__14254__B1 _18653_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ _09537_/A vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11163__S0 _11293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10815__B1 _09912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09468_ _09468_/A vssd1 vssd1 vccd1 vccd1 _14749_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_145_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12280__A2 _12273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14557__A1 _14554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09399_ _09399_/A vssd1 vssd1 vccd1 vccd1 _11697_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14336__C _18674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ _19913_/Q _19527_/Q _19977_/Q _19096_/Q _11356_/X _11357_/X vssd1 vssd1 vccd1
+ vccd1 _11431_/B sky130_fd_sc_hd__mux4_1
XFILLER_138_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11361_ _11351_/X _11353_/X _11360_/X _09817_/A vssd1 vssd1 vccd1 vccd1 _11361_/Y
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__11041__B _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15729__A _16298_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16324__S _16330_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ _10312_/A _10312_/B vssd1 vssd1 vccd1 vccd1 _10312_/Y sky130_fd_sc_hd__nor2_1
X_13100_ _13100_/A vssd1 vssd1 vccd1 vccd1 _18432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14080_ _14088_/A _14080_/B _14080_/C vssd1 vssd1 vccd1 vccd1 _18602_/D sky130_fd_sc_hd__nor3_1
X_11292_ _18836_/Q _09536_/A _11281_/X _11291_/Y vssd1 vssd1 vccd1 vccd1 _11292_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_152_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13249__A _17049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10243_ _10246_/B _10242_/X vssd1 vssd1 vccd1 vccd1 _11647_/A sky130_fd_sc_hd__or2b_1
X_13031_ _18796_/Q _11841_/A _11817_/X _18763_/Q _13030_/X vssd1 vssd1 vccd1 vccd1
+ _13031_/X sky130_fd_sc_hd__a221o_1
XFILLER_65_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15809__B2 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A io_ibus_inst[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ _10162_/X _10165_/X _10169_/X _10173_/X _09822_/A vssd1 vssd1 vccd1 vccd1
+ _10174_/X sky130_fd_sc_hd__a311o_1
XFILLER_152_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17155__S _17161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17770_ _17770_/A vssd1 vssd1 vccd1 vccd1 _19764_/D sky130_fd_sc_hd__clkbuf_1
X_14982_ _14979_/X _14980_/X _15132_/S vssd1 vssd1 vccd1 vccd1 _14982_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_89_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16721_ _19332_/Q _13797_/X _16725_/S vssd1 vssd1 vccd1 vccd1 _16722_/A sky130_fd_sc_hd__mux2_1
X_13933_ _13936_/B _13936_/C _11884_/X vssd1 vssd1 vccd1 vccd1 _13933_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17431__A0 _17103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19440_ _19996_/CLK _19440_/D vssd1 vssd1 vccd1 vccd1 _19440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16652_ _16345_/X _19302_/Q _16652_/S vssd1 vssd1 vccd1 vccd1 _16653_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13864_ _14577_/A _13864_/B vssd1 vssd1 vccd1 vccd1 _13865_/A sky130_fd_sc_hd__and2_1
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15603_ _13256_/B _18915_/Q _15611_/S vssd1 vssd1 vccd1 vccd1 _15604_/A sky130_fd_sc_hd__mux2_1
X_19371_ _19706_/CLK _19371_/D vssd1 vssd1 vccd1 vccd1 _19371_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14796__A1 _12866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ _18485_/Q _12010_/X _12530_/A vssd1 vssd1 vccd1 vccd1 _12815_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16583_ _19271_/Q _13806_/X _16591_/S vssd1 vssd1 vccd1 vccd1 _16584_/A sky130_fd_sc_hd__mux2_1
X_13795_ _18497_/Q _13794_/X _13804_/S vssd1 vssd1 vccd1 vccd1 _13796_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18322_ _17694_/X _19995_/Q _18324_/S vssd1 vssd1 vccd1 vccd1 _18323_/A sky130_fd_sc_hd__mux2_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _15071_/X _15069_/X _15533_/X vssd1 vssd1 vccd1 vccd1 _15534_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12746_ _12743_/A _12745_/Y _12770_/S vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__mux2_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _18253_/A vssd1 vssd1 vccd1 vccd1 _19964_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13431__B _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15465_ _15522_/A _15465_/B _15465_/C vssd1 vssd1 vccd1 vccd1 _15465_/X sky130_fd_sc_hd__and3_1
X_12677_ _12338_/A _12675_/X _12676_/Y vssd1 vssd1 vccd1 vccd1 _12677_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17204_ _17208_/A _17204_/B vssd1 vssd1 vccd1 vccd1 _17205_/A sky130_fd_sc_hd__and2_1
XANTENNA__11232__A _11344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14416_ _14422_/C _14419_/C _14366_/X vssd1 vssd1 vccd1 vccd1 _14416_/Y sky130_fd_sc_hd__a21oi_1
X_18184_ _18184_/A vssd1 vssd1 vccd1 vccd1 _19933_/D sky130_fd_sc_hd__clkbuf_1
X_11628_ _11628_/A _11628_/B _11628_/C _11628_/D vssd1 vssd1 vccd1 vccd1 _11631_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15396_ _15366_/X _15392_/Y _15395_/X _15353_/X vssd1 vssd1 vccd1 vccd1 _15399_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12047__B _12583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17135_ _17672_/A vssd1 vssd1 vccd1 vccd1 _17135_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13858__S _13858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14347_ _14350_/B _14350_/C _14332_/X vssd1 vssd1 vccd1 vccd1 _14347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11559_ _19223_/Q _19814_/Q _19976_/Q _19191_/Q _11553_/X _11565_/A vssd1 vssd1 vccd1
+ vccd1 _11559_/X sky130_fd_sc_hd__mux4_2
XANTENNA__16234__S _16236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17066_ _19475_/Q _17065_/X _17072_/S vssd1 vssd1 vccd1 vccd1 _17067_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09637__A _09637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14278_ _18653_/Q _14278_/B _18651_/Q _14278_/D vssd1 vssd1 vccd1 vccd1 _14279_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__11209__S1 _11208_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16017_ _16017_/A vssd1 vssd1 vccd1 vccd1 _19038_/D sky130_fd_sc_hd__clkbuf_1
X_13229_ _13458_/A _11714_/Y _13227_/Y _13228_/Y _13307_/A vssd1 vssd1 vccd1 vccd1
+ _13229_/X sky130_fd_sc_hd__a311o_1
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _19852_/Q _17010_/X _17976_/S vssd1 vssd1 vccd1 vccd1 _17969_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09372__A _18952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19707_ _19996_/CLK _19707_/D vssd1 vssd1 vccd1 vccd1 _19707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11298__B1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16919_ _16919_/A vssd1 vssd1 vccd1 vccd1 _19420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17899_ _17899_/A vssd1 vssd1 vccd1 vccd1 _19821_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11393__S0 _11154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19638_ _19767_/CLK _19638_/D vssd1 vssd1 vccd1 vccd1 _19638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19569_ _19569_/CLK _19569_/D vssd1 vssd1 vccd1 vccd1 _19569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16409__S _16413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ _09322_/A vssd1 vssd1 vccd1 vccd1 _17098_/A sky130_fd_sc_hd__buf_4
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09253_ _18992_/Q _09284_/A _09282_/B _11951_/B vssd1 vssd1 vccd1 vccd1 _09502_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA__16933__A _16990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09184_ _09282_/B vssd1 vssd1 vccd1 vccd1 _09313_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12014__A2 _12012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15549__A _15602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16144__S _16144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10981__A _11270_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12970__B1 _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09547__A _09547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09813__S1 _09895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15267__A2 _15270_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_90_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11289__B1 _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10930_ _09560_/A _10927_/Y _10929_/Y _09873_/A vssd1 vssd1 vccd1 vccd1 _10930_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_29_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10861_ _09830_/A _10860_/X _11493_/A vssd1 vssd1 vccd1 vccd1 _10861_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15975__B1 _15955_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13532__A _13660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ _18540_/Q vssd1 vssd1 vccd1 vccd1 _12601_/A sky130_fd_sc_hd__buf_2
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17004__A _17004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13580_ _13580_/A _18874_/Q _13580_/C vssd1 vssd1 vccd1 vccd1 _13593_/B sky130_fd_sc_hd__or3_1
X_10792_ _10905_/A vssd1 vssd1 vccd1 vccd1 _10858_/A sky130_fd_sc_hd__clkbuf_2
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12531_ _12508_/A _12532_/C _18776_/Q vssd1 vssd1 vccd1 vccd1 _12531_/Y sky130_fd_sc_hd__a21oi_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16843__A _17203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15250_ _15254_/A _15254_/B vssd1 vssd1 vccd1 vccd1 _15250_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12462_ _15952_/C _18914_/Q _12517_/S vssd1 vssd1 vccd1 vccd1 _14880_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11439__S1 _11357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14201_ _14239_/A _14207_/C vssd1 vssd1 vccd1 vccd1 _14201_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11413_ _19655_/Q _19421_/Q _18486_/Q _19751_/Q _11328_/X _11073_/A vssd1 vssd1 vccd1
+ vccd1 _11414_/B sky130_fd_sc_hd__mux4_1
X_15181_ _15181_/A _15181_/B vssd1 vssd1 vccd1 vccd1 _15181_/Y sky130_fd_sc_hd__nand2_1
X_12393_ _12393_/A _12393_/B _12393_/C _12393_/D vssd1 vssd1 vccd1 vccd1 _12393_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_126_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _14133_/B _14133_/C _18617_/Q vssd1 vssd1 vccd1 vccd1 _14134_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12961__B1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11344_ _11344_/A _11344_/B vssd1 vssd1 vccd1 vccd1 _11344_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11198__S _11367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14063_ _14062_/A _14062_/C _18596_/Q vssd1 vssd1 vccd1 vccd1 _14064_/C sky130_fd_sc_hd__a21oi_1
X_18940_ _18975_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _18940_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_165_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11275_ _19658_/Q _19424_/Q _18489_/Q _19754_/Q _11049_/S _10973_/A vssd1 vssd1 vccd1
+ vccd1 _11275_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13014_ _18838_/Q _13542_/B _13215_/S vssd1 vssd1 vccd1 vccd1 _13014_/X sky130_fd_sc_hd__mux2_1
X_10226_ _10388_/S vssd1 vssd1 vccd1 vccd1 _10330_/S sky130_fd_sc_hd__buf_2
XANTENNA_output151_A _12510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18871_ _19001_/CLK _18871_/D vssd1 vssd1 vccd1 vccd1 _18871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10157_ _10434_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _10157_/X sky130_fd_sc_hd__or2_1
X_17822_ _17822_/A vssd1 vssd1 vccd1 vccd1 _19787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10088_ _10093_/A _10088_/B vssd1 vssd1 vccd1 vccd1 _10088_/Y sky130_fd_sc_hd__nor2_1
X_17753_ _17753_/A vssd1 vssd1 vccd1 vccd1 _19756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14965_ _14965_/A _15243_/A vssd1 vssd1 vccd1 vccd1 _14965_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17613__S _17617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__A _11227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13916_ _18595_/Q _18597_/Q _18596_/Q _14056_/A vssd1 vssd1 vccd1 vccd1 _14065_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16704_ _16704_/A vssd1 vssd1 vccd1 vccd1 _19324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15922__A _15946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17684_ _17684_/A vssd1 vssd1 vccd1 vccd1 _17684_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14896_ _14927_/A vssd1 vssd1 vccd1 vccd1 _14933_/S sky130_fd_sc_hd__clkbuf_2
X_19423_ _20012_/CLK _19423_/D vssd1 vssd1 vccd1 vccd1 _19423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16635_ _16320_/X _19294_/Q _16641_/S vssd1 vssd1 vccd1 vccd1 _16636_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _13847_/A vssd1 vssd1 vccd1 vccd1 _18513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11127__S0 _11258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19354_ _19979_/CLK _19354_/D vssd1 vssd1 vccd1 vccd1 _19354_/Q sky130_fd_sc_hd__dfxtp_1
X_16566_ _16566_/A vssd1 vssd1 vccd1 vccd1 _19263_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13441__A1 _13223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13778_ _17014_/A vssd1 vssd1 vccd1 vccd1 _13778_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10255__A1 _09597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18305_ _17668_/X _19987_/Q _18313_/S vssd1 vssd1 vccd1 vccd1 _18306_/A sky130_fd_sc_hd__mux2_1
X_15517_ _15517_/A _15520_/A vssd1 vssd1 vccd1 vccd1 _15517_/X sky130_fd_sc_hd__or2_1
XANTENNA__10277__S _10277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19285_ _19876_/CLK _19285_/D vssd1 vssd1 vccd1 vccd1 _19285_/Q sky130_fd_sc_hd__dfxtp_1
X_12729_ _12729_/A _12729_/B _12729_/C vssd1 vssd1 vccd1 vccd1 _12729_/X sky130_fd_sc_hd__and3_1
X_16497_ _19233_/Q _13787_/X _16497_/S vssd1 vssd1 vccd1 vccd1 _16498_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12058__A _18457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18236_ _18236_/A vssd1 vssd1 vccd1 vccd1 _19956_/D sky130_fd_sc_hd__clkbuf_1
X_15448_ _15366_/X _15445_/Y _15447_/X _15353_/X vssd1 vssd1 vccd1 vccd1 _15451_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18167_ _17678_/X _19926_/Q _18169_/S vssd1 vssd1 vccd1 vccd1 _18168_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15379_ _18849_/Q _15363_/X _15378_/X vssd1 vssd1 vccd1 vccd1 _18849_/D sky130_fd_sc_hd__o21a_1
XFILLER_128_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17118_ _17118_/A vssd1 vssd1 vccd1 vccd1 _19495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18098_ _18115_/A vssd1 vssd1 vccd1 vccd1 _18112_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__16899__S _16903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17049_ _17049_/A vssd1 vssd1 vccd1 vccd1 _17049_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09940_ _09940_/A vssd1 vssd1 vccd1 vccd1 _09940_/X sky130_fd_sc_hd__buf_2
XFILLER_104_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11507__B2 _11506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12704__B1 _12860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _19526_/Q vssd1 vssd1 vccd1 vccd1 _09872_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_112_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10494__A1 _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09830__A _09830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15957__B1 _15955_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10976__A _11409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09305_ _11941_/A _09233_/Y _09292_/X _09535_/B vssd1 vssd1 vccd1 vccd1 _09305_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10341__S1 _10223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_37_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ _18991_/Q _18988_/Q _18987_/Q _18986_/Q vssd1 vssd1 vccd1 vccd1 _09276_/C
+ sky130_fd_sc_hd__or4_2
XANTENNA__13196__B1 _13192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15279__A _15458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09167_ _09282_/B vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16602__S _16602_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13499__A1 _12874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11060_ _09560_/A _11047_/X _11051_/X _11059_/X _11133_/A vssd1 vssd1 vccd1 vccd1
+ _11060_/X sky130_fd_sc_hd__a311o_2
XFILLER_135_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15726__B _15732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10011_ _10011_/A vssd1 vssd1 vccd1 vccd1 _10153_/A sky130_fd_sc_hd__buf_2
XFILLER_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12171__B2 _12170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12431__A _12514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14750_ _14750_/A _14750_/B _09471_/C vssd1 vssd1 vccd1 vccd1 _14750_/X sky130_fd_sc_hd__or3b_1
X_11962_ _09292_/X _11962_/B _14758_/A vssd1 vssd1 vccd1 vccd1 _12039_/A sky130_fd_sc_hd__and3b_2
XFILLER_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13701_ _13714_/C _13699_/Y _13700_/X vssd1 vssd1 vccd1 vccd1 _13701_/Y sky130_fd_sc_hd__a21oi_1
X_10913_ _10900_/A _10910_/X _10912_/X _09792_/A vssd1 vssd1 vccd1 vccd1 _10913_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09970__S0 _09657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14681_ _18793_/Q _11801_/A _14683_/S vssd1 vssd1 vccd1 vccd1 _14682_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16049__S _16053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ _18606_/Q _11851_/X _11852_/X _18638_/Q vssd1 vssd1 vccd1 vccd1 _11893_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13262__A _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16420_ _19199_/Q _13781_/X _16424_/S vssd1 vssd1 vccd1 vccd1 _16421_/A sky130_fd_sc_hd__mux2_1
X_13632_ _13637_/B _13632_/B vssd1 vssd1 vccd1 vccd1 _13632_/Y sky130_fd_sc_hd__nand2_2
X_10844_ _19924_/Q _19538_/Q _19988_/Q _19107_/Q _10859_/S _11487_/A vssd1 vssd1 vccd1
+ vccd1 _10844_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16351_ _16351_/A vssd1 vssd1 vccd1 vccd1 _19175_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17669__A _17736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13563_ _13563_/A vssd1 vssd1 vccd1 vccd1 _14548_/A sky130_fd_sc_hd__buf_2
XFILLER_12_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10775_ _10775_/A vssd1 vssd1 vccd1 vccd1 _10776_/A sky130_fd_sc_hd__buf_2
XFILLER_13_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10332__S1 _10283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11985__A1 _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ _15302_/A _15306_/A vssd1 vssd1 vccd1 vccd1 _15302_/X sky130_fd_sc_hd__or2_1
X_12514_ _12514_/A _12514_/B _15397_/A _12458_/A vssd1 vssd1 vccd1 vccd1 _12515_/B
+ sky130_fd_sc_hd__or4b_2
X_19070_ _20017_/CLK _19070_/D vssd1 vssd1 vccd1 vccd1 _19070_/Q sky130_fd_sc_hd__dfxtp_1
X_16282_ _16282_/A vssd1 vssd1 vccd1 vccd1 _16291_/S sky130_fd_sc_hd__buf_4
XFILLER_40_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13494_ _18677_/Q _11815_/X _12890_/X _14124_/B vssd1 vssd1 vccd1 vccd1 _13494_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18021_ _18021_/A vssd1 vssd1 vccd1 vccd1 _19876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15233_ _15209_/X _15230_/Y _15232_/X _15216_/X vssd1 vssd1 vccd1 vccd1 _15236_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12445_ _12446_/A _12446_/B vssd1 vssd1 vccd1 vccd1 _12447_/A sky130_fd_sc_hd__nor2_1
XFILLER_126_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15164_ _15546_/A vssd1 vssd1 vccd1 vccd1 _15478_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12376_ _13650_/A _12371_/X _12372_/X _12375_/Y vssd1 vssd1 vccd1 vccd1 _12377_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14115_ _18725_/Q _18724_/Q _18726_/Q _14471_/A vssd1 vssd1 vccd1 vccd1 _14480_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11327_ _09559_/A _11317_/X _11321_/X _11326_/X _09549_/A vssd1 vssd1 vccd1 vccd1
+ _11327_/X sky130_fd_sc_hd__a311o_1
XANTENNA__15917__A _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10126__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19972_ _19972_/CLK _19972_/D vssd1 vssd1 vccd1 vccd1 _19972_/Q sky130_fd_sc_hd__dfxtp_1
X_15095_ _14905_/X _14979_/X _15189_/S vssd1 vssd1 vccd1 vccd1 _15095_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output76_A _12390_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ _14046_/A _14051_/C vssd1 vssd1 vccd1 vccd1 _14046_/Y sky130_fd_sc_hd__nor2_1
X_18923_ _18923_/CLK _18923_/D vssd1 vssd1 vccd1 vccd1 _18923_/Q sky130_fd_sc_hd__dfxtp_1
X_11258_ _19229_/Q _19724_/Q _11258_/S vssd1 vssd1 vccd1 vccd1 _11258_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10209_ _19250_/Q _19745_/Q _10209_/S vssd1 vssd1 vccd1 vccd1 _10210_/B sky130_fd_sc_hd__mux2_1
X_18854_ _19025_/CLK _18854_/D vssd1 vssd1 vccd1 vccd1 _18854_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11189_ _11157_/A _11186_/X _11188_/X vssd1 vssd1 vccd1 vccd1 _11189_/Y sky130_fd_sc_hd__a21oi_1
X_17805_ _17805_/A vssd1 vssd1 vccd1 vccd1 _19780_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12060__B _12060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15997_ _15997_/A vssd1 vssd1 vccd1 vccd1 _19029_/D sky130_fd_sc_hd__clkbuf_1
X_18785_ _18819_/CLK _18785_/D vssd1 vssd1 vccd1 vccd1 _18785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17736_ _17735_/X _19750_/Q _17736_/S vssd1 vssd1 vccd1 vccd1 _17737_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14948_ _15474_/B _15219_/B _14948_/S vssd1 vssd1 vccd1 vccd1 _14948_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09866__B1 _09568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18050__A0 _18839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09650__A _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17667_ _17667_/A vssd1 vssd1 vccd1 vccd1 _19728_/D sky130_fd_sc_hd__clkbuf_1
X_14879_ _14879_/A vssd1 vssd1 vccd1 vccd1 _15338_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14268__A _14479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19406_ _19993_/CLK _19406_/D vssd1 vssd1 vccd1 vccd1 _19406_/Q sky130_fd_sc_hd__dfxtp_1
X_16618_ _16618_/A vssd1 vssd1 vccd1 vccd1 _19287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17598_ _17147_/X _19702_/Q _17606_/S vssd1 vssd1 vccd1 vccd1 _17599_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13414__A1 _18481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10228__A1 _10438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19337_ _20026_/CLK _19337_/D vssd1 vssd1 vccd1 vccd1 _19337_/Q sky130_fd_sc_hd__dfxtp_1
X_16549_ _16617_/S vssd1 vssd1 vccd1 vccd1 _16558_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__18174__S _18180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19268_ _20021_/CLK _19268_/D vssd1 vssd1 vccd1 vccd1 _19268_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15706__A3 _13700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18219_ _19949_/Q _17649_/A _18219_/S vssd1 vssd1 vccd1 vccd1 _18220_/A sky130_fd_sc_hd__mux2_1
X_19199_ _19949_/CLK _19199_/D vssd1 vssd1 vccd1 vccd1 _19199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18105__A1 _13685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16116__A0 _13238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10036__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16422__S _16424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09923_ _19156_/Q _19417_/Q _19316_/Q _19651_/Q _09659_/S _09647_/A vssd1 vssd1 vccd1
+ vccd1 _09924_/B sky130_fd_sc_hd__mux4_1
XFILLER_160_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11566__S _11566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10470__S _10470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09854_ _11533_/A _09853_/X _09933_/A vssd1 vssd1 vccd1 vccd1 _09854_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11361__C1 _09817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09785_ _09903_/A vssd1 vssd1 vccd1 vccd1 _11553_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11339__S0 _10618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12456__A2 _12848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09560__A _09560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13082__A _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13810__A _17046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10560_ _10553_/X _10555_/X _10557_/X _10559_/X _09875_/A vssd1 vssd1 vccd1 vccd1
+ _10560_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09219_ _09285_/C vssd1 vssd1 vccd1 vccd1 _09436_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_154_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10491_ _19370_/Q _19705_/Q _10493_/S vssd1 vssd1 vccd1 vccd1 _10492_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12230_ _18765_/Q vssd1 vssd1 vccd1 vccd1 _12231_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12161_ _18763_/Q _12161_/B vssd1 vssd1 vccd1 vccd1 _12162_/B sky130_fd_sc_hd__nor2_1
XFILLER_163_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11112_ _10854_/A _11110_/X _11227_/A vssd1 vssd1 vccd1 vccd1 _11112_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12092_ _12092_/A _12092_/B vssd1 vssd1 vccd1 vccd1 _12215_/A sky130_fd_sc_hd__nor2_2
XFILLER_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13257__A _13257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09454__B _09454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11043_ _19523_/Q vssd1 vssd1 vccd1 vccd1 _11322_/A sky130_fd_sc_hd__clkbuf_2
X_15920_ _15920_/A vssd1 vssd1 vccd1 vccd1 _15982_/A sky130_fd_sc_hd__buf_2
XANTENNA__10155__B1 _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12161__A _18763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13892__A1 _12501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13892__B2 _12484_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15851_ _15861_/A _17204_/B vssd1 vssd1 vccd1 vccd1 _15852_/A sky130_fd_sc_hd__and2_1
XFILLER_65_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18259__S _18263_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14802_ _15147_/A vssd1 vssd1 vccd1 vccd1 _15954_/A sky130_fd_sc_hd__buf_4
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18570_ _20005_/CLK _18570_/D vssd1 vssd1 vccd1 vccd1 _18570_/Q sky130_fd_sc_hd__dfxtp_1
X_15782_ _12260_/A _11867_/X _15781_/X _13885_/X vssd1 vssd1 vccd1 vccd1 _18959_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12994_ _18837_/Q _13529_/B _13215_/S vssd1 vssd1 vccd1 vccd1 _12994_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09470__A _18990_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17521_ _17521_/A vssd1 vssd1 vccd1 vccd1 _19666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14733_ _14733_/A vssd1 vssd1 vccd1 vccd1 _18816_/D sky130_fd_sc_hd__clkbuf_1
X_11945_ _11945_/A _12822_/B vssd1 vssd1 vccd1 vccd1 _11945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output114_A _12843_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14088__A _14088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17452_/A vssd1 vssd1 vccd1 vccd1 _19633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14664_ _14664_/A vssd1 vssd1 vccd1 vccd1 _18787_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11876_ _18573_/Q _11869_/Y _11873_/X _11875_/X vssd1 vssd1 vccd1 vccd1 _11877_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _16459_/A vssd1 vssd1 vccd1 vccd1 _16472_/S sky130_fd_sc_hd__buf_6
XANTENNA__10615__A1_N _18849_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13615_ _13630_/C _13615_/B vssd1 vssd1 vccd1 vccd1 _13615_/Y sky130_fd_sc_hd__nand2_2
X_10827_ _10832_/A _10827_/B vssd1 vssd1 vccd1 vccd1 _10827_/Y sky130_fd_sc_hd__nor2_1
X_17383_ _19603_/Q _17033_/X _17387_/S vssd1 vssd1 vccd1 vccd1 _17384_/A sky130_fd_sc_hd__mux2_1
X_14595_ _14595_/A _14595_/B vssd1 vssd1 vccd1 vccd1 _14596_/A sky130_fd_sc_hd__and2_1
XANTENNA__14816__A _14927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11958__A1 _11945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16346__A0 _16345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19122_ _19873_/CLK _19122_/D vssd1 vssd1 vccd1 vccd1 _19122_/Q sky130_fd_sc_hd__dfxtp_1
X_16334_ _16332_/X _19170_/Q _16346_/S vssd1 vssd1 vccd1 vccd1 _16335_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15149__A1 _12094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13546_ _13528_/X _13542_/X _13545_/Y _13532_/X _18999_/Q vssd1 vssd1 vccd1 vccd1
+ _13546_/X sky130_fd_sc_hd__a32o_4
X_10758_ _09882_/A _10746_/X _10757_/X _09912_/A _10735_/Y vssd1 vssd1 vccd1 vccd1
+ _12843_/A sky130_fd_sc_hd__o32a_4
XFILLER_119_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10091__C1 _09823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19053_ _20006_/CLK _19053_/D vssd1 vssd1 vccd1 vccd1 _19053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16265_ _13250_/X _19145_/Q _16269_/S vssd1 vssd1 vccd1 vccd1 _16266_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ _12897_/X _13486_/B _13476_/X _09532_/A vssd1 vssd1 vccd1 vccd1 _13477_/X
+ sky130_fd_sc_hd__a31o_1
X_10689_ _19239_/Q _19734_/Q _10691_/S vssd1 vssd1 vccd1 vccd1 _10690_/B sky130_fd_sc_hd__mux2_1
XFILLER_139_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18004_ _18004_/A vssd1 vssd1 vccd1 vccd1 _19868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12907__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15216_ _15268_/A vssd1 vssd1 vccd1 vccd1 _15216_/X sky130_fd_sc_hd__clkbuf_2
X_12428_ _12428_/A vssd1 vssd1 vccd1 vccd1 _14763_/C sky130_fd_sc_hd__buf_2
X_16196_ _16196_/A vssd1 vssd1 vccd1 vccd1 _19115_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12383__A1 _18911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15147_ _15147_/A vssd1 vssd1 vccd1 vccd1 _15920_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12359_ _12360_/A _14883_/A vssd1 vssd1 vccd1 vccd1 _12361_/A sky130_fd_sc_hd__and2_1
XANTENNA__12770__S _12770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10394__B1 _10382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19955_ _19957_/CLK _19955_/D vssd1 vssd1 vccd1 vccd1 _19955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15078_ _15165_/S _15078_/B vssd1 vssd1 vccd1 vccd1 _15078_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13332__B1 _14672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15872__A2 _15856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18906_ _19488_/CLK _18906_/D vssd1 vssd1 vccd1 vccd1 _18906_/Q sky130_fd_sc_hd__dfxtp_1
X_14029_ _14029_/A vssd1 vssd1 vccd1 vccd1 _14034_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_171_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19886_ _19888_/CLK _19886_/D vssd1 vssd1 vccd1 vccd1 _19886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18837_ _18972_/CLK _18837_/D vssd1 vssd1 vccd1 vccd1 _18837_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11894__B1 _11776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18169__S _18169_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09570_ _11325_/A vssd1 vssd1 vccd1 vccd1 _11278_/A sky130_fd_sc_hd__buf_2
XFILLER_82_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09839__B1 _11574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18768_ _19899_/CLK _18768_/D vssd1 vssd1 vccd1 vccd1 _18768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17719_ _17719_/A vssd1 vssd1 vccd1 vccd1 _19744_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09934__S0 _09668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18699_ _18744_/CLK _18699_/D vssd1 vssd1 vccd1 vccd1 _18699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14899__A0 _15078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15560__B2 _12812_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13776__S _13788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clock_A clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17248__S _17254_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14461__A _14495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19379__CLK _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__A _09555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15312__A1 _18845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09906_ _09957_/A _09906_/B vssd1 vssd1 vccd1 vccd1 _09906_/X sky130_fd_sc_hd__or2_1
XFILLER_99_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20026_ _20026_/CLK _20026_/D vssd1 vssd1 vccd1 vccd1 _20026_/Q sky130_fd_sc_hd__dfxtp_1
X_09837_ _09837_/A vssd1 vssd1 vccd1 vccd1 _09837_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09768_ _09824_/A vssd1 vssd1 vccd1 vccd1 _09768_/X sky130_fd_sc_hd__buf_2
XANTENNA__12429__A2 _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09925__S0 _09659_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09699_ _09699_/A vssd1 vssd1 vccd1 vccd1 _09699_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17711__S _17714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11730_ _11730_/A vssd1 vssd1 vccd1 vccd1 _13656_/A sky130_fd_sc_hd__buf_2
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15379__A1 _18849_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11667_/C _11656_/Y _11657_/Y _11660_/Y vssd1 vssd1 vccd1 vccd1 _11661_/X
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16327__S _16330_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ _18608_/Q _11851_/X _13194_/X _18740_/Q vssd1 vssd1 vccd1 vccd1 _13400_/X
+ sky130_fd_sc_hd__a22o_1
X_10612_ _10674_/A _10611_/X _09562_/A vssd1 vssd1 vccd1 vccd1 _10612_/Y sky130_fd_sc_hd__o21ai_1
X_14380_ _18690_/Q _14384_/C vssd1 vssd1 vccd1 vccd1 _14382_/B sky130_fd_sc_hd__nor2_1
X_11592_ _11592_/A _11624_/A _11592_/C vssd1 vssd1 vccd1 vccd1 _11594_/A sky130_fd_sc_hd__and3_1
XFILLER_10_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14355__B _14355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10612__A1 _10674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _19903_/Q _13373_/B _09405_/A _18700_/Q _11869_/Y vssd1 vssd1 vccd1 vccd1
+ _13331_/X sky130_fd_sc_hd__a221o_1
XFILLER_167_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10543_ _19241_/Q _19736_/Q _10543_/S vssd1 vssd1 vccd1 vccd1 _10543_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16050_ _16050_/A vssd1 vssd1 vccd1 vccd1 _19053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13262_ _17052_/A vssd1 vssd1 vccd1 vccd1 _17694_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10474_ _19147_/Q _19408_/Q _19307_/Q _19642_/Q _09729_/A _10473_/X vssd1 vssd1 vccd1
+ vccd1 _10474_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_160_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19063_/CLK sky130_fd_sc_hd__clkbuf_16
X_15001_ _15305_/A vssd1 vssd1 vccd1 vccd1 _15181_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17158__S _17161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12213_ _12213_/A _14871_/A vssd1 vssd1 vccd1 vccd1 _12214_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13562__B1 _13660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13193_ _18660_/Q _12889_/X _11852_/X _18628_/Q vssd1 vssd1 vccd1 vccd1 _13193_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09465__A _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ _12080_/B _12209_/C _12208_/A vssd1 vssd1 vccd1 vccd1 _12145_/B sky130_fd_sc_hd__o21ai_2
XFILLER_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_2_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13314__B1 _13082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19740_ _19868_/CLK _19740_/D vssd1 vssd1 vccd1 vccd1 _19740_/Q sky130_fd_sc_hd__dfxtp_1
X_16952_ _16952_/A vssd1 vssd1 vccd1 vccd1 _19434_/D sky130_fd_sc_hd__clkbuf_1
X_12075_ _13508_/A _12057_/X _12058_/X _12074_/X _12402_/B vssd1 vssd1 vccd1 vccd1
+ _12076_/B sky130_fd_sc_hd__a311o_1
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_6_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_175_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18878_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_159_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ _19136_/Q _19397_/Q _19296_/Q _19631_/Q _10962_/X _11022_/X vssd1 vssd1 vccd1
+ vccd1 _11027_/B sky130_fd_sc_hd__mux4_1
X_15903_ _15916_/A vssd1 vssd1 vccd1 vccd1 _15946_/A sky130_fd_sc_hd__clkbuf_4
X_19671_ _19767_/CLK _19671_/D vssd1 vssd1 vccd1 vccd1 _19671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11876__B1 _11873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16883_ _16905_/A vssd1 vssd1 vccd1 vccd1 _16892_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__16298__A _16691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18622_ _18655_/CLK _18622_/D vssd1 vssd1 vccd1 vccd1 _18622_/Q sky130_fd_sc_hd__dfxtp_1
X_15834_ _15834_/A vssd1 vssd1 vccd1 vccd1 _15834_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18553_ _18688_/CLK _18553_/D vssd1 vssd1 vccd1 vccd1 _18553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15765_ _15765_/A vssd1 vssd1 vccd1 vccd1 _15765_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12977_ _17004_/A vssd1 vssd1 vccd1 vccd1 _17646_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14249__C _14279_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17504_ _19658_/Q vssd1 vssd1 vccd1 vccd1 _17505_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11928_ hold2/A _12084_/S _12085_/A _11927_/X vssd1 vssd1 vccd1 vccd1 _11928_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14716_ _18809_/Q _13661_/X _14716_/S vssd1 vssd1 vccd1 vccd1 _14717_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18484_ _18544_/CLK _18484_/D vssd1 vssd1 vccd1 vccd1 _18484_/Q sky130_fd_sc_hd__dfxtp_2
X_15696_ _15696_/A vssd1 vssd1 vccd1 vccd1 _18924_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17435_ _17109_/X _19626_/Q _17437_/S vssd1 vssd1 vccd1 vccd1 _17436_/A sky130_fd_sc_hd__mux2_1
X_14647_ _14647_/A vssd1 vssd1 vccd1 vccd1 _18782_/D sky130_fd_sc_hd__clkbuf_1
X_11859_ _11731_/X _11857_/X _11858_/Y _11723_/X _19006_/Q vssd1 vssd1 vccd1 vccd1
+ _11860_/D sky130_fd_sc_hd__a32o_4
Xclkbuf_leaf_113_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19683_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14578_ _14578_/A vssd1 vssd1 vccd1 vccd1 _18762_/D sky130_fd_sc_hd__clkbuf_1
X_17366_ _17366_/A vssd1 vssd1 vccd1 vccd1 _19595_/D sky130_fd_sc_hd__clkbuf_1
X_19105_ _19986_/CLK _19105_/D vssd1 vssd1 vccd1 vccd1 _19105_/Q sky130_fd_sc_hd__dfxtp_1
X_16317_ _16400_/S vssd1 vssd1 vccd1 vccd1 _16330_/S sky130_fd_sc_hd__clkbuf_4
X_13529_ hold6/A _13529_/B vssd1 vssd1 vccd1 vccd1 _13529_/X sky130_fd_sc_hd__or2_1
XFILLER_174_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17297_ _17297_/A vssd1 vssd1 vccd1 vccd1 _19564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19036_ _19664_/CLK _19036_/D vssd1 vssd1 vccd1 vccd1 _19036_/Q sky130_fd_sc_hd__dfxtp_1
X_16248_ _16248_/A vssd1 vssd1 vccd1 vccd1 _19137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_128_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19487_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput103 _09188_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[0] sky130_fd_sc_hd__buf_2
Xoutput114 _12843_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[14] sky130_fd_sc_hd__buf_2
X_16179_ _16179_/A vssd1 vssd1 vccd1 vccd1 _19107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10367__B1 _09566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput125 _12856_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[24] sky130_fd_sc_hd__buf_2
XFILLER_154_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput136 _12829_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[5] sky130_fd_sc_hd__buf_2
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput147 _12403_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[14] sky130_fd_sc_hd__buf_2
XANTENNA__09375__A _18952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput158 _12656_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[24] sky130_fd_sc_hd__buf_2
XFILLER_115_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput169 _12140_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[5] sky130_fd_sc_hd__buf_2
XANTENNA__13609__B _13609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19938_ _20002_/CLK _19938_/D vssd1 vssd1 vccd1 vccd1 _19938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19869_ _20031_/CLK _19869_/D vssd1 vssd1 vccd1 vccd1 _19869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09622_ _10929_/A vssd1 vssd1 vccd1 vccd1 _10886_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10968__B _12835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _10502_/A vssd1 vssd1 vccd1 vccd1 _10194_/A sky130_fd_sc_hd__buf_2
XFILLER_71_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10517__S1 _10011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09484_ _09496_/A _14812_/B vssd1 vssd1 vccd1 vccd1 _12193_/A sky130_fd_sc_hd__or2_2
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11190__S1 _11108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13360__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12898__A2 _12892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 _19940_/CLK sky130_fd_sc_hd__clkbuf_16
X_10190_ _19154_/Q _19415_/Q _19314_/Q _19649_/Q _10449_/S _10185_/A vssd1 vssd1 vccd1
+ vccd1 _10191_/B sky130_fd_sc_hd__mux4_1
XFILLER_133_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10373__A3 _10372_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_160_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12900_ _12997_/A vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20009_ _20010_/CLK _20009_/D vssd1 vssd1 vccd1 vccd1 _20009_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17007__A _17007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16797__A0 _16345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13880_ _15833_/A vssd1 vssd1 vccd1 vccd1 _14447_/B sky130_fd_sc_hd__buf_4
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12831_ _12831_/A _12831_/B vssd1 vssd1 vccd1 vccd1 _12831_/Y sky130_fd_sc_hd__nor2_4
XFILLER_62_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16846__A _18937_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15550_ _18863_/Q _15547_/X _15567_/S vssd1 vssd1 vccd1 vccd1 _15551_/A sky130_fd_sc_hd__mux2_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12762_/A _15531_/B vssd1 vssd1 vccd1 vccd1 _12763_/B sky130_fd_sc_hd__and2_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_30_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _20015_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14501_/A _18734_/Q _14501_/C vssd1 vssd1 vccd1 vccd1 _14503_/B sky130_fd_sc_hd__and3_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _14398_/B _11698_/Y _11711_/X _11712_/Y vssd1 vssd1 vccd1 vccd1 _11713_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15481_ _15481_/A vssd1 vssd1 vccd1 vccd1 _18857_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16057__S _16057_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A vssd1 vssd1 vccd1 vccd1 _12693_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__14366__A _14427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17220_ _17220_/A vssd1 vssd1 vccd1 vccd1 _19530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _14452_/A _14432_/B _14432_/C vssd1 vssd1 vccd1 vccd1 _18704_/D sky130_fd_sc_hd__nor3_1
X_11644_ _11644_/A _11644_/B vssd1 vssd1 vccd1 vccd1 _11645_/C sky130_fd_sc_hd__nand2_1
XFILLER_35_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15772__A1 _09261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17151_ _17688_/A vssd1 vssd1 vccd1 vccd1 _17151_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_45_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19637_/CLK sky130_fd_sc_hd__clkbuf_16
X_14363_ _18678_/Q _14363_/B _14363_/C vssd1 vssd1 vccd1 vccd1 _14373_/D sky130_fd_sc_hd__and3_1
Xinput16 io_dbus_rdata[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_85_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11575_ _11563_/X _11574_/X _09702_/X _09843_/X _18864_/Q vssd1 vssd1 vccd1 vccd1
+ _12866_/C sky130_fd_sc_hd__a32o_4
XANTENNA__18272__S _18274_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput27 io_dbus_rdata[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_2
X_16102_ _16148_/S vssd1 vssd1 vccd1 vccd1 _16111_/S sky130_fd_sc_hd__buf_2
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput38 io_ibus_inst[13] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_4
X_13314_ _18571_/Q _13070_/A _13082_/X _18735_/Q vssd1 vssd1 vccd1 vccd1 _13314_/X
+ sky130_fd_sc_hd__a22o_1
X_10526_ _19673_/Q _19439_/Q _18504_/Q _19769_/Q _10216_/A _10218_/A vssd1 vssd1 vccd1
+ vccd1 _10527_/B sky130_fd_sc_hd__mux4_1
X_17082_ _19480_/Q _17081_/X _17088_/S vssd1 vssd1 vccd1 vccd1 _17083_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput49 io_ibus_inst[23] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14294_ _18664_/Q _18663_/Q _14297_/D vssd1 vssd1 vccd1 vccd1 _14295_/B sky130_fd_sc_hd__and3_1
X_16033_ _16044_/A vssd1 vssd1 vccd1 vccd1 _16042_/S sky130_fd_sc_hd__buf_6
XFILLER_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13245_ _13245_/A _13245_/B _11745_/Y vssd1 vssd1 vccd1 vccd1 _13245_/X sky130_fd_sc_hd__or3b_2
X_10457_ _19932_/Q _19546_/Q _19996_/Q _19115_/Q _10180_/S _09610_/A vssd1 vssd1 vccd1
+ vccd1 _10458_/B sky130_fd_sc_hd__mux4_1
XFILLER_124_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10349__B1 _09884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ _13268_/A _13172_/X _13175_/X vssd1 vssd1 vccd1 vccd1 _13176_/X sky130_fd_sc_hd__a21bo_1
X_10388_ _19373_/Q _19708_/Q _10388_/S vssd1 vssd1 vccd1 vccd1 _10388_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12127_ _18522_/Q _12128_/C _18523_/Q vssd1 vssd1 vccd1 vccd1 _12129_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__15925__A _15940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17984_ _17984_/A vssd1 vssd1 vccd1 vccd1 _19859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19723_ _20013_/CLK _19723_/D vssd1 vssd1 vccd1 vccd1 _19723_/Q sky130_fd_sc_hd__dfxtp_1
X_12058_ _18457_/Q _12472_/A vssd1 vssd1 vccd1 vccd1 _12058_/X sky130_fd_sc_hd__or2_1
X_16935_ _16935_/A vssd1 vssd1 vccd1 vccd1 _19426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12510__A1 _12501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10747__S1 _10626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ _19526_/Q vssd1 vssd1 vccd1 vccd1 _11133_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19654_ _19856_/CLK _19654_/D vssd1 vssd1 vccd1 vccd1 _19654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_6_0_clock_A clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16866_ _16323_/X _19396_/Q _16870_/S vssd1 vssd1 vccd1 vccd1 _16867_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18605_ _19941_/CLK _18605_/D vssd1 vssd1 vccd1 vccd1 _18605_/Q sky130_fd_sc_hd__dfxtp_1
X_15817_ _12003_/A _15816_/X _15798_/X input63/X vssd1 vssd1 vccd1 vccd1 _15818_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13164__B _13164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19585_ _19942_/CLK _19585_/D vssd1 vssd1 vccd1 vccd1 _19585_/Q sky130_fd_sc_hd__dfxtp_1
X_16797_ _16345_/X _19366_/Q _16797_/S vssd1 vssd1 vccd1 vccd1 _16798_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18536_ _18911_/CLK _18536_/D vssd1 vssd1 vccd1 vccd1 _18536_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _18945_/Q _15760_/B vssd1 vssd1 vccd1 vccd1 _15748_/X sky130_fd_sc_hd__or2_1
XFILLER_33_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ _18526_/CLK _18467_/D vssd1 vssd1 vccd1 vccd1 _18467_/Q sky130_fd_sc_hd__dfxtp_1
X_15679_ _15690_/A vssd1 vssd1 vccd1 vccd1 _15688_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17418_ _19619_/Q _17084_/X _17420_/S vssd1 vssd1 vccd1 vccd1 _17419_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18398_ _18409_/A vssd1 vssd1 vccd1 vccd1 _18407_/S sky130_fd_sc_hd__buf_4
XFILLER_119_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17349_ _17349_/A vssd1 vssd1 vccd1 vccd1 _19588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10683__S0 _10521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15515__A1 _18860_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19019_ _19023_/CLK _19019_/D vssd1 vssd1 vccd1 vccd1 _19019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10435__S0 _10469_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09833__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09605_ _10048_/A vssd1 vssd1 vccd1 vccd1 _09606_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18357__S _18363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17261__S _17265_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09536_ _09536_/A vssd1 vssd1 vccd1 vccd1 _09537_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11163__S1 _11015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10815__A1 _09882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09467_ _18981_/Q vssd1 vssd1 vccd1 vccd1 _09467_/X sky130_fd_sc_hd__buf_4
XFILLER_25_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_107_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15754__A1 _12032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ _11705_/A _11785_/A vssd1 vssd1 vccd1 vccd1 _09402_/C sky130_fd_sc_hd__nor2_1
XFILLER_40_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16605__S _16613_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11360_ _11309_/A _11354_/X _11359_/X _09789_/A vssd1 vssd1 vccd1 vccd1 _11360_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10311_ _19677_/Q _19443_/Q _18508_/Q _19773_/Q _09655_/A _10260_/A vssd1 vssd1 vccd1
+ vccd1 _10312_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11291_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11291_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12434__A _14966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13030_ _18460_/Q _12943_/A _12944_/A _18684_/Q _13029_/X vssd1 vssd1 vccd1 vccd1
+ _13030_/X sky130_fd_sc_hd__a221o_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10242_ _15972_/C _12858_/B vssd1 vssd1 vccd1 vccd1 _10242_/X sky130_fd_sc_hd__or2_1
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09694__A1_N _18863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15809__A2 _11860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10173_ _10335_/A _10170_/X _10172_/X _10159_/X vssd1 vssd1 vccd1 vccd1 _10173_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16340__S _16346_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09743__A _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input38_A io_ibus_inst[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14981_ _15016_/A vssd1 vssd1 vccd1 vccd1 _15132_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_59_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_5_0_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_16720_ _16720_/A vssd1 vssd1 vccd1 vccd1 _19331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13932_ _18551_/Q _13925_/C _13931_/Y vssd1 vssd1 vccd1 vccd1 _18551_/D sky130_fd_sc_hd__o21a_1
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16651_ _16651_/A vssd1 vssd1 vccd1 vccd1 _19301_/D sky130_fd_sc_hd__clkbuf_1
X_13863_ _13910_/A vssd1 vssd1 vccd1 vccd1 _14577_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15442__A0 _18854_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17171__S _17177_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ _12812_/Y _12813_/Y _12814_/S vssd1 vssd1 vccd1 vccd1 _12814_/X sky130_fd_sc_hd__mux2_1
X_15602_ _15602_/A vssd1 vssd1 vccd1 vccd1 _15611_/S sky130_fd_sc_hd__buf_2
X_19370_ _19995_/CLK _19370_/D vssd1 vssd1 vccd1 vccd1 _19370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13794_ _17030_/A vssd1 vssd1 vccd1 vccd1 _13794_/X sky130_fd_sc_hd__clkbuf_2
X_16582_ _16604_/A vssd1 vssd1 vccd1 vccd1 _16591_/S sky130_fd_sc_hd__buf_4
XFILLER_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18321_ _18321_/A vssd1 vssd1 vccd1 vccd1 _19994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15533_ _15236_/A _15530_/X _15532_/Y _15400_/A vssd1 vssd1 vccd1 vccd1 _15533_/X
+ sky130_fd_sc_hd__a31o_1
X_12745_ _12745_/A _12768_/C vssd1 vssd1 vccd1 vccd1 _12745_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11513__A _15947_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18252_ _19964_/Q _17697_/A _18252_/S vssd1 vssd1 vccd1 vccd1 _18253_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ _15384_/X _15459_/Y _15463_/Y vssd1 vssd1 vccd1 vccd1 _15465_/C sky130_fd_sc_hd__a21oi_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _18479_/Q _12556_/X _12557_/X vssd1 vssd1 vccd1 vccd1 _12676_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12559__A1 _12338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17203_ _17203_/A _17203_/B vssd1 vssd1 vccd1 vccd1 _19523_/D sky130_fd_sc_hd__nor2_1
X_14415_ _18700_/Q vssd1 vssd1 vccd1 vccd1 _14422_/C sky130_fd_sc_hd__clkbuf_1
X_11627_ _11626_/Y _11517_/X _10540_/A _11594_/A vssd1 vssd1 vccd1 vccd1 _11628_/D
+ sky130_fd_sc_hd__o22a_1
X_18183_ _17700_/X _19933_/Q _18191_/S vssd1 vssd1 vccd1 vccd1 _18184_/A sky130_fd_sc_hd__mux2_1
X_15395_ _15368_/X _15397_/B _15369_/X _15394_/X vssd1 vssd1 vccd1 vccd1 _15395_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16515__S _16519_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17134_ _17134_/A vssd1 vssd1 vccd1 vccd1 _19500_/D sky130_fd_sc_hd__clkbuf_1
X_14346_ _14356_/A _14346_/B _14350_/C vssd1 vssd1 vccd1 vccd1 _18679_/D sky130_fd_sc_hd__nor3_1
XANTENNA__10665__S0 _10724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11558_ _11558_/A _11558_/B vssd1 vssd1 vccd1 vccd1 _11558_/X sky130_fd_sc_hd__or2_1
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17065_ _17065_/A vssd1 vssd1 vccd1 vccd1 _17065_/X sky130_fd_sc_hd__clkbuf_2
X_10509_ _19210_/Q _19801_/Q _19963_/Q _19178_/Q _10319_/A _10542_/A vssd1 vssd1 vccd1
+ vccd1 _10509_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14277_ _18659_/Q _14273_/B _14276_/Y vssd1 vssd1 vccd1 vccd1 _18659_/D sky130_fd_sc_hd__o21a_1
XFILLER_155_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11489_ _09830_/A _11488_/X _11502_/A vssd1 vssd1 vccd1 vccd1 _11489_/X sky130_fd_sc_hd__a21o_1
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16016_ _13161_/X _19038_/Q _16020_/S vssd1 vssd1 vccd1 vccd1 _16017_/A sky130_fd_sc_hd__mux2_1
X_13228_ _13360_/A _18849_/Q vssd1 vssd1 vccd1 vccd1 _13228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17346__S _17348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16250__S _16258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13159_ _09532_/X _13157_/X _13158_/X vssd1 vssd1 vccd1 vccd1 _17033_/A sky130_fd_sc_hd__o21a_4
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09653__A _09653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _18024_/S vssd1 vssd1 vccd1 vccd1 _17976_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19706_ _19706_/CLK _19706_/D vssd1 vssd1 vccd1 vccd1 _19706_/Q sky130_fd_sc_hd__dfxtp_1
X_16918_ _16399_/X _19420_/Q _16918_/S vssd1 vssd1 vccd1 vccd1 _16919_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09372__B _18951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17898_ _19821_/Q _17014_/X _17904_/S vssd1 vssd1 vccd1 vccd1 _17899_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11393__S1 _11107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19637_ _19637_/CLK _19637_/D vssd1 vssd1 vccd1 vccd1 _19637_/Q sky130_fd_sc_hd__dfxtp_1
X_16849_ _16905_/A vssd1 vssd1 vccd1 vccd1 _16918_/S sky130_fd_sc_hd__buf_6
XFILLER_66_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19568_ _19824_/CLK _19568_/D vssd1 vssd1 vccd1 vccd1 _19568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09321_ _18982_/Q vssd1 vssd1 vccd1 vccd1 _09468_/A sky130_fd_sc_hd__clkbuf_4
X_18519_ _19880_/CLK _18519_/D vssd1 vssd1 vccd1 vccd1 _18519_/Q sky130_fd_sc_hd__dfxtp_1
X_19499_ _19569_/CLK _19499_/D vssd1 vssd1 vccd1 vccd1 _19499_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11470__A1 _09607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ _09283_/B _18966_/Q _09283_/D vssd1 vssd1 vccd1 vccd1 _11951_/B sky130_fd_sc_hd__or3b_2
XFILLER_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ _18973_/Q vssd1 vssd1 vccd1 vccd1 _11919_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16160__S _16162_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09563__A _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_33_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11289__A1 _11278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__A _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13813__A _17049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10860_ _19235_/Q _19730_/Q _11488_/S vssd1 vssd1 vccd1 vccd1 _10860_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11136__S1 _11050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09519_ _14811_/B vssd1 vssd1 vccd1 vccd1 _09525_/A sky130_fd_sc_hd__inv_2
XFILLER_13_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10791_ _10952_/A vssd1 vssd1 vccd1 vccd1 _10905_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12530_/A vssd1 vssd1 vccd1 vccd1 _12530_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_158_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15727__A1 hold2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12461_ _15385_/A _12461_/B vssd1 vssd1 vccd1 vccd1 _12464_/A sky130_fd_sc_hd__xnor2_1
XFILLER_32_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14200_ _18639_/Q _14200_/B vssd1 vssd1 vccd1 vccd1 _14207_/C sky130_fd_sc_hd__and2_1
XFILLER_32_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11412_ _11199_/A _11409_/X _11411_/X vssd1 vssd1 vccd1 vccd1 _11412_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12410__A0 _15947_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17020__A _17020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09738__A _11157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15180_ _14991_/X _15181_/B _15179_/X _15105_/X vssd1 vssd1 vccd1 vccd1 _15180_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12392_ _12416_/B _12392_/B vssd1 vssd1 vccd1 vccd1 _12393_/D sky130_fd_sc_hd__xor2_1
XFILLER_126_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14131_ _14133_/B _14133_/C _14130_/Y vssd1 vssd1 vccd1 vccd1 _18616_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17955__A _18011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ _19915_/Q _19529_/Q _19979_/Q _19098_/Q _10618_/A _11086_/A vssd1 vssd1 vccd1
+ vccd1 _11344_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12961__B2 _12906_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14062_ _14062_/A _18596_/Q _14062_/C vssd1 vssd1 vccd1 vccd1 _14064_/B sky130_fd_sc_hd__and3_1
X_11274_ _11258_/S _11272_/Y _11273_/Y _11073_/X vssd1 vssd1 vccd1 vccd1 _11274_/X
+ sky130_fd_sc_hd__a211o_1
X_13013_ _13945_/B _13189_/A _13009_/X _13011_/X _13012_/X vssd1 vssd1 vccd1 vccd1
+ _13542_/B sky130_fd_sc_hd__a2111o_4
X_10225_ _10344_/A _10225_/B vssd1 vssd1 vccd1 vccd1 _10225_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18870_ _19001_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 _18870_/Q sky130_fd_sc_hd__dfxtp_1
X_17821_ _19787_/Q _17007_/X _17821_/S vssd1 vssd1 vccd1 vccd1 _17822_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10156_ _20036_/Q _19874_/Q _19283_/Q _19053_/Q _10141_/X _10283_/A vssd1 vssd1 vccd1
+ vccd1 _10157_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11508__A _15940_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17752_ _17652_/X _19756_/Q _17760_/S vssd1 vssd1 vccd1 vccd1 _17753_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10087_ _20033_/Q _19871_/Q _19280_/Q _19050_/Q _09939_/A _10278_/A vssd1 vssd1 vccd1
+ vccd1 _10088_/B sky130_fd_sc_hd__mux4_1
X_14964_ _15546_/A vssd1 vssd1 vccd1 vccd1 _15243_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16703_ _19324_/Q _13771_/X _16703_/S vssd1 vssd1 vccd1 vccd1 _16704_/A sky130_fd_sc_hd__mux2_1
X_13915_ _18593_/Q _18592_/Q _18594_/Q _14045_/A vssd1 vssd1 vccd1 vccd1 _14056_/A
+ sky130_fd_sc_hd__and4_1
X_17683_ _17683_/A vssd1 vssd1 vccd1 vccd1 _19733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14895_ _14895_/A vssd1 vssd1 vccd1 vccd1 _15100_/B sky130_fd_sc_hd__buf_2
XFILLER_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19422_ _19720_/CLK _19422_/D vssd1 vssd1 vccd1 vccd1 _19422_/Q sky130_fd_sc_hd__dfxtp_1
X_16634_ _16634_/A vssd1 vssd1 vccd1 vccd1 _19293_/D sky130_fd_sc_hd__clkbuf_1
X_13846_ _18513_/Q _13845_/X _13852_/S vssd1 vssd1 vccd1 vccd1 _13847_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11127__S1 _10983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19353_ _19979_/CLK _19353_/D vssd1 vssd1 vccd1 vccd1 _19353_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09645__A1 _09568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13777_ _13777_/A vssd1 vssd1 vccd1 vccd1 _18491_/D sky130_fd_sc_hd__clkbuf_1
X_16565_ _19263_/Q _13781_/X _16569_/S vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10989_ _11252_/A _10978_/Y _10984_/X _10988_/Y vssd1 vssd1 vccd1 vccd1 _10989_/X
+ sky130_fd_sc_hd__a31o_1
X_18304_ _18350_/S vssd1 vssd1 vccd1 vccd1 _18313_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__14257__C _14264_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15516_ _15520_/A _15520_/B vssd1 vssd1 vccd1 vccd1 _15516_/Y sky130_fd_sc_hd__nand2_1
X_19284_ _20037_/CLK _19284_/D vssd1 vssd1 vccd1 vccd1 _19284_/Q sky130_fd_sc_hd__dfxtp_1
X_12728_ _18545_/Q _12673_/X _12723_/X _12727_/X vssd1 vssd1 vccd1 vccd1 _12728_/X
+ sky130_fd_sc_hd__o22a_4
X_16496_ _16496_/A vssd1 vssd1 vccd1 vccd1 _19232_/D sky130_fd_sc_hd__clkbuf_1
X_18235_ _19956_/Q _17672_/A _18241_/S vssd1 vssd1 vccd1 vccd1 _18236_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10660__C1 _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12659_ _12753_/A _12857_/B vssd1 vssd1 vccd1 vccd1 _12659_/Y sky130_fd_sc_hd__nor2_1
X_15447_ _15368_/X _15449_/B _15369_/X _15446_/X vssd1 vssd1 vccd1 vccd1 _15447_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16245__S _16247_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09648__A _10921_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18166_ _18166_/A vssd1 vssd1 vccd1 vccd1 _19925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15378_ _12443_/Y _15364_/X _15377_/X _15360_/X vssd1 vssd1 vccd1 vccd1 _15378_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_117_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17117_ _17115_/X _19495_/Q _17129_/S vssd1 vssd1 vccd1 vccd1 _17118_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17340__A0 _17179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14329_ _18674_/Q _18673_/Q _18672_/Q _14329_/D vssd1 vssd1 vccd1 vccd1 _14338_/D
+ sky130_fd_sc_hd__and4_1
X_18097_ _18853_/Q _13667_/X _18101_/S vssd1 vssd1 vccd1 vccd1 _18097_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17048_ _17048_/A vssd1 vssd1 vccd1 vccd1 _19469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12704__A1 _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17076__S _17088_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12704__B2 _11945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09870_ _11538_/A _09869_/X _09690_/X vssd1 vssd1 vccd1 vccd1 _09870_/X sky130_fd_sc_hd__o21a_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09383__A _18952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__S0 _11486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ _19488_/CLK _18999_/D vssd1 vssd1 vccd1 vccd1 _18999_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_85_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17804__S _17804_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15957__B2 _15956_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16944__A _16990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13432__A2 _12943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ _09542_/B _09542_/C _09303_/X vssd1 vssd1 vccd1 vccd1 _09535_/B sky130_fd_sc_hd__nor3b_2
XFILLER_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11153__A _11153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10877__S0 _10703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09235_ _09273_/A vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13779__S _13788_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10629__S0 _10691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ _09247_/B vssd1 vssd1 vccd1 vccd1 _09282_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__09558__A _11003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15994__S _15998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18370__S _18374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10010_ _10010_/A vssd1 vssd1 vccd1 vccd1 _10011_/A sky130_fd_sc_hd__buf_2
XANTENNA__09293__A _18937_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09999_ _09567_/A _09984_/X _09992_/X _09998_/X _09555_/A vssd1 vssd1 vccd1 vccd1
+ _09999_/X sky130_fd_sc_hd__a311o_1
XFILLER_77_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17714__S _17714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11961_ _11961_/A _11961_/B _11961_/C vssd1 vssd1 vccd1 vccd1 _11962_/B sky130_fd_sc_hd__or3_1
XFILLER_151_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10912_ _10952_/A _10912_/B vssd1 vssd1 vccd1 vccd1 _10912_/X sky130_fd_sc_hd__or2_1
X_13700_ _13700_/A vssd1 vssd1 vccd1 vccd1 _13700_/X sky130_fd_sc_hd__buf_4
XFILLER_151_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14680_ _14680_/A vssd1 vssd1 vccd1 vccd1 _18792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09970__S1 _09637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ _18814_/Q _11841_/X _11843_/X _18781_/Q _11891_/X vssd1 vssd1 vccd1 vccd1
+ _11892_/X sky130_fd_sc_hd__a221o_1
XANTENNA__15948__A1 _19009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13631_ _13630_/A _13630_/C _13207_/A vssd1 vssd1 vccd1 vccd1 _13632_/B sky130_fd_sc_hd__o21ai_1
X_10843_ _10843_/A _10843_/B vssd1 vssd1 vccd1 vccd1 _10843_/X sky130_fd_sc_hd__or2_1
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16350_ _16348_/X _19175_/Q _16362_/S vssd1 vssd1 vccd1 vccd1 _16351_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13562_ _11717_/X _13560_/X _13561_/Y _13660_/A _19001_/Q vssd1 vssd1 vccd1 vccd1
+ _13563_/A sky130_fd_sc_hd__a32o_2
X_10774_ _10824_/A _10774_/B vssd1 vssd1 vccd1 vccd1 _10774_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13689__S _13689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15301_ _15306_/A _15306_/B vssd1 vssd1 vccd1 vccd1 _15301_/Y sky130_fd_sc_hd__nand2_1
X_12513_ _12513_/A vssd1 vssd1 vccd1 vccd1 _15410_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_158_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16281_ _16281_/A vssd1 vssd1 vccd1 vccd1 _19152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13493_ _18745_/Q vssd1 vssd1 vccd1 vccd1 _14124_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18020_ _19876_/Q _17087_/X _18020_/S vssd1 vssd1 vccd1 vccd1 _18021_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09468__A _09468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12444_ _18534_/Q vssd1 vssd1 vccd1 vccd1 _12446_/A sky130_fd_sc_hd__buf_2
X_15232_ _15139_/A _15234_/A _15212_/X _15231_/X vssd1 vssd1 vccd1 vccd1 _15232_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_166_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11737__A2 _11732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17685__A _17717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15163_ _15151_/X _15153_/X _15162_/X _15005_/X vssd1 vssd1 vccd1 vccd1 _15163_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12375_ _12344_/A _12373_/Y _12424_/C _12285_/A vssd1 vssd1 vccd1 vccd1 _12375_/Y
+ sky130_fd_sc_hd__o31ai_1
XANTENNA__10407__A _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10945__B1 _09774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14114_ _18721_/Q _18723_/Q _18722_/Q _14462_/A vssd1 vssd1 vccd1 vccd1 _14471_/A
+ sky130_fd_sc_hd__and4_1
X_11326_ _11332_/A _11323_/X _11325_/X _11058_/A vssd1 vssd1 vccd1 vccd1 _11326_/X
+ sky130_fd_sc_hd__o211a_1
X_19971_ _19971_/CLK _19971_/D vssd1 vssd1 vccd1 vccd1 _19971_/Q sky130_fd_sc_hd__dfxtp_1
X_15094_ _15094_/A vssd1 vssd1 vccd1 vccd1 _15189_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14045_ _14045_/A vssd1 vssd1 vccd1 vccd1 _14051_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18922_ _18923_/CLK _18922_/D vssd1 vssd1 vccd1 vccd1 _18922_/Q sky130_fd_sc_hd__dfxtp_1
X_11257_ _11257_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11257_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10208_ _10208_/A vssd1 vssd1 vccd1 vccd1 _10209_/S sky130_fd_sc_hd__buf_4
XFILLER_122_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18853_ _19350_/CLK _18853_/D vssd1 vssd1 vccd1 vccd1 _18853_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__10173__A1 _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ _11237_/A _11187_/X _11311_/A vssd1 vssd1 vccd1 vccd1 _11188_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17624__S _17628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17804_ _17729_/X _19780_/Q _17804_/S vssd1 vssd1 vccd1 vccd1 _17805_/A sky130_fd_sc_hd__mux2_1
X_10139_ _18860_/Q _09539_/A _09547_/X _10138_/X vssd1 vssd1 vccd1 vccd1 _15974_/B
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__10142__A _10473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18784_ _19910_/CLK _18784_/D vssd1 vssd1 vccd1 vccd1 _18784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15996_ _12978_/X _19029_/Q _15998_/S vssd1 vssd1 vccd1 vccd1 _15997_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17735_ _17735_/A vssd1 vssd1 vccd1 vccd1 _17735_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14947_ _12664_/A _15177_/B _14956_/S vssd1 vssd1 vccd1 vccd1 _14947_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13662__A2 _13661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18050__A1 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17666_ _17665_/X _19728_/Q _17666_/S vssd1 vssd1 vccd1 vccd1 _17667_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15939__A1 _19006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14878_ _15355_/B _15373_/B _14948_/S vssd1 vssd1 vccd1 vccd1 _14878_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19405_ _19828_/CLK _19405_/D vssd1 vssd1 vccd1 vccd1 _19405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16617_ _19287_/Q _13857_/X _16617_/S vssd1 vssd1 vccd1 vccd1 _16618_/A sky130_fd_sc_hd__mux2_1
X_13829_ _17065_/A vssd1 vssd1 vccd1 vccd1 _13829_/X sky130_fd_sc_hd__clkbuf_2
X_17597_ _17619_/A vssd1 vssd1 vccd1 vccd1 _17606_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__14611__A1 _13629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13414__A2 _12943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19336_ _19828_/CLK _19336_/D vssd1 vssd1 vccd1 vccd1 _19336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16548_ _16604_/A vssd1 vssd1 vccd1 vccd1 _16617_/S sky130_fd_sc_hd__buf_6
XFILLER_149_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19267_ _19990_/CLK _19267_/D vssd1 vssd1 vccd1 vccd1 _19267_/Q sky130_fd_sc_hd__dfxtp_1
X_16479_ _16479_/A vssd1 vssd1 vccd1 vccd1 _19224_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13178__A1 _12967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18218_ _18218_/A vssd1 vssd1 vccd1 vccd1 _19948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19198_ _19853_/CLK _19198_/D vssd1 vssd1 vccd1 vccd1 _19198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17313__A0 _17141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__S0 _11121_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18149_ _18206_/S vssd1 vssd1 vccd1 vccd1 _18158_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__16703__S _16703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09922_ _10069_/A _09917_/X _09919_/X _09921_/X vssd1 vssd1 vccd1 vccd1 _09922_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13886__C1 _13885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09853_ _19253_/Q _19748_/Q _11534_/S vssd1 vssd1 vccd1 vccd1 _09853_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15843__A _15879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09784_ _10094_/S vssd1 vssd1 vccd1 vccd1 _09903_/A sky130_fd_sc_hd__buf_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14602__A1 _11860_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09218_ _09283_/D vssd1 vssd1 vccd1 vccd1 _09435_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _15958_/C _12850_/B vssd1 vssd1 vccd1 vccd1 _11626_/A sky130_fd_sc_hd__or2_2
XFILLER_154_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11275__S0 _11049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16613__S _16613_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12160_ _18763_/Q _12161_/B vssd1 vssd1 vccd1 vccd1 _12162_/A sky130_fd_sc_hd__and2_1
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _11111_/A vssd1 vssd1 vccd1 vccd1 _11227_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_2_2_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ _12091_/A _14914_/A vssd1 vssd1 vccd1 vccd1 _12092_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13877__C1 _13946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13341__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11042_ _11325_/A vssd1 vssd1 vccd1 vccd1 _11257_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10155__A1 _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09640__S0 _09635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15850_ _11982_/X _15842_/X _15843_/X input42/X vssd1 vssd1 vccd1 vccd1 _17204_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input20_A io_dbus_rdata[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ _14801_/A vssd1 vssd1 vccd1 vccd1 _18832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15781_ _18959_/Q _15783_/B vssd1 vssd1 vccd1 vccd1 _15781_/X sky130_fd_sc_hd__or2_1
XFILLER_29_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12993_ _14355_/B _11847_/X _12983_/X _12986_/X _12992_/X vssd1 vssd1 vccd1 vccd1
+ _13529_/B sky130_fd_sc_hd__a2111o_2
X_17520_ _19666_/Q vssd1 vssd1 vccd1 vccd1 _17521_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14732_ _18816_/Q _13710_/X _14738_/S vssd1 vssd1 vccd1 vccd1 _14733_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09943__S1 _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ _09702_/A _11438_/X _11449_/X _09842_/A _09347_/X vssd1 vssd1 vccd1 vccd1
+ _12822_/B sky130_fd_sc_hd__a32oi_4
XFILLER_45_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _17131_/X _19633_/Q _17459_/S vssd1 vssd1 vccd1 vccd1 _17452_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14663_ _14663_/A _14663_/B vssd1 vssd1 vccd1 vccd1 _14664_/A sky130_fd_sc_hd__and2_1
XFILLER_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11875_ _18737_/Q _12890_/A _09402_/D _18605_/Q _11874_/X vssd1 vssd1 vccd1 vccd1
+ _11875_/X sky130_fd_sc_hd__a221o_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output107_A _12866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _16692_/A _18208_/B vssd1 vssd1 vccd1 vccd1 _16459_/A sky130_fd_sc_hd__nor2_2
XFILLER_32_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10826_ _19139_/Q _19400_/Q _19299_/Q _19634_/Q _11467_/S _10820_/A vssd1 vssd1 vccd1
+ vccd1 _10827_/B sky130_fd_sc_hd__mux4_1
X_13614_ _18878_/Q _13614_/B vssd1 vssd1 vccd1 vccd1 _13615_/B sky130_fd_sc_hd__nand2_1
X_17382_ _17382_/A vssd1 vssd1 vccd1 vccd1 _19602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14594_ _12283_/A _13591_/X _14598_/S vssd1 vssd1 vccd1 vccd1 _14595_/B sky130_fd_sc_hd__mux2_1
XFILLER_13_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19121_ _20002_/CLK _19121_/D vssd1 vssd1 vccd1 vccd1 _19121_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_2_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16333_ _16400_/S vssd1 vssd1 vccd1 vccd1 _16346_/S sky130_fd_sc_hd__buf_4
X_10757_ _10579_/A _10748_/Y _10752_/Y _10756_/Y _09805_/A vssd1 vssd1 vccd1 vccd1
+ _10757_/X sky130_fd_sc_hd__o311a_2
X_13545_ _13589_/A _18999_/Q vssd1 vssd1 vccd1 vccd1 _13545_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_155_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11521__A _15966_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19052_ _19971_/CLK _19052_/D vssd1 vssd1 vccd1 vccd1 _19052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16264_ _16264_/A vssd1 vssd1 vccd1 vccd1 _19144_/D sky130_fd_sc_hd__clkbuf_1
X_13476_ _18895_/Q _13476_/B vssd1 vssd1 vccd1 vccd1 _13476_/X sky130_fd_sc_hd__or2_1
X_10688_ _19670_/Q _19436_/Q _18501_/Q _19766_/Q _10691_/S _10638_/A vssd1 vssd1 vccd1
+ vccd1 _10688_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18003_ _19868_/Q _17062_/X _18009_/S vssd1 vssd1 vccd1 vccd1 _18004_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12907__A1 _12874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12907__B2 _12906_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12427_ _12416_/C _12415_/X _12421_/Y _12426_/Y vssd1 vssd1 vccd1 vccd1 _12427_/X
+ sky130_fd_sc_hd__o22a_2
X_15215_ _15211_/X _15219_/B _15212_/X _15214_/X vssd1 vssd1 vccd1 vccd1 _15215_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15928__A _15928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16195_ _13283_/X _19115_/Q _16195_/S vssd1 vssd1 vccd1 vccd1 _16196_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10137__A _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18304__A _18350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15146_ _15458_/A vssd1 vssd1 vccd1 vccd1 _15146_/X sky130_fd_sc_hd__clkbuf_2
X_12358_ _15940_/C _18910_/Q _12358_/S vssd1 vssd1 vccd1 vccd1 _14883_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10394__A1 _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11309_ _11309_/A _11309_/B vssd1 vssd1 vccd1 vccd1 _11309_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19954_ _20017_/CLK _19954_/D vssd1 vssd1 vccd1 vccd1 _19954_/Q sky130_fd_sc_hd__dfxtp_1
X_15077_ _15366_/A vssd1 vssd1 vccd1 vccd1 _15077_/X sky130_fd_sc_hd__clkbuf_2
X_12289_ _12323_/A _15270_/A _12323_/C _12322_/A vssd1 vssd1 vccd1 vccd1 _12294_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13868__C1 _17203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13332__A1 _18476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ _14044_/A _14028_/B _14028_/C vssd1 vssd1 vccd1 vccd1 _18584_/D sky130_fd_sc_hd__nor3_1
X_18905_ _19001_/CLK _18905_/D vssd1 vssd1 vccd1 vccd1 _18905_/Q sky130_fd_sc_hd__dfxtp_1
X_19885_ _19885_/CLK _19885_/D vssd1 vssd1 vccd1 vccd1 _19885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18836_ _19324_/CLK _18836_/D vssd1 vssd1 vccd1 vccd1 _18836_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09661__A _10972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18767_ _19899_/CLK _18767_/D vssd1 vssd1 vccd1 vccd1 _18767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15979_ _19023_/Q _14803_/X _15978_/X vssd1 vssd1 vccd1 vccd1 _19023_/D sky130_fd_sc_hd__a21o_1
XFILLER_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17718_ _17716_/X _19744_/Q _17730_/S vssd1 vssd1 vccd1 vccd1 _17719_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09934__S1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18698_ _18744_/CLK _18698_/D vssd1 vssd1 vccd1 vccd1 _18698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17649_ _17649_/A vssd1 vssd1 vccd1 vccd1 _17649_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18185__S _18191_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16585__A1 _13810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19319_ _19846_/CLK _19319_/D vssd1 vssd1 vccd1 vccd1 _19319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12527__A _18473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14899__A1 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16433__S _16435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10047__A _15970_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17837__A1 _17030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15848__B1 _15789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09905_ _19157_/Q _19418_/Q _19317_/Q _19652_/Q _09903_/A _09824_/A vssd1 vssd1 vccd1
+ vccd1 _09906_/B sky130_fd_sc_hd__mux4_1
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13792__S _13804_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20025_ _20025_/CLK _20025_/D vssd1 vssd1 vccd1 vccd1 _20025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10232__S1 _10013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09836_ _19685_/Q _19451_/Q _18516_/Q _19781_/Q _09733_/X _09768_/X vssd1 vssd1 vccd1
+ vccd1 _09836_/X sky130_fd_sc_hd__mux4_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09571__A _11278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _09940_/A vssd1 vssd1 vccd1 vccd1 _09824_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14189__A _14189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16025__A0 _13238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__S1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _09698_/A _09698_/B _09698_/C vssd1 vssd1 vccd1 vccd1 _09698_/X sky130_fd_sc_hd__and3_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11660_ _11660_/A _14812_/A vssd1 vssd1 vccd1 vccd1 _11660_/Y sky130_fd_sc_hd__nand2_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15784__C1 _13885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10611_ _18440_/Q _19469_/Q _19506_/Q _19080_/Q _10655_/S _09607_/A vssd1 vssd1 vccd1
+ vccd1 _10611_/X sky130_fd_sc_hd__mux4_1
X_11591_ _11591_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13330_ _18779_/Q _14555_/B vssd1 vssd1 vccd1 vccd1 _13330_/X sky130_fd_sc_hd__and2_1
X_10542_ _10542_/A _10542_/B vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__and2_1
XANTENNA__15536__C1 _15954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ _13261_/A _13261_/B vssd1 vssd1 vccd1 vccd1 _17052_/A sky130_fd_sc_hd__nor2_4
X_10473_ _10473_/A vssd1 vssd1 vccd1 vccd1 _10473_/X sky130_fd_sc_hd__buf_2
XFILLER_10_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13011__B1 _11794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16343__S _16346_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12212_ _11459_/A _18905_/Q _12358_/S vssd1 vssd1 vccd1 vccd1 _14871_/A sky130_fd_sc_hd__mux2_1
X_15000_ _15384_/A vssd1 vssd1 vccd1 vccd1 _15305_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09746__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13562__A1 _11717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13192_ _18804_/Q _11841_/X _11843_/X _12399_/A _13191_/X vssd1 vssd1 vccd1 vccd1
+ _13192_/X sky130_fd_sc_hd__a221o_2
XFILLER_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input68_A io_irq_spi_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15839__B1 _15789_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ _12143_/A _15160_/A vssd1 vssd1 vccd1 vccd1 _12209_/C sky130_fd_sc_hd__or2_1
XANTENNA__09465__B _12260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16951_ _16342_/X _19434_/Q _16953_/S vssd1 vssd1 vccd1 vccd1 _16952_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12074_ _18760_/Q _12059_/X _12072_/Y _13595_/A vssd1 vssd1 vccd1 vccd1 _12074_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17174__S _17177_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15902_ _15902_/A vssd1 vssd1 vccd1 vccd1 _18994_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15483__A _15487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ _11145_/A _11016_/X _11018_/X _11024_/Y vssd1 vssd1 vccd1 vccd1 _11025_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_19670_ _19993_/CLK _19670_/D vssd1 vssd1 vccd1 vccd1 _19670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16882_ _16882_/A vssd1 vssd1 vccd1 vccd1 _19403_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11420__S0 _09586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16298__B _16474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18621_ _18653_/CLK _18621_/D vssd1 vssd1 vccd1 vccd1 _18621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15833_ _15833_/A vssd1 vssd1 vccd1 vccd1 _15871_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14099__A _14099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17902__S _17904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18552_ _18693_/CLK _18552_/D vssd1 vssd1 vccd1 vccd1 _18552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _09454_/B _15752_/X _15763_/X _15756_/X vssd1 vssd1 vccd1 vccd1 _18951_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _12967_/X _12975_/X _12906_/A input26/X vssd1 vssd1 vccd1 vccd1 _17004_/A
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _17503_/A vssd1 vssd1 vccd1 vccd1 _19657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _14715_/A vssd1 vssd1 vccd1 vccd1 _18808_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16567__A1 _13784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11927_ _15847_/A _12033_/S _12175_/A _09468_/A _14821_/A vssd1 vssd1 vccd1 vccd1
+ _11927_/X sky130_fd_sc_hd__a221o_1
X_18483_ _18544_/CLK _18483_/D vssd1 vssd1 vccd1 vccd1 _18483_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__15930__B _15930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15695_ _18924_/Q _18545_/Q _15699_/S vssd1 vssd1 vccd1 vccd1 _15696_/A sky130_fd_sc_hd__mux2_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17203__A _17203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17434_ _17434_/A vssd1 vssd1 vccd1 vccd1 _19625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14646_ _14646_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14647_/A sky130_fd_sc_hd__and2_1
X_11858_ _13726_/A _19006_/Q vssd1 vssd1 vccd1 vccd1 _11858_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10809_ _19140_/Q _19401_/Q _19300_/Q _19635_/Q _10797_/X _10793_/X vssd1 vssd1 vccd1
+ vccd1 _10809_/X sky130_fd_sc_hd__mux4_1
X_17365_ _19595_/Q _17007_/X _17365_/S vssd1 vssd1 vccd1 vccd1 _17366_/A sky130_fd_sc_hd__mux2_1
X_11789_ _18789_/Q _11778_/Y _11782_/X _11788_/X vssd1 vssd1 vccd1 vccd1 _11796_/A
+ sky130_fd_sc_hd__a211o_2
X_14577_ _14577_/A _14577_/B vssd1 vssd1 vccd1 vccd1 _14578_/A sky130_fd_sc_hd__and2_1
XFILLER_158_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19104_ _19986_/CLK _19104_/D vssd1 vssd1 vccd1 vccd1 _19104_/Q sky130_fd_sc_hd__dfxtp_1
X_16316_ _17652_/A vssd1 vssd1 vccd1 vccd1 _16316_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11800__A1 _18997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13528_ _13656_/A vssd1 vssd1 vccd1 vccd1 _13528_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11800__B2 _11831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17296_ _17115_/X _19564_/Q _17304_/S vssd1 vssd1 vccd1 vccd1 _17297_/A sky130_fd_sc_hd__mux2_1
X_19035_ _19824_/CLK _19035_/D vssd1 vssd1 vccd1 vccd1 _19035_/Q sky130_fd_sc_hd__dfxtp_1
X_16247_ _13115_/X _19137_/Q _16247_/S vssd1 vssd1 vccd1 vccd1 _16248_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13459_ _12956_/A _09914_/Y _13458_/Y _13145_/A vssd1 vssd1 vccd1 vccd1 _13460_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput104 _14791_/A vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[1] sky130_fd_sc_hd__buf_2
X_16178_ _13150_/X _19107_/Q _16184_/S vssd1 vssd1 vccd1 vccd1 _16179_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput115 _12844_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[15] sky130_fd_sc_hd__buf_2
XFILLER_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput126 _12857_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[25] sky130_fd_sc_hd__buf_2
XFILLER_142_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput137 _12830_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[6] sky130_fd_sc_hd__buf_2
XFILLER_126_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15129_ _14951_/X _14939_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _15129_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput148 _12427_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[15] sky130_fd_sc_hd__buf_2
Xoutput159 _12681_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[25] sky130_fd_sc_hd__buf_2
XFILLER_130_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19937_ _20032_/CLK _19937_/D vssd1 vssd1 vccd1 vccd1 _19937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15393__A _15393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19868_ _19868_/CLK _19868_/D vssd1 vssd1 vccd1 vccd1 _19868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09391__A _18950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ _11006_/A vssd1 vssd1 vccd1 vccd1 _10929_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18819_ _18819_/CLK _18819_/D vssd1 vssd1 vccd1 vccd1 _18819_/Q sky130_fd_sc_hd__dfxtp_1
X_19799_ _19976_/CLK _19799_/D vssd1 vssd1 vccd1 vccd1 _19799_/Q sky130_fd_sc_hd__dfxtp_1
X_09552_ _10668_/A vssd1 vssd1 vccd1 vccd1 _10502_/A sky130_fd_sc_hd__buf_2
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09483_ _11941_/B vssd1 vssd1 vccd1 vccd1 _14812_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12292__A1 _09467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18209__A _18265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13360__B _18857_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17259__S _17265_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16730__A1 _13810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14472__A _14472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__A _09566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10358__A1 _10200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14191__B _14197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15297__A1 _18844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_103_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13816__A _17052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11402__S0 _11356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15049__B2 _11971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20008_ _20040_/CLK _20008_/D vssd1 vssd1 vccd1 vccd1 _20008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09819_ _09819_/A vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__buf_2
XFILLER_59_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10530__A1 _10424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12830_ _12831_/A _12830_/B vssd1 vssd1 vccd1 vccd1 _12830_/Y sky130_fd_sc_hd__nor2_8
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16846__B _16846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12762_/A _15531_/B vssd1 vssd1 vccd1 vccd1 _12786_/A sky130_fd_sc_hd__nor2_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14501_/A _14501_/C _14499_/Y vssd1 vssd1 vccd1 vccd1 _18733_/D sky130_fd_sc_hd__o21a_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17023__A _17023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11712_ _11869_/A _11712_/B vssd1 vssd1 vccd1 vccd1 _11712_/Y sky130_fd_sc_hd__nor2_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11491__C1 _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _18857_/Q _15479_/X _15480_/S vssd1 vssd1 vccd1 vccd1 _15481_/A sky130_fd_sc_hd__mux2_1
X_12692_ _12729_/B _12692_/B vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__xnor2_4
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11643_ _11643_/A vssd1 vssd1 vccd1 vccd1 _11644_/B sky130_fd_sc_hd__inv_2
XANTENNA__13270__B _13290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _18704_/Q _14433_/C _14431_/C vssd1 vssd1 vccd1 vccd1 _14432_/C sky130_fd_sc_hd__and3_1
XANTENNA__10386__S _10470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13232__B1 _13093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10046__B1 _09913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17150_ _17150_/A vssd1 vssd1 vccd1 vccd1 _19505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ _11574_/A _11574_/B _11574_/C vssd1 vssd1 vccd1 vccd1 _11574_/X sky130_fd_sc_hd__or3_1
Xclkbuf_opt_1_0_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_14362_ _18685_/Q _18684_/Q _18679_/Q vssd1 vssd1 vccd1 vccd1 _14363_/C sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_28_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 io_dbus_rdata[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16101_ _16101_/A vssd1 vssd1 vccd1 vccd1 _19073_/D sky130_fd_sc_hd__clkbuf_1
Xinput28 io_dbus_rdata[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_4
Xinput39 io_ibus_inst[14] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_8
X_10525_ _10516_/Y _10518_/Y _10520_/Y _10524_/Y _09821_/A vssd1 vssd1 vccd1 vccd1
+ _10525_/X sky130_fd_sc_hd__o221a_1
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13313_ _18667_/Q _13081_/X _11687_/X _18635_/Q vssd1 vssd1 vccd1 vccd1 _13313_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17081_ _17081_/A vssd1 vssd1 vccd1 vccd1 _17081_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14293_ _14479_/A vssd1 vssd1 vccd1 vccd1 _14319_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16032_ _16032_/A vssd1 vssd1 vccd1 vccd1 _19045_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09476__A _15139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ _13642_/A _13256_/C _12897_/X vssd1 vssd1 vccd1 vccd1 _13244_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_171_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10456_ _09566_/A _10451_/X _10453_/X _10455_/X _10194_/A vssd1 vssd1 vccd1 vccd1
+ _10456_/X sky130_fd_sc_hd__a221o_1
XFILLER_143_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13175_ _13175_/A _13175_/B _13183_/B vssd1 vssd1 vccd1 vccd1 _13175_/X sky130_fd_sc_hd__or3_1
X_10387_ _10424_/A _10387_/B vssd1 vssd1 vccd1 vccd1 _10387_/X sky130_fd_sc_hd__and2_1
XFILLER_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12126_ _18523_/Q _12303_/B vssd1 vssd1 vccd1 vccd1 _12139_/A sky130_fd_sc_hd__or2_1
XFILLER_2_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17983_ _19859_/Q _17033_/X _17987_/S vssd1 vssd1 vccd1 vccd1 _17984_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15925__B _15955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19722_ _20013_/CLK _19722_/D vssd1 vssd1 vccd1 vccd1 _19722_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15417__S _15480_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _12791_/A _12046_/Y _12054_/X _12056_/X vssd1 vssd1 vccd1 vccd1 _12057_/X
+ sky130_fd_sc_hd__a211o_1
X_16934_ _16316_/X _19426_/Q _16942_/S vssd1 vssd1 vccd1 vccd1 _16935_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16102__A _16148_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11849__B2 _18690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11008_ _11001_/A _11007_/X _09683_/A vssd1 vssd1 vccd1 vccd1 _11008_/Y sky130_fd_sc_hd__o21ai_1
X_19653_ _20007_/CLK _19653_/D vssd1 vssd1 vccd1 vccd1 _19653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16865_ _16865_/A vssd1 vssd1 vccd1 vccd1 _19395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17632__S _17632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18604_ _19941_/CLK _18604_/D vssd1 vssd1 vccd1 vccd1 _18604_/Q sky130_fd_sc_hd__dfxtp_1
X_15816_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15816_/X sky130_fd_sc_hd__clkbuf_2
X_19584_ _20034_/CLK _19584_/D vssd1 vssd1 vccd1 vccd1 _19584_/Q sky130_fd_sc_hd__dfxtp_1
X_16796_ _16796_/A vssd1 vssd1 vccd1 vccd1 _19365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18535_ _19001_/CLK _18535_/D vssd1 vssd1 vccd1 vccd1 _18535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _15747_/A vssd1 vssd1 vccd1 vccd1 _15760_/B sky130_fd_sc_hd__clkbuf_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09675__C1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12959_ _18867_/Q vssd1 vssd1 vccd1 vccd1 _13504_/A sky130_fd_sc_hd__buf_2
XANTENNA__13471__B1 _11776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18466_ _18994_/CLK _18466_/D vssd1 vssd1 vccd1 vccd1 _18466_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15678_ _15678_/A vssd1 vssd1 vccd1 vccd1 _18916_/D sky130_fd_sc_hd__clkbuf_1
X_17417_ _17417_/A vssd1 vssd1 vccd1 vccd1 _19618_/D sky130_fd_sc_hd__clkbuf_1
X_14629_ _14629_/A _14629_/B vssd1 vssd1 vccd1 vccd1 _14630_/A sky130_fd_sc_hd__and2_1
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18397_ _18397_/A vssd1 vssd1 vccd1 vccd1 _20028_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12077__A _12077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17348_ _17192_/X _19588_/Q _17348_/S vssd1 vssd1 vccd1 vccd1 _17349_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17079__S _17088_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17279_ _17279_/A vssd1 vssd1 vccd1 vccd1 _19557_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16712__A1 _13784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19018_ _19973_/CLK _19018_/D vssd1 vssd1 vccd1 vccd1 _19018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12524__B _18537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10435__S1 _10163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09604_ _10709_/A vssd1 vssd1 vccd1 vccd1 _10048_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09535_ _09909_/A _09535_/B vssd1 vssd1 vccd1 vccd1 _09536_/A sky130_fd_sc_hd__and2_1
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16158__S _16162_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10995__A _11409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _09466_/A _11920_/C _09514_/C vssd1 vssd1 vccd1 vccd1 _12055_/C sky130_fd_sc_hd__or3_2
XFILLER_19_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09397_ _09403_/A vssd1 vssd1 vccd1 vccd1 _11785_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13214__B1 _13211_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_174_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18911_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12715__A _12715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _10107_/X _10303_/Y _10305_/Y _10307_/Y _10309_/Y vssd1 vssd1 vccd1 vccd1
+ _10310_/X sky130_fd_sc_hd__o32a_1
XFILLER_152_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11290_ _11283_/Y _11285_/Y _11287_/Y _11289_/Y _09549_/A vssd1 vssd1 vccd1 vccd1
+ _11291_/B sky130_fd_sc_hd__o221a_1
XFILLER_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_189_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19524_/CLK sky130_fd_sc_hd__clkbuf_16
X_10241_ _15972_/C _12858_/B vssd1 vssd1 vccd1 vccd1 _10246_/B sky130_fd_sc_hd__and2_1
XANTENNA__10235__A _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10172_ _10172_/A _10172_/B vssd1 vssd1 vccd1 vccd1 _10172_/X sky130_fd_sc_hd__or2_1
XFILLER_106_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10751__A1 _10690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_112_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _20037_/CLK sky130_fd_sc_hd__clkbuf_16
X_14980_ _14903_/X _14979_/X _15117_/S vssd1 vssd1 vccd1 vccd1 _14980_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13931_ _13967_/A _13936_/C vssd1 vssd1 vccd1 vccd1 _13931_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16650_ _16342_/X _19301_/Q _16652_/S vssd1 vssd1 vccd1 vccd1 _16651_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13862_ _13862_/A vssd1 vssd1 vccd1 vccd1 _18518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15442__A1 _15441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_127_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19010_/CLK sky130_fd_sc_hd__clkbuf_16
X_15601_ _15601_/A vssd1 vssd1 vccd1 vccd1 _18882_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12813_ _18549_/Q _12813_/B vssd1 vssd1 vccd1 vccd1 _12813_/Y sky130_fd_sc_hd__xnor2_1
X_16581_ _16581_/A vssd1 vssd1 vccd1 vccd1 _19270_/D sky130_fd_sc_hd__clkbuf_1
X_13793_ _13793_/A vssd1 vssd1 vccd1 vccd1 _18496_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13453__B1 _12984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18320_ _17691_/X _19994_/Q _18324_/S vssd1 vssd1 vccd1 vccd1 _18321_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ _15181_/A _15527_/Y _15531_/Y vssd1 vssd1 vccd1 vccd1 _15532_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _18546_/Q vssd1 vssd1 vccd1 vccd1 _12745_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18392__A0 _17691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _18251_/A vssd1 vssd1 vccd1 vccd1 _19963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11513__B _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15463_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18283__S _18291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _15482_/A _12674_/Y _12697_/S vssd1 vssd1 vccd1 vccd1 _12675_/X sky130_fd_sc_hd__mux2_1
X_17202_ _17202_/A vssd1 vssd1 vccd1 vccd1 _19522_/D sky130_fd_sc_hd__clkbuf_1
X_14414_ _18699_/Q _14410_/C _14413_/Y vssd1 vssd1 vccd1 vccd1 _18699_/D sky130_fd_sc_hd__o21a_1
XANTENNA__14953__A0 _12783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18182_ _18193_/A vssd1 vssd1 vccd1 vccd1 _18191_/S sky130_fd_sc_hd__buf_4
XFILLER_129_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11626_ _11626_/A vssd1 vssd1 vccd1 vccd1 _11626_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15394_ _15506_/A _15397_/A vssd1 vssd1 vccd1 vccd1 _15394_/X sky130_fd_sc_hd__or2_1
XFILLER_128_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17133_ _17131_/X _19500_/Q _17145_/S vssd1 vssd1 vccd1 vccd1 _17134_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14345_ _18679_/Q _14345_/B _14373_/C vssd1 vssd1 vccd1 vccd1 _14350_/C sky130_fd_sc_hd__and3_1
XFILLER_7_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10665__S1 _10820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11557_ _18455_/Q _19484_/Q _19521_/Q _19095_/Q _11553_/X _11565_/A vssd1 vssd1 vccd1
+ vccd1 _11558_/B sky130_fd_sc_hd__mux4_2
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17064_ _17064_/A vssd1 vssd1 vccd1 vccd1 _19474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ _10508_/A _10508_/B vssd1 vssd1 vccd1 vccd1 _10508_/Y sky130_fd_sc_hd__nor2_1
X_11488_ _19237_/Q _19732_/Q _11488_/S vssd1 vssd1 vccd1 vccd1 _11488_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output99_A _12150_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14276_ _14288_/A _14287_/D vssd1 vssd1 vccd1 vccd1 _14276_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16015_ _16015_/A vssd1 vssd1 vccd1 vccd1 _19037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10439_ _20029_/Q _19867_/Q _19276_/Q _19046_/Q _10141_/X _10283_/A vssd1 vssd1 vccd1
+ vccd1 _10439_/X sky130_fd_sc_hd__mux4_1
X_13227_ _13227_/A vssd1 vssd1 vccd1 vccd1 _13227_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14840__A _14966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13158_ input4/X _13091_/X _13094_/X vssd1 vssd1 vccd1 vccd1 _13158_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _12108_/A _12108_/B _12059_/X vssd1 vssd1 vccd1 vccd1 _12109_/X sky130_fd_sc_hd__o21a_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17966_ _17966_/A vssd1 vssd1 vccd1 vccd1 _19851_/D sky130_fd_sc_hd__clkbuf_1
X_13089_ _13175_/A _13089_/B _13131_/C vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__or3_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19705_ _20027_/CLK _19705_/D vssd1 vssd1 vccd1 vccd1 _19705_/Q sky130_fd_sc_hd__dfxtp_1
X_16917_ _16917_/A vssd1 vssd1 vccd1 vccd1 _19419_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09372__C _18950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17897_ _17897_/A vssd1 vssd1 vccd1 vccd1 _19820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19636_ _19636_/CLK _19636_/D vssd1 vssd1 vccd1 vccd1 _19636_/Q sky130_fd_sc_hd__dfxtp_1
X_16848_ _17426_/B _17954_/B vssd1 vssd1 vccd1 vccd1 _16905_/A sky130_fd_sc_hd__or2_2
XFILLER_66_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13444__A0 _13443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19567_ _19567_/CLK _19567_/D vssd1 vssd1 vccd1 vccd1 _19567_/Q sky130_fd_sc_hd__dfxtp_1
X_16779_ _16779_/A vssd1 vssd1 vccd1 vccd1 _19357_/D sky130_fd_sc_hd__clkbuf_1
X_09320_ _18939_/Q vssd1 vssd1 vccd1 vccd1 _12913_/A sky130_fd_sc_hd__inv_2
XFILLER_34_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18518_ _19880_/CLK _18518_/D vssd1 vssd1 vccd1 vccd1 _18518_/Q sky130_fd_sc_hd__dfxtp_1
X_19498_ _20017_/CLK _19498_/D vssd1 vssd1 vccd1 vccd1 _19498_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10353__S0 _10356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_91_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 _20031_/CLK sky130_fd_sc_hd__clkbuf_16
X_09251_ _09306_/A _11919_/C _09246_/X _09248_/X _09516_/A vssd1 vssd1 vccd1 vccd1
+ _11932_/B sky130_fd_sc_hd__o32a_1
X_18449_ _20033_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16706__S _16714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14944__A0 _12715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09182_ _09492_/A vssd1 vssd1 vccd1 vccd1 _14813_/A sky130_fd_sc_hd__inv_8
XFILLER_147_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11758__B1 _14555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12970__A2 _11776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13380__C1 _13376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19990_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18368__S _18374_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17272__S _17276_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09518_ _11941_/A vssd1 vssd1 vccd1 vccd1 _14805_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_59_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19995_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_140_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10790_ _10843_/A _10790_/B vssd1 vssd1 vccd1 vccd1 _10790_/Y sky130_fd_sc_hd__nor2_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _11950_/A _09272_/A _09279_/X _09521_/A vssd1 vssd1 vccd1 vccd1 _11983_/S
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12460_ _12514_/A _12458_/Y _12515_/A vssd1 vssd1 vccd1 vccd1 _12461_/B sky130_fd_sc_hd__o21ai_1
XFILLER_166_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11411_ _11320_/A _11410_/X _11335_/A vssd1 vssd1 vccd1 vccd1 _11411_/X sky130_fd_sc_hd__a21o_1
X_12391_ _18532_/Q vssd1 vssd1 vccd1 vccd1 _12416_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12445__A _12446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11342_ _11344_/A _11341_/X _09789_/A vssd1 vssd1 vccd1 vccd1 _11342_/Y sky130_fd_sc_hd__o21ai_1
X_14130_ _14133_/B _14133_/C _14102_/X vssd1 vssd1 vccd1 vccd1 _14130_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14061_ _14062_/A _14062_/C _14060_/Y vssd1 vssd1 vccd1 vccd1 _18595_/D sky130_fd_sc_hd__o21a_1
X_11273_ _11273_/A _19227_/Q vssd1 vssd1 vccd1 vccd1 _11273_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10224_ _19154_/Q _19415_/Q _19314_/Q _19649_/Q _10166_/S _10223_/X vssd1 vssd1 vccd1
+ vccd1 _10225_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input50_A io_ibus_inst[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13012_ _18587_/Q _11851_/A _11855_/B _18719_/Q vssd1 vssd1 vccd1 vccd1 _13012_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17820_ _17820_/A vssd1 vssd1 vccd1 vccd1 _19786_/D sky130_fd_sc_hd__clkbuf_1
X_10155_ _10335_/A _10154_/X _09779_/A vssd1 vssd1 vccd1 vccd1 _10155_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17751_ _17808_/S vssd1 vssd1 vccd1 vccd1 _17760_/S sky130_fd_sc_hd__clkbuf_4
X_10086_ _10007_/A _10085_/X _09837_/A vssd1 vssd1 vccd1 vccd1 _10086_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11508__B _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14963_ _14858_/X _14922_/X _14962_/X vssd1 vssd1 vccd1 vccd1 _14965_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__18278__S _18278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output137_A _12830_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16702_ _16702_/A vssd1 vssd1 vccd1 vccd1 _19323_/D sky130_fd_sc_hd__clkbuf_1
X_13914_ _18589_/Q _18591_/Q _18590_/Q _14037_/A vssd1 vssd1 vccd1 vccd1 _14045_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_75_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17682_ _17681_/X _19733_/Q _17682_/S vssd1 vssd1 vccd1 vccd1 _17683_/A sky130_fd_sc_hd__mux2_1
X_14894_ _14876_/X _14891_/X _15202_/S vssd1 vssd1 vccd1 vccd1 _14894_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19421_ _19720_/CLK _19421_/D vssd1 vssd1 vccd1 vccd1 _19421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16633_ _16316_/X _19293_/Q _16641_/S vssd1 vssd1 vccd1 vccd1 _16634_/A sky130_fd_sc_hd__mux2_1
X_13845_ _17081_/A vssd1 vssd1 vccd1 vccd1 _13845_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13426__B1 _13368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13215__S _13215_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19352_ _19979_/CLK _19352_/D vssd1 vssd1 vccd1 vccd1 _19352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16564_ _16564_/A vssd1 vssd1 vccd1 vccd1 _19262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13776_ _18491_/Q _13774_/X _13788_/S vssd1 vssd1 vccd1 vccd1 _13777_/A sky130_fd_sc_hd__mux2_1
X_10988_ _11278_/A _10988_/B vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__nor2_1
X_18303_ _18303_/A vssd1 vssd1 vccd1 vccd1 _19986_/D sky130_fd_sc_hd__clkbuf_1
X_15515_ _18860_/Q _15457_/X _15514_/X vssd1 vssd1 vccd1 vccd1 _18860_/D sky130_fd_sc_hd__o21a_1
X_19283_ _20036_/CLK _19283_/D vssd1 vssd1 vccd1 vccd1 _19283_/Q sky130_fd_sc_hd__dfxtp_1
X_12727_ _12170_/X _12725_/X _12726_/Y _12234_/B vssd1 vssd1 vccd1 vccd1 _12727_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__16526__S _16530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16495_ _19232_/Q _13784_/X _16497_/S vssd1 vssd1 vccd1 vccd1 _16496_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17211__A _17267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18234_ _18234_/A vssd1 vssd1 vccd1 vccd1 _19955_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09929__A _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15446_ _15506_/A _15449_/A vssd1 vssd1 vccd1 vccd1 _15446_/X sky130_fd_sc_hd__or2_1
X_12658_ _12658_/A vssd1 vssd1 vccd1 vccd1 _12753_/A sky130_fd_sc_hd__buf_2
XFILLER_157_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18165_ _17675_/X _19925_/Q _18169_/S vssd1 vssd1 vccd1 vccd1 _18166_/A sky130_fd_sc_hd__mux2_1
X_11609_ _11609_/A _11269_/X vssd1 vssd1 vccd1 vccd1 _11611_/B sky130_fd_sc_hd__or2b_1
XFILLER_117_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15377_ _15329_/X _15349_/X _15376_/X _15342_/X vssd1 vssd1 vccd1 vccd1 _15377_/X
+ sky130_fd_sc_hd__o211a_1
X_12589_ _12634_/A _12854_/B vssd1 vssd1 vccd1 vccd1 _12589_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17116_ _17199_/S vssd1 vssd1 vccd1 vccd1 _17129_/S sky130_fd_sc_hd__clkbuf_4
X_14328_ _14479_/A vssd1 vssd1 vccd1 vccd1 _14413_/A sky130_fd_sc_hd__buf_2
XFILLER_143_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18096_ _18096_/A vssd1 vssd1 vccd1 vccd1 _19900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17357__S _17365_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17047_ _19469_/Q _17046_/X _17056_/S vssd1 vssd1 vccd1 vccd1 _17048_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16261__S _16269_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14259_ _14265_/A _14259_/B vssd1 vssd1 vccd1 vccd1 _14259_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09664__A _09664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09383__B _18951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10603__A _10836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__S1 _10625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ _18998_/CLK _18998_/D vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17949_ _17949_/A vssd1 vssd1 vccd1 vccd1 _19844_/D sky130_fd_sc_hd__clkbuf_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15605__S _15611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16474__C_N _16298_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19619_ _20037_/CLK _19619_/D vssd1 vssd1 vccd1 vccd1 _19619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11428__C1 _19526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09303_ _18977_/Q _09322_/A _09301_/X _09302_/Y _18827_/Q vssd1 vssd1 vccd1 vccd1
+ _09303_/X sky130_fd_sc_hd__o221a_1
XFILLER_55_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12964__S _13003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10877__S1 _10663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14745__A _14745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09234_ _18990_/Q _18989_/Q vssd1 vssd1 vccd1 vccd1 _09273_/A sky130_fd_sc_hd__or2_1
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18108__A0 _18856_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09165_ _18964_/Q _18963_/Q _18962_/Q _18961_/Q vssd1 vssd1 vccd1 vccd1 _09247_/B
+ sky130_fd_sc_hd__or4bb_2
XFILLER_147_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10629__S1 _10626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13795__S _13804_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16171__S _16173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15893__A1 _12260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09574__A _11473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15893__B2 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09998_ _09973_/A _09993_/X _09997_/X _09980_/X vssd1 vssd1 vccd1 vccd1 _09998_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11960_ _11960_/A vssd1 vssd1 vccd1 vccd1 _11960_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10911_ _19138_/Q _19399_/Q _19298_/Q _19633_/Q _10954_/S _10893_/A vssd1 vssd1 vccd1
+ vccd1 _10912_/B sky130_fd_sc_hd__mux4_1
XFILLER_45_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11891_ _19905_/Q _11845_/X _11847_/X _18702_/Q _11890_/X vssd1 vssd1 vccd1 vccd1
+ _11891_/X sky130_fd_sc_hd__a221o_1
XANTENNA__15948__A2 _15921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17730__S _17730_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11344__A _11344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13630_ _13630_/A _18880_/Q _13630_/C vssd1 vssd1 vccd1 vccd1 _13637_/B sky130_fd_sc_hd__or3_1
X_10842_ _18435_/Q _19464_/Q _19501_/Q _19075_/Q _10797_/X _10793_/X vssd1 vssd1 vccd1
+ vccd1 _10843_/B sky130_fd_sc_hd__mux4_1
XFILLER_60_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10317__S0 _10354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ _14560_/A _19001_/Q vssd1 vssd1 vccd1 vccd1 _13561_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16346__S _16346_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ _19925_/Q _19539_/Q _19989_/Q _19108_/Q _10704_/A _10048_/A vssd1 vssd1 vccd1
+ vccd1 _10774_/B sky130_fd_sc_hd__mux4_1
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15300_ _14978_/X _15123_/X _15097_/X vssd1 vssd1 vccd1 vccd1 _15415_/B sky130_fd_sc_hd__o21a_1
XANTENNA__14908__A0 _15219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12512_ _11904_/X _12850_/B _12511_/Y vssd1 vssd1 vccd1 vccd1 _12513_/A sky130_fd_sc_hd__a21oi_1
X_16280_ _13365_/X _19152_/Q _16280_/S vssd1 vssd1 vccd1 vccd1 _16281_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13492_ _13924_/B _11683_/X _11733_/X _18645_/Q vssd1 vssd1 vccd1 vccd1 _13492_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15231_ _15286_/A _15234_/B vssd1 vssd1 vccd1 vccd1 _15231_/X sky130_fd_sc_hd__or2_1
X_12443_ _12443_/A vssd1 vssd1 vccd1 vccd1 _12443_/Y sky130_fd_sc_hd__inv_6
XFILLER_173_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15162_ _15438_/A _15162_/B _15162_/C vssd1 vssd1 vccd1 vccd1 _15162_/X sky130_fd_sc_hd__and3_1
X_12374_ _18770_/Q _18769_/Q _12374_/C vssd1 vssd1 vccd1 vccd1 _12424_/C sky130_fd_sc_hd__and3_2
XFILLER_154_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17177__S _17177_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14113_ _18719_/Q _18718_/Q _18720_/Q _14453_/A vssd1 vssd1 vccd1 vccd1 _14462_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11325_ _11325_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11325_/X sky130_fd_sc_hd__or2_1
X_19970_ _20002_/CLK _19970_/D vssd1 vssd1 vccd1 vccd1 _19970_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16081__S _16089_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12147__A0 _15923_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15093_ _15405_/A vssd1 vssd1 vccd1 vccd1 _15093_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15884__A1 _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11256_ _19660_/Q _19426_/Q _18491_/Q _19756_/Q _11212_/X _11208_/X vssd1 vssd1 vccd1
+ vccd1 _11257_/B sky130_fd_sc_hd__mux4_2
X_14044_ _14044_/A _14044_/B _14044_/C vssd1 vssd1 vccd1 vccd1 _18590_/D sky130_fd_sc_hd__nor3_1
X_18921_ _18924_/CLK _18921_/D vssd1 vssd1 vccd1 vccd1 _18921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10207_ _10207_/A _10207_/B vssd1 vssd1 vccd1 vccd1 _10207_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11519__A _15962_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ _19228_/Q _19723_/Q _11295_/S vssd1 vssd1 vccd1 vccd1 _11187_/X sky130_fd_sc_hd__mux2_1
X_18852_ _18858_/CLK _18852_/D vssd1 vssd1 vccd1 vccd1 _18852_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11113__A1_N _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11370__A1 _11045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_151_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _10194_/A _10120_/X _10137_/X vssd1 vssd1 vccd1 vccd1 _10138_/X sky130_fd_sc_hd__a21bo_1
X_17803_ _17803_/A vssd1 vssd1 vccd1 vccd1 _19779_/D sky130_fd_sc_hd__clkbuf_1
X_18783_ _19910_/CLK _18783_/D vssd1 vssd1 vccd1 vccd1 _18783_/Q sky130_fd_sc_hd__dfxtp_1
X_15995_ _15995_/A vssd1 vssd1 vccd1 vccd1 _19028_/D sky130_fd_sc_hd__clkbuf_1
X_17734_ _17734_/A vssd1 vssd1 vccd1 vccd1 _19749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10069_ _10069_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _10069_/Y sky130_fd_sc_hd__nor2_1
X_14946_ _14943_/X _14944_/X _15014_/S vssd1 vssd1 vccd1 vccd1 _14946_/X sky130_fd_sc_hd__mux2_1
X_17665_ _17665_/A vssd1 vssd1 vccd1 vccd1 _17665_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15939__A2 _15921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14877_ _14877_/A vssd1 vssd1 vccd1 vccd1 _15355_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_165_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19404_ _19767_/CLK _19404_/D vssd1 vssd1 vccd1 vccd1 _19404_/Q sky130_fd_sc_hd__dfxtp_1
X_16616_ _16616_/A vssd1 vssd1 vccd1 vccd1 _19286_/D sky130_fd_sc_hd__clkbuf_1
X_13828_ _13828_/A vssd1 vssd1 vccd1 vccd1 _18507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17596_ _17596_/A vssd1 vssd1 vccd1 vccd1 _19701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10308__S0 _09655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19335_ _19828_/CLK _19335_/D vssd1 vssd1 vccd1 vccd1 _19335_/Q sky130_fd_sc_hd__dfxtp_1
X_16547_ _18208_/A _18352_/C vssd1 vssd1 vccd1 vccd1 _16604_/A sky130_fd_sc_hd__nor2_2
XANTENNA__16256__S _16258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ _13858_/S vssd1 vssd1 vccd1 vccd1 _13772_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__12622__A1 _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14565__A _14577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19266_ _20021_/CLK _19266_/D vssd1 vssd1 vccd1 vccd1 _19266_/Q sky130_fd_sc_hd__dfxtp_1
X_16478_ _19224_/Q _13754_/X _16486_/S vssd1 vssd1 vccd1 vccd1 _16479_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18217_ _19948_/Q _17646_/A _18219_/S vssd1 vssd1 vccd1 vccd1 _18218_/A sky130_fd_sc_hd__mux2_1
X_15429_ _15419_/X _15283_/X _15427_/X _15428_/X vssd1 vssd1 vccd1 vccd1 _15429_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19197_ _19950_/CLK _19197_/D vssd1 vssd1 vccd1 vccd1 _19197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_76_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11189__A1 _11157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18148_ _18148_/A vssd1 vssd1 vccd1 vccd1 _19917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11284__S1 _11077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18079_ _18079_/A vssd1 vssd1 vccd1 vccd1 _19895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09921_ _09614_/A _09920_/X _10073_/A vssd1 vssd1 vccd1 vccd1 _09921_/X sky130_fd_sc_hd__a21o_1
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09394__A _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13628__B _19009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17815__S _17821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ _09920_/S vssd1 vssd1 vccd1 vccd1 _11534_/S sky130_fd_sc_hd__clkbuf_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09783_ _09891_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09783_/X sky130_fd_sc_hd__or2_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17116__A _17199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10547__S0 _09653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16955__A _16977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11164__A _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15260__C1 _15951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09217_ _09217_/A vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__inv_2
XANTENNA__10508__A _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18381__S _18385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11275__S1 _10973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13819__A _17055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11110_ _19359_/Q _19694_/Q _11348_/S vssd1 vssd1 vccd1 vccd1 _11110_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12090_ _12091_/A _14914_/A vssd1 vssd1 vccd1 vccd1 _12092_/A sky130_fd_sc_hd__and2_1
XFILLER_1_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11041_ _11459_/A _12834_/A vssd1 vssd1 vccd1 vccd1 _11462_/B sky130_fd_sc_hd__nand2_4
XFILLER_150_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09640__S1 _09639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10560__C1 _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14800_ _14800_/A _14800_/B vssd1 vssd1 vccd1 vccd1 _14801_/A sky130_fd_sc_hd__and2_1
XANTENNA__17026__A _17026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _14750_/B _11867_/X _15779_/X _13885_/X vssd1 vssd1 vccd1 vccd1 _18958_/D
+ sky130_fd_sc_hd__o211a_1
X_12992_ _14278_/D _12889_/A _12989_/X _12991_/X vssd1 vssd1 vccd1 vccd1 _12992_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input13_A io_dbus_rdata[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ _14731_/A vssd1 vssd1 vccd1 vccd1 _18815_/D sky130_fd_sc_hd__clkbuf_1
X_11943_ _18968_/Q _12831_/A _11936_/X _11942_/Y vssd1 vssd1 vccd1 vccd1 _11943_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _17496_/S vssd1 vssd1 vccd1 vccd1 _17459_/S sky130_fd_sc_hd__buf_2
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _12799_/A _13742_/X _14667_/S vssd1 vssd1 vccd1 vccd1 _14663_/B sky130_fd_sc_hd__mux2_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _18637_/Q _09405_/B _13335_/B _18669_/Q vssd1 vssd1 vccd1 vccd1 _11874_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _16401_/A vssd1 vssd1 vccd1 vccd1 _19191_/D sky130_fd_sc_hd__clkbuf_1
X_13613_ _18878_/Q _13614_/B vssd1 vssd1 vccd1 vccd1 _13630_/C sky130_fd_sc_hd__or2_4
X_10825_ _11477_/A _10820_/Y _10822_/Y _10824_/Y vssd1 vssd1 vccd1 vccd1 _10825_/X
+ sky130_fd_sc_hd__a31o_1
X_17381_ _19602_/Q _17030_/X _17387_/S vssd1 vssd1 vccd1 vccd1 _17382_/A sky130_fd_sc_hd__mux2_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12604__A1 _12338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14593_ _14593_/A vssd1 vssd1 vccd1 vccd1 _18766_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14385__A _14385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19120_ _19583_/CLK _19120_/D vssd1 vssd1 vccd1 vccd1 _19120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16332_ _17668_/A vssd1 vssd1 vccd1 vccd1 _16332_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10615__B1 _09547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13544_ _14560_/A vssd1 vssd1 vccd1 vccd1 _13589_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09479__A _13307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ _10748_/A _10753_/X _10755_/X vssd1 vssd1 vccd1 vccd1 _10756_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19051_ _20033_/CLK _19051_/D vssd1 vssd1 vccd1 vccd1 _19051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16263_ _13238_/X _19144_/Q _16269_/S vssd1 vssd1 vccd1 vccd1 _16264_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11521__B _12855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18291__S _18291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13475_ _18895_/Q _13476_/B vssd1 vssd1 vccd1 vccd1 _13486_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16804__S _16808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10687_ _10680_/Y _10682_/Y _10684_/Y _10686_/Y _09820_/A vssd1 vssd1 vccd1 vccd1
+ _10687_/X sky130_fd_sc_hd__o221a_2
X_18002_ _18002_/A vssd1 vssd1 vccd1 vccd1 _19867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15214_ _15302_/A _15219_/A vssd1 vssd1 vccd1 vccd1 _15214_/X sky130_fd_sc_hd__or2_1
XFILLER_173_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12426_ _12422_/X _12423_/Y _12483_/C _12425_/X vssd1 vssd1 vccd1 vccd1 _12426_/Y
+ sky130_fd_sc_hd__o31ai_4
X_16194_ _16194_/A vssd1 vssd1 vccd1 vccd1 _19114_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15145_ _14830_/X _15135_/X _15144_/X _15089_/X vssd1 vssd1 vccd1 vccd1 _15145_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11040__B1 _09912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ _15321_/A _12357_/B vssd1 vssd1 vccd1 vccd1 _12360_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__15857__A1 _12082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output81_A _12521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15857__B2 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ _20012_/Q _19850_/Q _19259_/Q _19029_/Q _11155_/A _11108_/A vssd1 vssd1 vccd1
+ vccd1 _11309_/B sky130_fd_sc_hd__mux4_1
XFILLER_114_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19953_ _20017_/CLK _19953_/D vssd1 vssd1 vccd1 vccd1 _19953_/Q sky130_fd_sc_hd__dfxtp_1
X_15076_ _15099_/A vssd1 vssd1 vccd1 vccd1 _15366_/A sky130_fd_sc_hd__clkbuf_2
X_12288_ _12288_/A vssd1 vssd1 vccd1 vccd1 _12288_/X sky130_fd_sc_hd__buf_4
XFILLER_84_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18904_ _19001_/CLK _18904_/D vssd1 vssd1 vccd1 vccd1 _18904_/Q sky130_fd_sc_hd__dfxtp_1
X_14027_ _14026_/A _14026_/B _18584_/Q vssd1 vssd1 vccd1 vccd1 _14028_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__13332__A2 _13511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10153__A _10153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ _11296_/A _11238_/X _11340_/A vssd1 vssd1 vccd1 vccd1 _11239_/X sky130_fd_sc_hd__a21o_1
X_19884_ _19885_/CLK _19884_/D vssd1 vssd1 vccd1 vccd1 _19884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10777__S0 _10776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09942__A _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18835_ _18972_/CLK _18835_/D vssd1 vssd1 vccd1 vccd1 _18835_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11894__A2 _13189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18766_ _19899_/CLK _18766_/D vssd1 vssd1 vccd1 vccd1 _18766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15978_ _15978_/A _15978_/B _15978_/C vssd1 vssd1 vccd1 vccd1 _15978_/X sky130_fd_sc_hd__and3_1
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17717_ _17717_/A vssd1 vssd1 vccd1 vccd1 _17730_/S sky130_fd_sc_hd__buf_4
X_14929_ _12467_/A _15355_/B _14937_/S vssd1 vssd1 vccd1 vccd1 _14929_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18697_ _18744_/CLK _18697_/D vssd1 vssd1 vccd1 vccd1 _18697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17370__S _17376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17648_ _17648_/A vssd1 vssd1 vccd1 vccd1 _19722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13399__A2 _12889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17579_ _17579_/A vssd1 vssd1 vccd1 vccd1 _19693_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14295__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19318_ _20007_/CLK _19318_/D vssd1 vssd1 vccd1 vccd1 _19318_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12527__B _12556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14348__A1 _14350_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19249_ _19747_/CLK _19249_/D vssd1 vssd1 vccd1 vccd1 _19249_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16714__S _16714_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10909__A1 _10788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10047__B _12857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09904_ _19349_/Q _19620_/Q _19844_/Q _19588_/Q _11566_/S _09826_/A vssd1 vssd1 vccd1
+ vccd1 _09904_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20024_ _20024_/CLK _20024_/D vssd1 vssd1 vccd1 vccd1 _20024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09852__A _09920_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input5_A io_dbus_rdata[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09835_ _09833_/X _09834_/X _09942_/A vssd1 vssd1 vccd1 vccd1 _09835_/X sky130_fd_sc_hd__a21o_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09766_ _09942_/A vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13093__B _13093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _18827_/Q _09697_/B _09697_/C _09697_/D vssd1 vssd1 vccd1 vccd1 _09697_/X
+ sky130_fd_sc_hd__and4_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17280__S _17280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10845__B1 _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10670_/A _10610_/B vssd1 vssd1 vccd1 vccd1 _10610_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ _11626_/A _11589_/C _11589_/A vssd1 vssd1 vccd1 vccd1 _11591_/B sky130_fd_sc_hd__a21oi_1
XFILLER_22_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _19369_/Q _19704_/Q _10543_/S vssd1 vssd1 vccd1 vccd1 _10542_/B sky130_fd_sc_hd__mux2_1
XANTENNA__15536__B1 _15535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16624__S _16630_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13260_ _13068_/X _13255_/Y _13256_/X _13259_/X _13223_/A vssd1 vssd1 vccd1 vccd1
+ _13261_/B sky130_fd_sc_hd__o311a_1
X_10472_ _10207_/A _10469_/X _10471_/X vssd1 vssd1 vccd1 vccd1 _10472_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_136_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12211_ _15234_/A _12211_/B vssd1 vssd1 vccd1 vccd1 _12213_/A sky130_fd_sc_hd__xor2_1
XFILLER_170_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13191_ _18468_/Q _13511_/A _11847_/X _18692_/Q _13190_/X vssd1 vssd1 vccd1 vccd1
+ _13191_/X sky130_fd_sc_hd__a221o_1
XFILLER_163_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12142_ _12209_/B vssd1 vssd1 vccd1 vccd1 _15178_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_150_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12172__B _12234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17455__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13314__A2 _13070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16950_ _16950_/A vssd1 vssd1 vccd1 vccd1 _19433_/D sky130_fd_sc_hd__clkbuf_1
X_12073_ _13518_/A vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09762__A _10001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15901_ _18994_/Q _15900_/X _15901_/S vssd1 vssd1 vccd1 vccd1 _15902_/A sky130_fd_sc_hd__mux2_1
X_11024_ _11022_/X _11023_/X _09755_/A vssd1 vssd1 vccd1 vccd1 _11024_/Y sky130_fd_sc_hd__a21oi_1
X_16881_ _16345_/X _19403_/Q _16881_/S vssd1 vssd1 vccd1 vccd1 _16882_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15483__B _15487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11420__S1 _11208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11876__A2 _11869_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16298__C _16298_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15832_ _15832_/A vssd1 vssd1 vccd1 vccd1 _18972_/D sky130_fd_sc_hd__clkbuf_1
X_18620_ _18653_/CLK _18620_/D vssd1 vssd1 vccd1 vccd1 _18620_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10701__A _15947_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _18951_/Q _15775_/B vssd1 vssd1 vccd1 vccd1 _15763_/X sky130_fd_sc_hd__or2_1
X_18551_ _18745_/CLK _18551_/D vssd1 vssd1 vccd1 vccd1 _18551_/Q sky130_fd_sc_hd__dfxtp_1
X_12975_ _12936_/A _12971_/X _13015_/C _12974_/Y vssd1 vssd1 vccd1 vccd1 _12975_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17190__S _17193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__S0 _11171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _18808_/Q _11764_/X _14716_/S vssd1 vssd1 vccd1 vccd1 _14715_/A sky130_fd_sc_hd__mux2_1
X_17502_ _19657_/Q vssd1 vssd1 vccd1 vccd1 _17503_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_45_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15703__S _15703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _12587_/A _12033_/S vssd1 vssd1 vccd1 vccd1 _12175_/A sky130_fd_sc_hd__nor2_2
X_18482_ _18544_/CLK _18482_/D vssd1 vssd1 vccd1 vccd1 _18482_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ _15694_/A vssd1 vssd1 vccd1 vccd1 _18923_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15224__C1 _15951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17106_/X _19625_/Q _17437_/S vssd1 vssd1 vccd1 vccd1 _17434_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _18782_/Q _13704_/X _14649_/S vssd1 vssd1 vccd1 vccd1 _14646_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13731__B _13731_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _19006_/Q _11857_/B _11857_/C _11857_/D vssd1 vssd1 vccd1 vccd1 _11857_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_61_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10808_ _10009_/A _10805_/X _10807_/X vssd1 vssd1 vccd1 vccd1 _10808_/Y sky130_fd_sc_hd__a21oi_1
X_17364_ _17364_/A vssd1 vssd1 vccd1 vccd1 _19594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14576_ _12165_/A _13546_/X _14581_/S vssd1 vssd1 vccd1 vccd1 _14577_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11788_ _18756_/Q _14547_/A _13269_/A _18793_/Q _11787_/X vssd1 vssd1 vccd1 vccd1
+ _11788_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16315_ _16315_/A vssd1 vssd1 vccd1 vccd1 _19164_/D sky130_fd_sc_hd__clkbuf_1
X_19103_ _20016_/CLK _19103_/D vssd1 vssd1 vccd1 vccd1 _19103_/Q sky130_fd_sc_hd__dfxtp_1
X_13527_ _18457_/Q _13517_/X _16072_/B _13526_/Y vssd1 vssd1 vccd1 vccd1 _18457_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10739_ _10748_/A _10739_/B vssd1 vssd1 vccd1 vccd1 _10739_/Y sky130_fd_sc_hd__nor2_1
X_17295_ _17352_/S vssd1 vssd1 vccd1 vccd1 _17304_/S sky130_fd_sc_hd__buf_2
XFILLER_159_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18315__A _18337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19034_ _19567_/CLK _19034_/D vssd1 vssd1 vccd1 vccd1 _19034_/Q sky130_fd_sc_hd__dfxtp_1
X_16246_ _16246_/A vssd1 vssd1 vccd1 vccd1 _19136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13458_ _13458_/A _13731_/B vssd1 vssd1 vccd1 vccd1 _13458_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12409_ _12409_/A vssd1 vssd1 vccd1 vccd1 _12517_/S sky130_fd_sc_hd__buf_2
XFILLER_161_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16177_ _16177_/A vssd1 vssd1 vccd1 vccd1 _19106_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13389_ input19/X _13318_/X _13368_/X vssd1 vssd1 vccd1 vccd1 _13389_/Y sky130_fd_sc_hd__a21oi_1
Xoutput105 _14811_/A vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[2] sky130_fd_sc_hd__buf_2
Xoutput116 _12847_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[16] sky130_fd_sc_hd__buf_2
Xoutput127 _12858_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[26] sky130_fd_sc_hd__buf_2
Xoutput138 _12831_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[7] sky130_fd_sc_hd__buf_2
X_15128_ _15128_/A vssd1 vssd1 vccd1 vccd1 _18836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput149 _12454_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[16] sky130_fd_sc_hd__buf_2
XFILLER_5_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17365__S _17365_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19936_ _19936_/CLK _19936_/D vssd1 vssd1 vccd1 vccd1 _19936_/Q sky130_fd_sc_hd__dfxtp_1
X_15059_ _15057_/X _15058_/X _15199_/S vssd1 vssd1 vccd1 vccd1 _15059_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09672__A _09920_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19867_ _20031_/CLK _19867_/D vssd1 vssd1 vccd1 vccd1 _19867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09620_ _11140_/A vssd1 vssd1 vccd1 vccd1 _11006_/A sky130_fd_sc_hd__clkbuf_2
X_18818_ _18819_/CLK _18818_/D vssd1 vssd1 vccd1 vccd1 _18818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19798_ _19976_/CLK _19798_/D vssd1 vssd1 vccd1 vccd1 _19798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09551_ _09551_/A vssd1 vssd1 vccd1 vccd1 _10668_/A sky130_fd_sc_hd__buf_2
X_18749_ _19063_/CLK _18749_/D vssd1 vssd1 vccd1 vccd1 _18749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18196__S _18202_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__S0 _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09482_ _09480_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _11941_/B sky130_fd_sc_hd__and2b_2
XFILLER_37_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13241__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16444__S _16446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11004__B1 _11003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12273__A _12273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12504__A0 _12498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09582__A _10069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11402__S1 _11357_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20007_ _20007_/CLK _20007_/D vssd1 vssd1 vccd1 vccd1 _20007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09818_ _11166_/A vssd1 vssd1 vccd1 vccd1 _09819_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10521__A _10521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09749_ _19943_/Q _19557_/Q _20007_/Q _19126_/Q _09733_/X _09895_/A vssd1 vssd1 vccd1
+ vccd1 _09750_/B sky130_fd_sc_hd__mux4_1
XFILLER_36_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13832__A _17068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16846__C _16846_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12760_ _12760_/A vssd1 vssd1 vccd1 vccd1 _15531_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _18749_/Q _11677_/B _14555_/B _12452_/A _11710_/X vssd1 vssd1 vccd1 vccd1
+ _11711_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11653__C_N _11650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13551__B _13551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12729_/A _12645_/B _12670_/A _12690_/Y vssd1 vssd1 vccd1 vccd1 _12692_/B
+ sky130_fd_sc_hd__a31o_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13043__S _13116_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14433_/C _14431_/C _18704_/Q vssd1 vssd1 vccd1 vccd1 _14432_/B sky130_fd_sc_hd__a21oi_1
X_11642_ _11642_/A _11642_/B vssd1 vssd1 vccd1 vccd1 _11645_/B sky130_fd_sc_hd__or2_1
XFILLER_30_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10046__A1 _09884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14361_ _18683_/Q _18682_/Q _18681_/Q _18680_/Q vssd1 vssd1 vccd1 vccd1 _14363_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_35_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11573_ _11558_/A _11570_/X _11572_/X _09809_/X vssd1 vssd1 vccd1 vccd1 _11574_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 io_dbus_rdata[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_4
XFILLER_155_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16100_ _13115_/X _19073_/Q _16100_/S vssd1 vssd1 vccd1 vccd1 _16101_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12991__B1 _11791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ _18811_/Q _13071_/X _12984_/X _18778_/Q _13311_/X vssd1 vssd1 vccd1 vccd1
+ _13312_/X sky130_fd_sc_hd__a221o_2
Xinput29 io_dbus_rdata[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_156_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10524_ _10567_/A _10523_/X _09796_/A vssd1 vssd1 vccd1 vccd1 _10524_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_128_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17080_ _17080_/A vssd1 vssd1 vccd1 vccd1 _19479_/D sky130_fd_sc_hd__clkbuf_1
X_14292_ _14300_/D _14292_/B vssd1 vssd1 vccd1 vccd1 _18663_/D sky130_fd_sc_hd__nor2_1
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16031_ _13283_/X _19045_/Q _16031_/S vssd1 vssd1 vccd1 vccd1 _16032_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14732__A1 _13710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ _18882_/Q vssd1 vssd1 vccd1 vccd1 _13642_/A sky130_fd_sc_hd__clkbuf_2
X_10455_ _10415_/A _10454_/X _10192_/X vssd1 vssd1 vccd1 vccd1 _10455_/X sky130_fd_sc_hd__o21a_1
XFILLER_136_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09476__B _15942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13174_ _13174_/A _18878_/Q _13174_/C vssd1 vssd1 vccd1 vccd1 _13183_/B sky130_fd_sc_hd__and3_1
X_10386_ _19245_/Q _19740_/Q _10470_/S vssd1 vssd1 vccd1 vccd1 _10387_/B sky130_fd_sc_hd__mux2_1
XFILLER_112_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12125_ _12285_/A vssd1 vssd1 vccd1 vccd1 _12303_/B sky130_fd_sc_hd__clkbuf_2
X_17982_ _17982_/A vssd1 vssd1 vccd1 vccd1 _19858_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12911__A _14225_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13299__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15925__C _15925_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19721_ _20012_/CLK _19721_/D vssd1 vssd1 vccd1 vccd1 _19721_/Q sky130_fd_sc_hd__dfxtp_1
X_16933_ _16990_/S vssd1 vssd1 vccd1 vccd1 _16942_/S sky130_fd_sc_hd__clkbuf_4
X_12056_ _12154_/A vssd1 vssd1 vccd1 vccd1 _12056_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11849__A2 _11845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17913__S _17915_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _20017_/Q _19855_/Q _19264_/Q _19034_/Q _11048_/S _10978_/A vssd1 vssd1 vccd1
+ vccd1 _11007_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19652_ _20038_/CLK _19652_/D vssd1 vssd1 vccd1 vccd1 _19652_/Q sky130_fd_sc_hd__dfxtp_1
X_16864_ _16320_/X _19395_/Q _16870_/S vssd1 vssd1 vccd1 vccd1 _16865_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17985__A1 _17036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18603_ _20037_/CLK _18603_/D vssd1 vssd1 vccd1 vccd1 _18603_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14799__A1 _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15815_ _15883_/A vssd1 vssd1 vccd1 vccd1 _15831_/A sky130_fd_sc_hd__clkbuf_2
X_19583_ _19583_/CLK _19583_/D vssd1 vssd1 vccd1 vccd1 _19583_/Q sky130_fd_sc_hd__dfxtp_1
X_16795_ _16342_/X _19365_/Q _16797_/S vssd1 vssd1 vccd1 vccd1 _16796_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14838__A _14948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15746_ _09458_/A _15734_/X _15745_/X _15743_/X vssd1 vssd1 vccd1 vccd1 _18944_/D
+ sky130_fd_sc_hd__o211a_1
X_18534_ _19001_/CLK _18534_/D vssd1 vssd1 vccd1 vccd1 _18534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12958_ _12875_/X _13505_/B _12956_/Y _12957_/X vssd1 vssd1 vccd1 vccd1 _12958_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10904__S0 _10892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11909_ _13511_/B vssd1 vssd1 vccd1 vccd1 _14744_/B sky130_fd_sc_hd__buf_2
XFILLER_61_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18465_ _18526_/CLK _18465_/D vssd1 vssd1 vccd1 vccd1 _18465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15677_ _18916_/Q _18537_/Q _15677_/S vssd1 vssd1 vccd1 vccd1 _15678_/A sky130_fd_sc_hd__mux2_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _12889_/A vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17416_ _19618_/Q _17081_/X _17420_/S vssd1 vssd1 vccd1 vccd1 _17417_/A sky130_fd_sc_hd__mux2_1
X_14628_ _12562_/A _13667_/X _14632_/S vssd1 vssd1 vccd1 vccd1 _14629_/B sky130_fd_sc_hd__mux2_1
X_18396_ _17697_/X _20028_/Q _18396_/S vssd1 vssd1 vccd1 vccd1 _18397_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17347_ _17347_/A vssd1 vssd1 vccd1 vccd1 _19587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11234__B1 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14559_ _14559_/A vssd1 vssd1 vccd1 vccd1 _18757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09667__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _17195_/X _19557_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17279_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19017_ _19973_/CLK _19017_/D vssd1 vssd1 vccd1 vccd1 _19017_/Q sky130_fd_sc_hd__dfxtp_1
X_16229_ _16229_/A vssd1 vssd1 vccd1 vccd1 _19128_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14723__A1 _13685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13189__A _13189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17884__A _17952_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10606__A _10832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19919_ _20015_/CLK _19919_/D vssd1 vssd1 vccd1 vccd1 _19919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10199__S1 _10182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09603_ _10662_/A vssd1 vssd1 vccd1 vccd1 _10709_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14748__A _15762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11148__S0 _11017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ _09534_/A vssd1 vssd1 vccd1 vccd1 _19487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09465_ _12316_/A _12260_/A _09465_/C vssd1 vssd1 vccd1 vccd1 _09514_/C sky130_fd_sc_hd__or3_1
XFILLER_169_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09396_ _18952_/Q _18951_/Q _18949_/Q _18950_/Q vssd1 vssd1 vccd1 vccd1 _09403_/A
+ sky130_fd_sc_hd__or4b_2
XANTENNA__13798__S _13804_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10984__C1 _10983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09296__B _18939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14714__A1 _11764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15911__A0 _18997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10240_ _09884_/A _10229_/X _10238_/X _09913_/X _10239_/Y vssd1 vssd1 vccd1 vccd1
+ _12858_/B sky130_fd_sc_hd__o32a_4
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10171_ _19155_/Q _19416_/Q _19315_/Q _19650_/Q _10208_/A _10153_/A vssd1 vssd1 vccd1
+ vccd1 _10172_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17733__S _17736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13930_ _13938_/D vssd1 vssd1 vccd1 vccd1 _13936_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13861_ _14385_/A _18518_/Q _13861_/C vssd1 vssd1 vccd1 vccd1 _13862_/A sky130_fd_sc_hd__and3_1
XFILLER_47_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11139__S0 _11049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15600_ _13642_/A _18914_/Q _15600_/S vssd1 vssd1 vccd1 vccd1 _15601_/A sky130_fd_sc_hd__mux2_1
X_12812_ _12812_/A _12812_/B vssd1 vssd1 vccd1 vccd1 _12812_/Y sky130_fd_sc_hd__xnor2_4
X_16580_ _19270_/Q _13803_/X _16580_/S vssd1 vssd1 vccd1 vccd1 _16581_/A sky130_fd_sc_hd__mux2_1
X_13792_ _18496_/Q _13790_/X _13804_/S vssd1 vssd1 vccd1 vccd1 _13793_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15531_ _15531_/A _15531_/B vssd1 vssd1 vccd1 vccd1 _15531_/Y sky130_fd_sc_hd__nor2_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12743_ _12743_/A vssd1 vssd1 vccd1 vccd1 _12743_/Y sky130_fd_sc_hd__inv_6
XFILLER_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _19963_/Q _17694_/A _18252_/S vssd1 vssd1 vccd1 vccd1 _18251_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11799__B1_N _11730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _15366_/X _15459_/Y _15461_/X _14998_/X vssd1 vssd1 vccd1 vccd1 _15465_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12674_/A _12695_/C vssd1 vssd1 vccd1 vccd1 _12674_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__13205__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17201_/A _17201_/B vssd1 vssd1 vccd1 vccd1 _17202_/A sky130_fd_sc_hd__and2_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14413_/A _14419_/C vssd1 vssd1 vccd1 vccd1 _14413_/Y sky130_fd_sc_hd__nor2_1
X_18181_ _18181_/A vssd1 vssd1 vccd1 vccd1 _19932_/D sky130_fd_sc_hd__clkbuf_1
X_11625_ _11624_/Y _11515_/X _10653_/A _11595_/X vssd1 vssd1 vccd1 vccd1 _11628_/C
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11216__B1 _09559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14953__A1 _14996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15393_ _15393_/A vssd1 vssd1 vccd1 vccd1 _15506_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_168_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14393__A _14413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17132_ _17199_/S vssd1 vssd1 vccd1 vccd1 _17145_/S sky130_fd_sc_hd__buf_2
XANTENNA__11810__A _12918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14344_ _14345_/B _14364_/A _18679_/Q vssd1 vssd1 vccd1 vccd1 _14346_/B sky130_fd_sc_hd__a21oi_1
X_11556_ _11572_/A _11556_/B vssd1 vssd1 vccd1 vccd1 _11556_/X sky130_fd_sc_hd__or2_1
X_17063_ _19474_/Q _17062_/X _17072_/S vssd1 vssd1 vccd1 vccd1 _17064_/A sky130_fd_sc_hd__mux2_1
X_10507_ _20027_/Q _19865_/Q _19274_/Q _19044_/Q _10125_/S _10492_/A vssd1 vssd1 vccd1
+ vccd1 _10508_/B sky130_fd_sc_hd__mux4_1
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14705__A1 _13621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14275_ _18659_/Q _18658_/Q _18657_/Q _14275_/D vssd1 vssd1 vccd1 vccd1 _14287_/D
+ sky130_fd_sc_hd__and4_1
X_11487_ _11487_/A _11487_/B vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__and2_1
X_16014_ _13150_/X _19037_/Q _16020_/S vssd1 vssd1 vccd1 vccd1 _16015_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13226_ _13226_/A vssd1 vssd1 vccd1 vccd1 _13458_/A sky130_fd_sc_hd__clkbuf_2
X_10438_ _10438_/A _10438_/B vssd1 vssd1 vccd1 vccd1 _10438_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15936__B _15936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10860__S _11488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _13154_/X _13156_/X _13359_/B vssd1 vssd1 vccd1 vccd1 _13157_/X sky130_fd_sc_hd__mux2_1
X_10369_ _10369_/A _10369_/B vssd1 vssd1 vccd1 vccd1 _10369_/X sky130_fd_sc_hd__or2_1
XANTENNA__12641__A _12641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16113__A _16135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _12108_/A _12108_/B vssd1 vssd1 vccd1 vccd1 _12108_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _19851_/Q _17007_/X _17965_/S vssd1 vssd1 vccd1 vccd1 _17966_/A sky130_fd_sc_hd__mux2_1
X_13088_ _18873_/Q _13088_/B vssd1 vssd1 vccd1 vccd1 _13131_/C sky130_fd_sc_hd__and2_1
XANTENNA__11378__S0 _11212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19704_ _20024_/CLK _19704_/D vssd1 vssd1 vccd1 vccd1 _19704_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15952__A _15966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16916_ _16396_/X _19419_/Q _16918_/S vssd1 vssd1 vccd1 vccd1 _16917_/A sky130_fd_sc_hd__mux2_1
X_12039_ _12039_/A vssd1 vssd1 vccd1 vccd1 _12179_/S sky130_fd_sc_hd__clkbuf_2
X_17896_ _19820_/Q _17010_/X _17904_/S vssd1 vssd1 vccd1 vccd1 _17897_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11152__C1 _11166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18080__A0 _18848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19635_ _19989_/CLK _19635_/D vssd1 vssd1 vccd1 vccd1 _19635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16847_ _17635_/B vssd1 vssd1 vccd1 vccd1 _17954_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__15969__B1 _15955_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14568__A _14577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19566_ _19951_/CLK _19566_/D vssd1 vssd1 vccd1 vccd1 _19566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16778_ _16316_/X _19357_/Q _16786_/S vssd1 vssd1 vccd1 vccd1 _16779_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18517_ _19842_/CLK _18517_/D vssd1 vssd1 vccd1 vccd1 _18517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15729_ _16298_/C _15745_/B vssd1 vssd1 vccd1 vccd1 _15729_/X sky130_fd_sc_hd__or2_1
XFILLER_34_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19497_ _19693_/CLK _19497_/D vssd1 vssd1 vccd1 vccd1 _19497_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10353__S1 _09636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09250_ _09290_/A vssd1 vssd1 vccd1 vccd1 _09516_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18448_ _19583_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _09287_/A vssd1 vssd1 vccd1 vccd1 _09492_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__14944__A1 _15160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18379_ _17672_/X _20020_/Q _18385_/S vssd1 vssd1 vccd1 vccd1 _18380_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_146_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11758__B2 _12508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__A _14552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10966__C1 _11166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14750__B _14750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17119__A _17656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12551__A _12551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11167__A _18839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12486__A2 _12849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18071__A0 _18845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__A _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11694__B1 _11687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16169__S _16173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14478__A _14495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09517_ _14813_/A _14804_/C _14813_/B _11949_/B vssd1 vssd1 vccd1 vccd1 _09527_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_71_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _15147_/A vssd1 vssd1 vccd1 vccd1 _15942_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_158_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09379_ _15760_/A _11777_/B _11777_/C vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__or3_1
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11410_ _19352_/Q _19687_/Q _11410_/S vssd1 vssd1 vccd1 vccd1 _11410_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12390_ _12390_/A vssd1 vssd1 vccd1 vccd1 _12390_/Y sky130_fd_sc_hd__inv_6
XFILLER_166_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11341_ _20011_/Q _19849_/Q _19258_/Q _19028_/Q _11155_/A _11108_/A vssd1 vssd1 vccd1
+ vccd1 _11341_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14060_ _14062_/A _14062_/C _14059_/X vssd1 vssd1 vccd1 vccd1 _14060_/Y sky130_fd_sc_hd__a21oi_1
X_11272_ _19722_/Q vssd1 vssd1 vccd1 vccd1 _11272_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13011_ _18651_/Q _11815_/A _11794_/X _14142_/B vssd1 vssd1 vccd1 vccd1 _13011_/X
+ sky130_fd_sc_hd__a22o_1
X_10223_ _10223_/A vssd1 vssd1 vccd1 vccd1 _10223_/X sky130_fd_sc_hd__buf_2
XFILLER_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input43_A io_ibus_inst[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _18451_/Q _19480_/Q _19517_/Q _19091_/Q _10152_/X _10153_/X vssd1 vssd1 vccd1
+ vccd1 _10154_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11077__A _11077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17750_ _17750_/A vssd1 vssd1 vccd1 vccd1 _19755_/D sky130_fd_sc_hd__clkbuf_1
X_14962_ _14923_/X _14941_/Y _14961_/Y _15068_/A vssd1 vssd1 vccd1 vccd1 _14962_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10085_ _18448_/Q _19477_/Q _19514_/Q _19088_/Q _10095_/S _10028_/X vssd1 vssd1 vccd1
+ vccd1 _10085_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__buf_2
XANTENNA__09878__B1 _09540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701_ _19323_/Q _13768_/X _16703_/S vssd1 vssd1 vccd1 vccd1 _16702_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13913_ _18587_/Q _18586_/Q _18588_/Q _14029_/A vssd1 vssd1 vccd1 vccd1 _14037_/A
+ sky130_fd_sc_hd__and4_1
X_17681_ _17681_/A vssd1 vssd1 vccd1 vccd1 _17681_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14893_ _15016_/A vssd1 vssd1 vccd1 vccd1 _15202_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_63_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19420_ _19622_/CLK _19420_/D vssd1 vssd1 vccd1 vccd1 _19420_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11805__A _15762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13844_ _13844_/A vssd1 vssd1 vccd1 vccd1 _18512_/D sky130_fd_sc_hd__clkbuf_1
X_16632_ _16689_/S vssd1 vssd1 vccd1 vccd1 _16641_/S sky130_fd_sc_hd__buf_2
XANTENNA__13426__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12229__A2 _12012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19351_ _19622_/CLK _19351_/D vssd1 vssd1 vccd1 vccd1 _19351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13775_ _13858_/S vssd1 vssd1 vccd1 vccd1 _13788_/S sky130_fd_sc_hd__clkbuf_4
X_16563_ _19262_/Q _13778_/X _16569_/S vssd1 vssd1 vccd1 vccd1 _16564_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18294__S _18302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ _19663_/Q _19429_/Q _18494_/Q _19759_/Q _11121_/S _10973_/A vssd1 vssd1 vccd1
+ vccd1 _10988_/B sky130_fd_sc_hd__mux4_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18302_ _17665_/X _19986_/Q _18302_/S vssd1 vssd1 vccd1 vccd1 _18303_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12726_ _12750_/B _12750_/C vssd1 vssd1 vccd1 vccd1 _12726_/Y sky130_fd_sc_hd__nand2_1
X_15514_ _12717_/X _15458_/X _15513_/X _15454_/X vssd1 vssd1 vccd1 vccd1 _15514_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_149_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19282_ _19939_/CLK _19282_/D vssd1 vssd1 vccd1 vccd1 _19282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16494_ _16494_/A vssd1 vssd1 vccd1 vccd1 _19231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18233_ _19955_/Q _17668_/A _18241_/S vssd1 vssd1 vccd1 vccd1 _18234_/A sky130_fd_sc_hd__mux2_1
X_15445_ _15449_/A _15449_/B vssd1 vssd1 vccd1 vccd1 _15445_/Y sky130_fd_sc_hd__nand2_1
X_12657_ _12657_/A vssd1 vssd1 vccd1 vccd1 _12657_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12937__B1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10099__S0 _10277_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11608_ _11454_/Y _11608_/B _11608_/C vssd1 vssd1 vccd1 vccd1 _11608_/Y sky130_fd_sc_hd__nand3b_1
X_18164_ _18164_/A vssd1 vssd1 vccd1 vccd1 _19924_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15376_ _15365_/X _15348_/X _15375_/X _15324_/X vssd1 vssd1 vccd1 vccd1 _15376_/X
+ sky130_fd_sc_hd__a211o_1
X_12588_ _12588_/A vssd1 vssd1 vccd1 vccd1 _12682_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17638__S _17650_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14327_ _18673_/Q _14327_/B _14327_/C vssd1 vssd1 vccd1 vccd1 _14327_/X sky130_fd_sc_hd__and3_1
X_17115_ _17652_/A vssd1 vssd1 vccd1 vccd1 _17115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11539_ _19351_/Q _19622_/Q _19846_/Q _19590_/Q _09635_/X _09639_/X vssd1 vssd1 vccd1
+ vccd1 _11539_/X sky130_fd_sc_hd__mux4_2
XANTENNA__15947__A _15966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18095_ _18094_/X _19900_/Q _18095_/S vssd1 vssd1 vccd1 vccd1 _18096_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17046_ _17046_/A vssd1 vssd1 vccd1 vccd1 _17046_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14258_ _14279_/B _14264_/D vssd1 vssd1 vccd1 vccd1 _14259_/B sky130_fd_sc_hd__and2_1
XFILLER_172_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13209_ _19896_/Q _13209_/B vssd1 vssd1 vccd1 vccd1 _13209_/X sky130_fd_sc_hd__and2_1
XFILLER_143_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14189_ _14189_/A _14189_/B _14190_/B vssd1 vssd1 vccd1 vccd1 _18635_/D sky130_fd_sc_hd__nor3_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _18997_/CLK _18997_/D vssd1 vssd1 vccd1 vccd1 _18997_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_85_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _19844_/Q _17087_/X _17948_/S vssd1 vssd1 vccd1 vccd1 _17949_/A sky130_fd_sc_hd__mux2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_173_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19001_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_72_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17879_ _17879_/A vssd1 vssd1 vccd1 vccd1 _19813_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14298__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19618_ _19810_/CLK _19618_/D vssd1 vssd1 vccd1 vccd1 _19618_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11715__A _19010_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19549_ _19935_/CLK _19549_/D vssd1 vssd1 vccd1 vccd1 _19549_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_188_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19523_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16717__S _16725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09302_ _18978_/Q _18938_/Q vssd1 vssd1 vccd1 vccd1 _09302_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11979__A1 _14931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10100__B1 _09798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09233_ _11939_/A _14758_/A vssd1 vssd1 vccd1 vccd1 _09233_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10765__S _10872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18108__A1 _11879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19587_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12928__B1 _12879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09855__A _09855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_126_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _18918_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18379__S _18385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ _10200_/A _09997_/B vssd1 vssd1 vccd1 vccd1 _09997_/X sky130_fd_sc_hd__or2_1
XFILLER_89_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10014__S0 _10275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10910_ _19330_/Q _19601_/Q _19825_/Q _19569_/Q _10787_/A _10856_/A vssd1 vssd1 vccd1
+ vccd1 _10910_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11890_ _18478_/Q _12943_/A _11772_/A _18711_/Q vssd1 vssd1 vccd1 vccd1 _11890_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ _09547_/A _10830_/X _10839_/X _10078_/X _10840_/Y vssd1 vssd1 vccd1 vccd1
+ _15936_/B sky130_fd_sc_hd__o32a_4
XFILLER_44_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10317__S1 _10185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ _19001_/Q _13560_/B vssd1 vssd1 vccd1 vccd1 _13560_/X sky130_fd_sc_hd__or2_1
X_10772_ _10712_/X _10763_/X _10767_/X _10771_/X _09551_/A vssd1 vssd1 vccd1 vccd1
+ _10772_/X sky130_fd_sc_hd__a311o_1
XFILLER_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12511_ _12082_/X _14763_/C _12318_/Y vssd1 vssd1 vccd1 vccd1 _12511_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__14908__A1 _15474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ _18613_/Q vssd1 vssd1 vccd1 vccd1 _13924_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15230_ _15234_/A _15234_/B vssd1 vssd1 vccd1 vccd1 _15230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12442_ _12442_/A _12442_/B vssd1 vssd1 vccd1 vccd1 _12443_/A sky130_fd_sc_hd__xnor2_4
XFILLER_138_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15581__A1 _18905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15161_ _15159_/X _15154_/Y _15160_/Y vssd1 vssd1 vccd1 vccd1 _15162_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__16362__S _16362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _12349_/A _12374_/C _18770_/Q vssd1 vssd1 vccd1 vccd1 _12373_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_165_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14112_ _18714_/Q _18715_/Q _18717_/Q _18716_/Q vssd1 vssd1 vccd1 vccd1 _14453_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11324_ _19130_/Q _19391_/Q _19290_/Q _19625_/Q _11328_/A _11322_/A vssd1 vssd1 vccd1
+ vccd1 _11325_/B sky130_fd_sc_hd__mux4_1
XFILLER_154_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15092_ _18835_/Q _15053_/X _15090_/X _15091_/Y vssd1 vssd1 vccd1 vccd1 _18835_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14043_ _14042_/A _14042_/C _18590_/Q vssd1 vssd1 vccd1 vccd1 _14044_/C sky130_fd_sc_hd__a21oi_1
X_18920_ _18924_/CLK _18920_/D vssd1 vssd1 vccd1 vccd1 _18920_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14541__C1 _14540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11255_ _11003_/X _11248_/Y _11250_/Y _11252_/Y _11254_/Y vssd1 vssd1 vccd1 vccd1
+ _11255_/X sky130_fd_sc_hd__o32a_1
XANTENNA__10704__A _10704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13895__A1 _18537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ _19378_/Q _19713_/Q _10469_/S vssd1 vssd1 vccd1 vccd1 _10207_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_90_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 _19999_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_133_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11519__B _12853_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18851_ _18851_/CLK _18851_/D vssd1 vssd1 vccd1 vccd1 _18851_/Q sky130_fd_sc_hd__dfxtp_4
X_11186_ _19356_/Q _19691_/Q _11186_/S vssd1 vssd1 vccd1 vccd1 _11186_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18289__S _18291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17193__S _17193_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17802_ _17726_/X _19779_/Q _17804_/S vssd1 vssd1 vccd1 vccd1 _17803_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10137_ _10502_/A _10137_/B _10137_/C vssd1 vssd1 vccd1 vccd1 _10137_/X sky130_fd_sc_hd__or3_1
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18782_ _19910_/CLK _18782_/D vssd1 vssd1 vccd1 vccd1 _18782_/Q sky130_fd_sc_hd__dfxtp_1
X_15994_ _12963_/X _19028_/Q _15998_/S vssd1 vssd1 vccd1 vccd1 _15995_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17733_ _17732_/X _19749_/Q _17736_/S vssd1 vssd1 vccd1 vccd1 _17734_/A sky130_fd_sc_hd__mux2_1
X_10068_ _19937_/Q _19551_/Q _20001_/Q _19120_/Q _09918_/S _09646_/A vssd1 vssd1 vccd1
+ vccd1 _10069_/B sky130_fd_sc_hd__mux4_1
XFILLER_36_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14945_ _15029_/A vssd1 vssd1 vccd1 vccd1 _15014_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_36_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17664_ _17664_/A vssd1 vssd1 vccd1 vccd1 _19727_/D sky130_fd_sc_hd__clkbuf_1
X_14876_ _14867_/X _14874_/X _15117_/S vssd1 vssd1 vccd1 vccd1 _14876_/X sky130_fd_sc_hd__mux2_1
X_19403_ _20020_/CLK _19403_/D vssd1 vssd1 vccd1 vccd1 _19403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16615_ _19286_/Q _13854_/X _16617_/S vssd1 vssd1 vccd1 vccd1 _16616_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13827_ _18507_/Q _13826_/X _13836_/S vssd1 vssd1 vccd1 vccd1 _13828_/A sky130_fd_sc_hd__mux2_1
X_17595_ _17144_/X _19701_/Q _17595_/S vssd1 vssd1 vccd1 vccd1 _17596_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16537__S _16541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10308__S1 _10185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19334_ _19828_/CLK _19334_/D vssd1 vssd1 vccd1 vccd1 _19334_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12083__A0 _09466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13758_ _13839_/A vssd1 vssd1 vccd1 vccd1 _13858_/S sky130_fd_sc_hd__buf_8
X_16546_ _16546_/A vssd1 vssd1 vccd1 vccd1 _19255_/D sky130_fd_sc_hd__clkbuf_1
X_12709_ _15974_/B vssd1 vssd1 vccd1 vccd1 _12709_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19265_ _19569_/CLK _19265_/D vssd1 vssd1 vccd1 vccd1 _19265_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12366__A _12368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16477_ _16545_/S vssd1 vssd1 vccd1 vccd1 _16486_/S sky130_fd_sc_hd__buf_2
X_13689_ _11879_/X _13688_/Y _13689_/S vssd1 vssd1 vccd1 vccd1 _13689_/X sky130_fd_sc_hd__mux2_1
X_18216_ _18216_/A vssd1 vssd1 vccd1 vccd1 _19947_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15572__A1 _18901_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clock_A _18998_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15428_ _15428_/A vssd1 vssd1 vccd1 vccd1 _15428_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19196_ _19949_/CLK _19196_/D vssd1 vssd1 vccd1 vccd1 _19196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13583__A0 _13579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19636_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17368__S _17376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18147_ _17649_/X _19917_/Q _18147_/S vssd1 vssd1 vccd1 vccd1 _18148_/A sky130_fd_sc_hd__mux2_1
X_15359_ _15329_/X _15348_/X _15358_/X _15342_/X vssd1 vssd1 vccd1 vccd1 _15359_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16272__S _16280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18078_ _18077_/X _19895_/Q _18078_/S vssd1 vssd1 vccd1 vccd1 _18079_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09920_ _19380_/Q _19715_/Q _09920_/S vssd1 vssd1 vccd1 vccd1 _09920_/X sky130_fd_sc_hd__mux2_1
X_17029_ _17029_/A vssd1 vssd1 vccd1 vccd1 _19463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_58_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19994_/CLK sky130_fd_sc_hd__clkbuf_16
X_20040_ _20040_/CLK _20040_/D vssd1 vssd1 vccd1 vccd1 _20040_/Q sky130_fd_sc_hd__dfxtp_1
X_09851_ _09851_/A _09851_/B vssd1 vssd1 vccd1 vccd1 _09851_/X sky130_fd_sc_hd__and2_1
XFILLER_113_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13925__A _13946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09782_ _19222_/Q _19813_/Q _19975_/Q _19190_/Q _09733_/X _09768_/X vssd1 vssd1 vccd1
+ vccd1 _09783_/B sky130_fd_sc_hd__mux4_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16301__A _16400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10547__S1 _10587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17132__A _17199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13660__A _13660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11821__B1 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09216_ _09342_/B _09215_/X input33/X vssd1 vssd1 vccd1 vccd1 _09217_/A sky130_fd_sc_hd__o21bai_1
XFILLER_167_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13574__A0 _13572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17278__S _17280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16182__S _16184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09585__A _10980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10483__S0 _10279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16910__S _16914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11040_ _09881_/A _11030_/X _11039_/X _09912_/A _11011_/Y vssd1 vssd1 vccd1 vccd1
+ _12834_/A sky130_fd_sc_hd__o32a_4
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13835__A _17071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13629__B2 _19009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09928__S0 _09659_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _14034_/B _11682_/A _11791_/A _18554_/Q vssd1 vssd1 vccd1 vccd1 _12991_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17741__S _17749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11942_ _09504_/C _11937_/X _11940_/X _12536_/B vssd1 vssd1 vccd1 vccd1 _11942_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_55_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14730_ _18815_/Q _13704_/X _14738_/S vssd1 vssd1 vccd1 vccd1 _14731_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14661_ _14661_/A vssd1 vssd1 vccd1 vccd1 _18786_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _12060_/B _11772_/A _09405_/A _18701_/Q _11872_/X vssd1 vssd1 vccd1 vccd1
+ _11873_/X sky130_fd_sc_hd__a221o_2
XFILLER_60_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14666__A _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18138__A _18206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _16399_/X _19191_/Q _16400_/S vssd1 vssd1 vccd1 vccd1 _16401_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13570__A _19002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13612_ _13587_/X _13609_/X _13611_/Y _13590_/X _19007_/Q vssd1 vssd1 vccd1 vccd1
+ _13612_/X sky130_fd_sc_hd__a32o_4
X_10824_ _10824_/A _10824_/B vssd1 vssd1 vccd1 vccd1 _10824_/Y sky130_fd_sc_hd__nor2_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17042__A _17042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ _17380_/A vssd1 vssd1 vccd1 vccd1 _19601_/D sky130_fd_sc_hd__clkbuf_1
X_14592_ _14595_/A _14592_/B vssd1 vssd1 vccd1 vccd1 _14593_/A sky130_fd_sc_hd__and2_1
XANTENNA__11407__A3 _11406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10076__C1 _09555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16331_ _16331_/A vssd1 vssd1 vccd1 vccd1 _19169_/D sky130_fd_sc_hd__clkbuf_1
X_13543_ _13747_/A vssd1 vssd1 vccd1 vccd1 _14560_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10755_ _09759_/A _10754_/X _09794_/A vssd1 vssd1 vccd1 vccd1 _10755_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16262_ _16262_/A vssd1 vssd1 vccd1 vccd1 _19143_/D sky130_fd_sc_hd__clkbuf_1
X_19050_ _19839_/CLK _19050_/D vssd1 vssd1 vccd1 vccd1 _19050_/Q sky130_fd_sc_hd__dfxtp_1
X_13474_ _13188_/X _13472_/X _13473_/X _13268_/A vssd1 vssd1 vccd1 vccd1 _13474_/X
+ sky130_fd_sc_hd__o211a_1
X_10686_ _10680_/A _10685_/X _09777_/A vssd1 vssd1 vccd1 vccd1 _10686_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18001_ _19867_/Q _17058_/X _18009_/S vssd1 vssd1 vccd1 vccd1 _18002_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15213_ _15393_/A vssd1 vssd1 vccd1 vccd1 _15302_/A sky130_fd_sc_hd__clkbuf_2
X_12425_ _12583_/A vssd1 vssd1 vccd1 vccd1 _12425_/X sky130_fd_sc_hd__clkbuf_4
X_16193_ _13263_/X _19114_/Q _16195_/S vssd1 vssd1 vccd1 vccd1 _16194_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16092__S _16100_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12914__A _18938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09495__A _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15144_ _15071_/X _15137_/X _15143_/X _15491_/A vssd1 vssd1 vccd1 vccd1 _15144_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11040__A1 _09881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12356_ _12406_/A _12406_/B _12459_/A vssd1 vssd1 vccd1 vccd1 _12357_/B sky130_fd_sc_hd__o21ai_1
XFILLER_153_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15857__A2 _15856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11307_ _11242_/A _11304_/X _11306_/X vssd1 vssd1 vccd1 vccd1 _11307_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_153_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19952_ _19982_/CLK _19952_/D vssd1 vssd1 vccd1 vccd1 _19952_/Q sky130_fd_sc_hd__dfxtp_1
X_15075_ _14858_/X _15073_/X _15074_/X vssd1 vssd1 vccd1 vccd1 _15075_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10434__A _10434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ _12287_/A _12287_/B vssd1 vssd1 vccd1 vccd1 _12288_/A sky130_fd_sc_hd__and2_1
XFILLER_84_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14026_ _14026_/A _14026_/B _18584_/Q vssd1 vssd1 vccd1 vccd1 _14028_/B sky130_fd_sc_hd__and3_1
X_18903_ _19001_/CLK _18903_/D vssd1 vssd1 vccd1 vccd1 _18903_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output74_A _12335_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ _19357_/Q _19692_/Q _11348_/S vssd1 vssd1 vccd1 vccd1 _11238_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19883_ _19883_/CLK _19883_/D vssd1 vssd1 vccd1 vccd1 _19883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18834_ _19485_/CLK _18834_/D vssd1 vssd1 vccd1 vccd1 _18834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11169_ _15925_/C _12831_/B _15923_/C _12830_/B vssd1 vssd1 vccd1 vccd1 _11609_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18765_ _19899_/CLK _18765_/D vssd1 vssd1 vccd1 vccd1 _18765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15977_ _19022_/Q _14803_/X _15976_/X vssd1 vssd1 vccd1 vccd1 _19022_/D sky130_fd_sc_hd__a21o_1
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17716_ _17716_/A vssd1 vssd1 vccd1 vccd1 _17716_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15960__A _15964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14279__C _14279_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14928_ _15385_/B _15338_/B _14937_/S vssd1 vssd1 vccd1 vccd1 _14928_/X sky130_fd_sc_hd__mux2_1
X_18696_ _19888_/CLK _18696_/D vssd1 vssd1 vccd1 vccd1 _18696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17647_ _17646_/X _19722_/Q _17650_/S vssd1 vssd1 vccd1 vccd1 _17648_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16267__S _16269_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14859_ _14859_/A vssd1 vssd1 vccd1 vccd1 _15291_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13480__A _17090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17578_ _17119_/X _19693_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17579_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10067__C1 _09876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19317_ _20038_/CLK _19317_/D vssd1 vssd1 vccd1 vccd1 _19317_/Q sky130_fd_sc_hd__dfxtp_1
X_16529_ _16529_/A vssd1 vssd1 vccd1 vccd1 _19247_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11712__B _11712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19248_ _20032_/CLK _19248_/D vssd1 vssd1 vccd1 vccd1 _19248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19179_ _19706_/CLK _19179_/D vssd1 vssd1 vccd1 vccd1 _19179_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12824__A _12824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12543__B _14860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17826__S _17832_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16730__S _16736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ _09903_/A vssd1 vssd1 vccd1 vccd1 _11566_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12531__A1 _12508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20023_ _20023_/CLK _20023_/D vssd1 vssd1 vccd1 vccd1 _20023_/Q sky130_fd_sc_hd__dfxtp_1
X_09834_ _19254_/Q _19749_/Q _09898_/S vssd1 vssd1 vccd1 vccd1 _09834_/X sky130_fd_sc_hd__mux2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _09765_/A vssd1 vssd1 vccd1 vccd1 _09942_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12819__C1 _13650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16966__A _16977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09696_ _09696_/A _09696_/B _09696_/C vssd1 vssd1 vccd1 vccd1 _09697_/D sky130_fd_sc_hd__and3_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10845__A1 _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15784__A1 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09999__C1 _09555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18392__S _18396_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _10540_/A _10540_/B vssd1 vssd1 vccd1 vccd1 _11592_/A sky130_fd_sc_hd__nor2_1
XANTENNA__15536__A1 _12766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_194_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10471_ _10424_/A _10470_/X _10376_/A vssd1 vssd1 vccd1 vccd1 _10471_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10953__S _10953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13011__A2 _11815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12210_ _12322_/A _12323_/A vssd1 vssd1 vccd1 vccd1 _12211_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13190_ _19895_/Q _13373_/B vssd1 vssd1 vccd1 vccd1 _13190_/X sky130_fd_sc_hd__and2_1
XFILLER_68_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17736__S _17736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ _12174_/A _12830_/B _12175_/A _09261_/A vssd1 vssd1 vccd1 vccd1 _12209_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10254__A _10254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12072_ _12070_/Y _12071_/X _12059_/X vssd1 vssd1 vccd1 vccd1 _12072_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15900_ _15899_/B _11967_/Y _11935_/X _15899_/Y vssd1 vssd1 vccd1 vccd1 _15900_/X
+ sky130_fd_sc_hd__o22a_2
X_11023_ _19360_/Q _19695_/Q _11023_/S vssd1 vssd1 vccd1 vccd1 _11023_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16880_ _16880_/A vssd1 vssd1 vccd1 vccd1 _19402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15831_ _15831_/A _15831_/B vssd1 vssd1 vccd1 vccd1 _15832_/A sky130_fd_sc_hd__and2_1
XFILLER_77_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10701__B _12844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18550_ _18745_/CLK _18550_/D vssd1 vssd1 vccd1 vccd1 _18550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _15762_/A vssd1 vssd1 vccd1 vccd1 _15775_/B sky130_fd_sc_hd__clkbuf_1
X_12974_ _13504_/A _12973_/B _13307_/A vssd1 vssd1 vccd1 vccd1 _12974_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09334__B_N _17098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17501_ _17501_/A vssd1 vssd1 vccd1 vccd1 _19656_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11184__S1 _11172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _14713_/A vssd1 vssd1 vccd1 vccd1 _18807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _11951_/A _11925_/B _09436_/C vssd1 vssd1 vccd1 vccd1 _12587_/A sky130_fd_sc_hd__nor3b_4
X_18481_ _18544_/CLK _18481_/D vssd1 vssd1 vccd1 vccd1 _18481_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output112_A _12841_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16087__S _16089_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15693_ _18923_/Q _18544_/Q _15699_/S vssd1 vssd1 vccd1 vccd1 _15694_/A sky130_fd_sc_hd__mux2_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _17432_/A vssd1 vssd1 vccd1 vccd1 _19624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11813__A _13656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14644_ _14644_/A vssd1 vssd1 vccd1 vccd1 _18781_/D sky130_fd_sc_hd__clkbuf_1
X_11856_ _18658_/Q _11815_/X _13189_/A _18562_/Q _11855_/X vssd1 vssd1 vccd1 vccd1
+ _11857_/D sky130_fd_sc_hd__a221o_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ _09830_/A _10806_/X _11493_/A vssd1 vssd1 vccd1 vccd1 _10807_/X sky130_fd_sc_hd__a21o_1
X_14575_ _14575_/A vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__clkbuf_1
X_17363_ _19594_/Q _17004_/X _17365_/S vssd1 vssd1 vccd1 vccd1 _17364_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15004__B _15004_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16815__S _16819_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10429__A _10434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11787_ _18681_/Q _11819_/A _11671_/A _18746_/Q _11786_/X vssd1 vssd1 vccd1 vccd1
+ _11787_/X sky130_fd_sc_hd__a221o_1
X_19102_ _20015_/CLK _19102_/D vssd1 vssd1 vccd1 vccd1 _19102_/Q sky130_fd_sc_hd__dfxtp_1
X_16314_ _16313_/X _19164_/Q _16314_/S vssd1 vssd1 vccd1 vccd1 _16315_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11261__A1 _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10738_ _19927_/Q _19541_/Q _19991_/Q _19110_/Q _09725_/A _10009_/A vssd1 vssd1 vccd1
+ vccd1 _10739_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13526_ _13526_/A _13526_/B vssd1 vssd1 vccd1 vccd1 _13526_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17294_ _17294_/A vssd1 vssd1 vccd1 vccd1 _19563_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13538__A0 hold7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19033_ _19949_/CLK _19033_/D vssd1 vssd1 vccd1 vccd1 _19033_/Q sky130_fd_sc_hd__dfxtp_1
X_16245_ _13098_/X _19136_/Q _16247_/S vssd1 vssd1 vccd1 vccd1 _16246_/A sky130_fd_sc_hd__mux2_1
X_13457_ _18579_/Q _13070_/X _13453_/X _13455_/X _13456_/X vssd1 vssd1 vccd1 vccd1
+ _13731_/B sky130_fd_sc_hd__a2111o_2
XFILLER_173_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10669_ _19928_/Q _19542_/Q _19992_/Q _19111_/Q _10586_/S _10656_/A vssd1 vssd1 vccd1
+ vccd1 _10670_/B sky130_fd_sc_hd__mux4_1
XFILLER_139_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12408_ _15355_/A _12408_/B vssd1 vssd1 vccd1 vccd1 _12411_/A sky130_fd_sc_hd__xnor2_4
XFILLER_12_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16176_ _13137_/X _19106_/Q _16184_/S vssd1 vssd1 vccd1 vccd1 _16177_/A sky130_fd_sc_hd__mux2_1
X_13388_ _13388_/A vssd1 vssd1 vccd1 vccd1 _18449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput106 _14782_/A vssd1 vssd1 vccd1 vccd1 io_dbus_rd_en sky130_fd_sc_hd__buf_2
XFILLER_154_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput117 _12848_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[17] sky130_fd_sc_hd__buf_2
XFILLER_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15955__A _15955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput128 _12861_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[27] sky130_fd_sc_hd__buf_2
X_12339_ _12340_/A _12340_/C _12340_/B vssd1 vssd1 vccd1 vccd1 _12341_/A sky130_fd_sc_hd__a21oi_1
X_15127_ _18836_/Q _15126_/X _15127_/S vssd1 vssd1 vccd1 vccd1 _15128_/A sky130_fd_sc_hd__mux2_1
Xoutput139 _12834_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[8] sky130_fd_sc_hd__buf_2
XANTENNA__16550__S _16558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19935_ _19935_/CLK _19935_/D vssd1 vssd1 vccd1 vccd1 _19935_/Q sky130_fd_sc_hd__dfxtp_1
X_15058_ _14930_/X _14882_/X _15118_/S vssd1 vssd1 vccd1 vccd1 _15058_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _18578_/Q _14013_/C vssd1 vssd1 vccd1 vccd1 _14010_/B sky130_fd_sc_hd__and2_1
XFILLER_68_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19866_ _19972_/CLK _19866_/D vssd1 vssd1 vccd1 vccd1 _19866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18817_ _19910_/CLK _18817_/D vssd1 vssd1 vccd1 vccd1 _18817_/Q sky130_fd_sc_hd__dfxtp_1
X_19797_ _19959_/CLK _19797_/D vssd1 vssd1 vccd1 vccd1 _19797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17381__S _17387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09550_ _09550_/A vssd1 vssd1 vccd1 vccd1 _09551_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15690__A _15690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18748_ _19063_/CLK _18748_/D vssd1 vssd1 vccd1 vccd1 _18748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11175__S1 _11015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ _09481_/A _09481_/B _09481_/C _09481_/D vssd1 vssd1 vccd1 vccd1 _09482_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__09693__A1 _09862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18679_ _18687_/CLK _18679_/D vssd1 vssd1 vccd1 vccd1 _18679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11723__A _11831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12538__B _12851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16725__S _16725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12837__A_N _12833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12554__A _12554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16460__S _16468_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13701__B1 _13700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20006_ _20006_/CLK _20006_/D vssd1 vssd1 vccd1 vccd1 _20006_/Q sky130_fd_sc_hd__dfxtp_1
X_09817_ _09817_/A vssd1 vssd1 vccd1 vccd1 _11166_/A sky130_fd_sc_hd__buf_2
XFILLER_74_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17291__S _17293_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _09940_/A vssd1 vssd1 vccd1 vccd1 _09895_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _10069_/A _09679_/B vssd1 vssd1 vccd1 vccd1 _09679_/X sky130_fd_sc_hd__or2_1
XFILLER_43_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13324__S _13366_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ _18470_/Q _12943_/A _14672_/A _18806_/Q _11709_/X vssd1 vssd1 vccd1 vccd1
+ _11710_/X sky130_fd_sc_hd__a221o_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15757__A1 _12082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12640_/A _12666_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _12690_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11491__B2 _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11524_/A _10301_/A _11634_/B _10106_/Y _11642_/A vssd1 vssd1 vccd1 vccd1
+ _11645_/A sky130_fd_sc_hd__a311o_1
XFILLER_14_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14360_ _18684_/Q _14356_/C _18685_/Q vssd1 vssd1 vccd1 vccd1 _14365_/B sky130_fd_sc_hd__a21oi_1
XFILLER_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11572_ _11572_/A _11572_/B vssd1 vssd1 vccd1 vccd1 _11572_/X sky130_fd_sc_hd__or2_1
XANTENNA__12586__A4 _15436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13311_ _18475_/Q _11755_/X _11847_/A _18699_/Q _13310_/X vssd1 vssd1 vccd1 vccd1
+ _13311_/X sky130_fd_sc_hd__a221o_1
XFILLER_168_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10523_ _19210_/Q _19801_/Q _19963_/Q _19178_/Q _10521_/X _10522_/X vssd1 vssd1 vccd1
+ vccd1 _10523_/X sky130_fd_sc_hd__mux4_1
Xinput19 io_dbus_rdata[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_6
XFILLER_7_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ _18663_/Q _14297_/D _14792_/A vssd1 vssd1 vccd1 vccd1 _14292_/B sky130_fd_sc_hd__o21ai_1
XFILLER_167_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16030_ _16030_/A vssd1 vssd1 vccd1 vccd1 _19044_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14193__B1 _14160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13242_ _18882_/Q _13256_/C vssd1 vssd1 vccd1 vccd1 _13267_/C sky130_fd_sc_hd__and2_1
X_10454_ _19339_/Q _19610_/Q _19834_/Q _19578_/Q _09995_/A _10400_/A vssd1 vssd1 vccd1
+ vccd1 _10454_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17466__S _17470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10203__C1 _09876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13173_ _13174_/A _13174_/C _18878_/Q vssd1 vssd1 vccd1 vccd1 _13175_/B sky130_fd_sc_hd__a21oi_1
X_10385_ _19676_/Q _19442_/Q _18507_/Q _19772_/Q _10209_/S _09745_/A vssd1 vssd1 vccd1
+ vccd1 _10385_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12124_ _12215_/C _12124_/B vssd1 vssd1 vccd1 vccd1 _12124_/X sky130_fd_sc_hd__xor2_4
X_17981_ _19858_/Q _17030_/X _17987_/S vssd1 vssd1 vccd1 vccd1 _17982_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19720_ _19720_/CLK _19720_/D vssd1 vssd1 vccd1 vccd1 _19720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12055_ _12055_/A _12055_/B _12055_/C _09471_/X vssd1 vssd1 vccd1 vccd1 _12154_/A
+ sky130_fd_sc_hd__nor4b_1
X_16932_ _16932_/A vssd1 vssd1 vccd1 vccd1 _19425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10712__A _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__B1 _10107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11006_ _11006_/A _11006_/B vssd1 vssd1 vccd1 vccd1 _11006_/Y sky130_fd_sc_hd__nor2_1
X_19651_ _19973_/CLK _19651_/D vssd1 vssd1 vccd1 vccd1 _19651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16863_ _16863_/A vssd1 vssd1 vccd1 vccd1 _19394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18602_ _20037_/CLK _18602_/D vssd1 vssd1 vccd1 vccd1 _18602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15814_ _15814_/A vssd1 vssd1 vccd1 vccd1 _18967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19582_ _20030_/CLK _19582_/D vssd1 vssd1 vccd1 vccd1 _19582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16794_ _16794_/A vssd1 vssd1 vccd1 vccd1 _19364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18533_ _18867_/CLK _18533_/D vssd1 vssd1 vccd1 vccd1 _18533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _18944_/Q _15745_/B vssd1 vssd1 vccd1 vccd1 _15745_/X sky130_fd_sc_hd__or2_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _12957_/A vssd1 vssd1 vccd1 vccd1 _12957_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13471__A2 _13120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ _12827_/A _14771_/A vssd1 vssd1 vccd1 vccd1 _11908_/Y sky130_fd_sc_hd__nor2_4
X_18464_ _18526_/CLK _18464_/D vssd1 vssd1 vccd1 vccd1 _18464_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ _15676_/A vssd1 vssd1 vccd1 vccd1 _18915_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _18582_/Q _11732_/X _12887_/X _18614_/Q vssd1 vssd1 vccd1 vccd1 _12888_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17415_ _17415_/A vssd1 vssd1 vccd1 vccd1 _19617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14627_ _14627_/A vssd1 vssd1 vccd1 vccd1 _18776_/D sky130_fd_sc_hd__clkbuf_1
X_18395_ _18395_/A vssd1 vssd1 vccd1 vccd1 _20027_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10159__A _10382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16545__S _16545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11839_ _12060_/B _14792_/B _11833_/X _11838_/X vssd1 vssd1 vccd1 vccd1 _18712_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18326__A _18337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ _17189_/X _19587_/Q _17348_/S vssd1 vssd1 vccd1 vccd1 _17347_/A sky130_fd_sc_hd__mux2_1
X_14558_ _15833_/A _14558_/B vssd1 vssd1 vccd1 vccd1 _14559_/A sky130_fd_sc_hd__or2_1
XANTENNA__14971__A2 _12812_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13509_ _13648_/A _13504_/Y _16069_/B vssd1 vssd1 vccd1 vccd1 _13509_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17277_ _17277_/A vssd1 vssd1 vccd1 vccd1 _19556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14489_ _14514_/A _14493_/C vssd1 vssd1 vccd1 vccd1 _14489_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19016_ _19973_/CLK _19016_/D vssd1 vssd1 vccd1 vccd1 _19016_/Q sky130_fd_sc_hd__dfxtp_1
X_16228_ _12909_/X _19128_/Q _16236_/S vssd1 vssd1 vccd1 vccd1 _16229_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12195__C1 _12154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17376__S _17376_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12734__A1 _09471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16280__S _16280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16159_ _16159_/A vssd1 vssd1 vccd1 vccd1 _19098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19918_ _19982_/CLK _19918_/D vssd1 vssd1 vccd1 vccd1 _19918_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10622__A _11486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_142_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19849_ _19947_/CLK _19849_/D vssd1 vssd1 vccd1 vccd1 _19849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09602_ _11050_/A vssd1 vssd1 vccd1 vccd1 _10662_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09533_ _09532_/X _14782_/A _15127_/S vssd1 vssd1 vccd1 vccd1 _09534_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11148__S1 _11015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09464_ _18991_/Q vssd1 vssd1 vccd1 vccd1 _12260_/A sky130_fd_sc_hd__buf_4
XFILLER_145_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09395_ _11777_/C _09407_/C vssd1 vssd1 vccd1 vccd1 _11671_/A sky130_fd_sc_hd__nor2_4
XANTENNA__16455__S _16457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10069__A _10069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13214__A2 _11732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_67_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17113__A0 _17112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10736__B1 _10078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09593__A _10493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10831__S0 _11467_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ _19347_/Q _19618_/Q _19842_/Q _19586_/Q _10152_/X _10153_/X vssd1 vssd1 vccd1
+ vccd1 _10170_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _16836_/A vssd1 vssd1 vccd1 vccd1 _14385_/A sky130_fd_sc_hd__buf_4
XFILLER_75_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11139__S1 _10973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _12811_/A _12811_/B vssd1 vssd1 vccd1 vccd1 _12812_/B sky130_fd_sc_hd__xnor2_2
X_13791_ _13858_/S vssd1 vssd1 vccd1 vccd1 _13804_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__12459__A _12459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13453__A2 _13071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _15077_/X _15527_/Y _15529_/X _15216_/X vssd1 vssd1 vccd1 vccd1 _15530_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_103_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12742_/A _12742_/B vssd1 vssd1 vccd1 vccd1 _12743_/A sky130_fd_sc_hd__xnor2_4
XFILLER_16_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12790_/A vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__buf_2
X_15461_ _15368_/X _15463_/B _15369_/X _15460_/X vssd1 vssd1 vccd1 vccd1 _15461_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14674__A _14742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13205__A2 _13091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17200_/A vssd1 vssd1 vccd1 vccd1 _19521_/D sky130_fd_sc_hd__clkbuf_1
X_11624_ _11624_/A vssd1 vssd1 vccd1 vccd1 _11624_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _14422_/D vssd1 vssd1 vccd1 vccd1 _14419_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18180_ _17697_/X _19932_/Q _18180_/S vssd1 vssd1 vccd1 vccd1 _18181_/A sky130_fd_sc_hd__mux2_1
X_15392_ _15397_/A _15397_/B vssd1 vssd1 vccd1 vccd1 _15392_/Y sky130_fd_sc_hd__nand2_1
X_17131_ _17668_/A vssd1 vssd1 vccd1 vccd1 _17131_/X sky130_fd_sc_hd__clkbuf_2
X_11555_ _19944_/Q _19558_/Q _20008_/Q _19127_/Q _11553_/X _11565_/A vssd1 vssd1 vccd1
+ vccd1 _11556_/B sky130_fd_sc_hd__mux4_1
X_14343_ _14345_/B _14364_/A _14342_/Y vssd1 vssd1 vccd1 vccd1 _18678_/D sky130_fd_sc_hd__o21a_1
XFILLER_7_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10506_ _09988_/A _10505_/X _10107_/A vssd1 vssd1 vccd1 vccd1 _10506_/Y sky130_fd_sc_hd__o21ai_1
X_17062_ _17062_/A vssd1 vssd1 vccd1 vccd1 _17062_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14274_ _18658_/Q _14270_/B _14273_/Y vssd1 vssd1 vccd1 vccd1 _18658_/D sky130_fd_sc_hd__o21a_1
X_11486_ _19365_/Q _19700_/Q _11486_/S vssd1 vssd1 vccd1 vccd1 _11487_/B sky130_fd_sc_hd__mux2_1
XFILLER_171_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16013_ _16013_/A vssd1 vssd1 vccd1 vccd1 _19036_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17196__S _17199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13225_ _13207_/A _13224_/C _18881_/Q vssd1 vssd1 vccd1 vccd1 _13225_/Y sky130_fd_sc_hd__a21oi_1
X_10437_ _19212_/Q _19803_/Q _19965_/Q _19180_/Q _10328_/S _10027_/A vssd1 vssd1 vccd1
+ vccd1 _10438_/B sky130_fd_sc_hd__mux4_1
XANTENNA__17104__A0 _17103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12922__A _13386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13156_ _13174_/A _13174_/C vssd1 vssd1 vccd1 vccd1 _13156_/X sky130_fd_sc_hd__xor2_1
X_10368_ _19213_/Q _19804_/Q _19966_/Q _19181_/Q _10058_/A _10261_/A vssd1 vssd1 vccd1
+ vccd1 _10369_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15666__A0 _18911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12107_/A _12107_/B vssd1 vssd1 vccd1 vccd1 _12108_/B sky130_fd_sc_hd__nand2_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17924__S _17926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11538__A _11538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _17964_/A vssd1 vssd1 vccd1 vccd1 _19850_/D sky130_fd_sc_hd__clkbuf_1
X_13087_ _13580_/A _13088_/B vssd1 vssd1 vccd1 vccd1 _13089_/B sky130_fd_sc_hd__nor2_1
X_10299_ _18856_/Q _09843_/X _09884_/X _10298_/X vssd1 vssd1 vccd1 vccd1 _12855_/B
+ sky130_fd_sc_hd__o2bb2a_4
X_19703_ _19960_/CLK _19703_/D vssd1 vssd1 vccd1 vccd1 _19703_/Q sky130_fd_sc_hd__dfxtp_1
X_16915_ _16915_/A vssd1 vssd1 vccd1 vccd1 _19418_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11378__S1 _11077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ _12038_/A _15103_/B vssd1 vssd1 vccd1 vccd1 _12042_/A sky130_fd_sc_hd__xnor2_1
XFILLER_78_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15952__B _15966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17895_ _17952_/S vssd1 vssd1 vccd1 vccd1 _17904_/S sky130_fd_sc_hd__buf_2
XFILLER_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19634_ _19637_/CLK _19634_/D vssd1 vssd1 vccd1 vccd1 _19634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18080__A1 _13629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16846_ _18937_/Q _16846_/B _16846_/C vssd1 vssd1 vccd1 vccd1 _17635_/B sky130_fd_sc_hd__or3_2
XFILLER_38_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19565_ _19951_/CLK _19565_/D vssd1 vssd1 vccd1 vccd1 _19565_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10588__S _10657_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16777_ _16834_/S vssd1 vssd1 vccd1 vccd1 _16786_/S sky130_fd_sc_hd__buf_2
XFILLER_93_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13989_ _18570_/Q _13990_/C _18571_/Q vssd1 vssd1 vccd1 vccd1 _13991_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11273__A _11273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18516_ _20039_/CLK _18516_/D vssd1 vssd1 vccd1 vccd1 _18516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ _16150_/B vssd1 vssd1 vccd1 vccd1 _16298_/C sky130_fd_sc_hd__buf_4
X_19496_ _20017_/CLK _19496_/D vssd1 vssd1 vccd1 vccd1 _19496_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12088__B _15183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18447_ _19936_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17591__A0 _17138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15659_ _15659_/A vssd1 vssd1 vccd1 vccd1 _18907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14584__A _14601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ _11919_/B _09282_/C _09311_/A vssd1 vssd1 vccd1 vccd1 _09287_/A sky130_fd_sc_hd__or3_1
X_18378_ _18378_/A vssd1 vssd1 vccd1 vccd1 _20019_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17329_ _17163_/X _19579_/Q _17337_/S vssd1 vssd1 vccd1 vccd1 _17330_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17895__A _17952_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11066__S0 _11063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13139__S _13203_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14759__A _15393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__B1 _09537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18071__A1 _11860_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12891__B1 _12890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14632__A1 _13677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14197__C _14197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09516_ _09516_/A _09516_/B vssd1 vssd1 vccd1 vccd1 _11949_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11614__C _11614_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _14665_/A _14771_/B vssd1 vssd1 vccd1 vccd1 _15147_/A sky130_fd_sc_hd__nand2_4
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13199__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ _09378_/A _14227_/A vssd1 vssd1 vccd1 vccd1 _11777_/C sky130_fd_sc_hd__or2_2
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10527__A _10572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11340_ _11340_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11340_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14699__A1 _11833_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13838__A _17074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11271_ _10983_/X _11270_/X _11425_/A vssd1 vssd1 vccd1 vccd1 _11271_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_153_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13010_ _18619_/Q vssd1 vssd1 vccd1 vccd1 _14142_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10222_ _10480_/A vssd1 vssd1 vccd1 vccd1 _10344_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _10153_/A vssd1 vssd1 vccd1 vccd1 _10153_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10280__S1 _10329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13123__A1 _18464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10084_ _10093_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10084_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_input36_A io_ibus_inst[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ _15165_/S _14951_/X _14960_/X vssd1 vssd1 vccd1 vccd1 _14961_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09878__B2 _18862_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16700_ _16700_/A vssd1 vssd1 vccd1 vccd1 _19322_/D sky130_fd_sc_hd__clkbuf_1
X_13912_ _18582_/Q _18583_/Q _18585_/Q _18584_/Q vssd1 vssd1 vccd1 vccd1 _14029_/A
+ sky130_fd_sc_hd__and4_1
X_17680_ _17680_/A vssd1 vssd1 vccd1 vccd1 _19732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14892_ _12753_/A _11981_/Y _11985_/X vssd1 vssd1 vccd1 vccd1 _15016_/A sky130_fd_sc_hd__o21ai_4
XFILLER_48_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16631_ _16631_/A vssd1 vssd1 vccd1 vccd1 _19292_/D sky130_fd_sc_hd__clkbuf_1
X_13843_ _18512_/Q _13842_/X _13852_/S vssd1 vssd1 vccd1 vccd1 _13844_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19350_ _19350_/CLK _19350_/D vssd1 vssd1 vccd1 vccd1 _19350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16562_ _16562_/A vssd1 vssd1 vccd1 vccd1 _19261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10986_ _11212_/A vssd1 vssd1 vccd1 vccd1 _11121_/S sky130_fd_sc_hd__buf_4
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13774_ _17010_/A vssd1 vssd1 vccd1 vccd1 _13774_/X sky130_fd_sc_hd__buf_2
XFILLER_90_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18301_ _18301_/A vssd1 vssd1 vccd1 vccd1 _19985_/D sky130_fd_sc_hd__clkbuf_1
X_15513_ _15419_/X _15137_/X _15512_/X _15428_/X vssd1 vssd1 vccd1 vccd1 _15513_/X
+ sky130_fd_sc_hd__o211a_1
X_19281_ _20002_/CLK _19281_/D vssd1 vssd1 vccd1 vccd1 _19281_/Q sky130_fd_sc_hd__dfxtp_1
X_12725_ _12750_/B _12750_/C vssd1 vssd1 vccd1 vccd1 _12725_/X sky130_fd_sc_hd__or2_1
XANTENNA__17573__A0 _17112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15179__A2 _15177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16493_ _19231_/Q _13781_/X _16497_/S vssd1 vssd1 vccd1 vccd1 _16494_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12917__A _15735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18232_ _18278_/S vssd1 vssd1 vccd1 vccd1 _18241_/S sky130_fd_sc_hd__buf_4
XFILLER_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09498__A _14782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15444_ _15444_/A vssd1 vssd1 vccd1 vccd1 _15522_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12656_ _18542_/Q _12553_/X _12651_/X _12655_/X vssd1 vssd1 vccd1 vccd1 _12656_/X
+ sky130_fd_sc_hd__o22a_2
XANTENNA__12636__B _15474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12937__A1 _12874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18163_ _17672_/X _19924_/Q _18169_/S vssd1 vssd1 vccd1 vccd1 _18164_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12937__B2 _12906_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ _11607_/A _11607_/B vssd1 vssd1 vccd1 vccd1 _11608_/C sky130_fd_sc_hd__nor2_1
XFILLER_90_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10099__S1 _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12587_ _12587_/A vssd1 vssd1 vccd1 vccd1 _12657_/A sky130_fd_sc_hd__clkbuf_2
X_15375_ _15399_/A _15375_/B _15375_/C vssd1 vssd1 vccd1 vccd1 _15375_/X sky130_fd_sc_hd__and3_1
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17114_ _17114_/A vssd1 vssd1 vccd1 vccd1 _19494_/D sky130_fd_sc_hd__clkbuf_1
X_14326_ _14356_/A _14326_/B _14336_/D vssd1 vssd1 vccd1 vccd1 _18673_/D sky130_fd_sc_hd__nor3_1
XFILLER_8_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11538_ _11538_/A _11538_/B vssd1 vssd1 vccd1 vccd1 _11538_/Y sky130_fd_sc_hd__nor2_1
X_18094_ _18852_/Q _13661_/X _18101_/S vssd1 vssd1 vccd1 vccd1 _18094_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15947__B _15966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17045_ _17045_/A vssd1 vssd1 vccd1 vccd1 _19468_/D sky130_fd_sc_hd__clkbuf_1
X_11469_ _09664_/A _11468_/X _10886_/A vssd1 vssd1 vccd1 vccd1 _11469_/X sky130_fd_sc_hd__a21o_1
X_14257_ _14315_/A _14257_/B _14264_/D vssd1 vssd1 vccd1 vccd1 _18653_/D sky130_fd_sc_hd__nor3_1
XANTENNA__16124__A _16135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13362__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13208_ _13207_/A _13224_/C _12957_/A vssd1 vssd1 vccd1 vccd1 _13208_/X sky130_fd_sc_hd__o21a_1
X_14188_ _18635_/Q _18634_/Q _14188_/C vssd1 vssd1 vccd1 vccd1 _14190_/B sky130_fd_sc_hd__and3_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17654__S _17666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13139_ _13137_/X _18434_/Q _13203_/S vssd1 vssd1 vccd1 vccd1 _13140_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ _19488_/CLK _18996_/D vssd1 vssd1 vccd1 vccd1 _18996_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_140_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09961__A _18861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17947_ _17947_/A vssd1 vssd1 vccd1 vccd1 _19843_/D sky130_fd_sc_hd__clkbuf_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14579__A _14665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17878_ _19813_/Q _17090_/X _17880_/S vssd1 vssd1 vccd1 vccd1 _17879_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19617_ _19942_/CLK _19617_/D vssd1 vssd1 vccd1 vccd1 _19617_/Q sky130_fd_sc_hd__dfxtp_1
X_16829_ _16829_/A vssd1 vssd1 vccd1 vccd1 _19380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11715__B _13227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19548_ _19966_/CLK _19548_/D vssd1 vssd1 vccd1 vccd1 _19548_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12625__A0 _12621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09301_ _18978_/Q _18938_/Q vssd1 vssd1 vccd1 vccd1 _09301_/X sky130_fd_sc_hd__and2_1
XFILLER_81_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11979__A2 _14865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19479_ _19873_/CLK _19479_/D vssd1 vssd1 vccd1 vccd1 _19479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09232_ _11939_/C vssd1 vssd1 vccd1 vccd1 _14758_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11731__A _13656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13050__B1 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15327__C1 _15275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13658__A _14552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13889__C1 _13885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14550__B1 _14507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11364__B1 _11452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10082__A _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09996_ _19153_/Q _19414_/Q _19313_/Q _19648_/Q _10356_/S _09636_/A vssd1 vssd1 vccd1
+ vccd1 _09997_/B sky130_fd_sc_hd__mux4_1
XFILLER_131_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09871__A _19526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10014__S1 _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14605__A1 _13612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16908__S _16914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15802__B1 _15798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10840_ _18844_/Q vssd1 vssd1 vccd1 vccd1 _10840_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10771_ _11481_/A _10768_/X _10770_/X _09685_/A vssd1 vssd1 vccd1 vccd1 _10771_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ _12501_/B _12415_/X _12506_/Y _12509_/X vssd1 vssd1 vccd1 vccd1 _12510_/X
+ sky130_fd_sc_hd__o22a_4
X_13490_ _19063_/Q _12878_/X _13488_/X _13489_/X vssd1 vssd1 vccd1 vccd1 _13490_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_157_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12441_ _12389_/A _12389_/B _12438_/Y _12440_/X vssd1 vssd1 vccd1 vccd1 _12442_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12372_ _18467_/Q _12372_/B vssd1 vssd1 vccd1 vccd1 _12372_/X sky130_fd_sc_hd__or2_1
X_15160_ _15160_/A _15160_/B vssd1 vssd1 vccd1 vccd1 _15160_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11323_ _19322_/Q _19593_/Q _19817_/Q _19561_/Q _09586_/A _11322_/X vssd1 vssd1 vccd1
+ vccd1 _11323_/X sky130_fd_sc_hd__mux4_1
X_14111_ _13924_/B _14108_/B _14110_/Y vssd1 vssd1 vccd1 vccd1 _18613_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10691__S _10691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15091_ _11994_/A _15482_/B _15457_/A vssd1 vssd1 vccd1 vccd1 _15091_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14042_ _14042_/A _18590_/Q _14042_/C vssd1 vssd1 vccd1 vccd1 _14044_/B sky130_fd_sc_hd__and3_1
X_11254_ _11287_/A _11253_/X _09559_/A vssd1 vssd1 vccd1 vccd1 _11254_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09643__S0 _09598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _10208_/A vssd1 vssd1 vccd1 vccd1 _10469_/S sky130_fd_sc_hd__buf_4
XFILLER_134_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18850_ _18851_/CLK _18850_/D vssd1 vssd1 vccd1 vccd1 _18850_/Q sky130_fd_sc_hd__dfxtp_4
X_11185_ _11225_/A _11185_/B vssd1 vssd1 vccd1 vccd1 _11185_/Y sky130_fd_sc_hd__nor2_1
X_17801_ _17801_/A vssd1 vssd1 vccd1 vccd1 _19778_/D sky130_fd_sc_hd__clkbuf_1
X_10136_ _10112_/A _10133_/X _10135_/X _10192_/A vssd1 vssd1 vccd1 vccd1 _10137_/C
+ sky130_fd_sc_hd__o211a_1
X_18781_ _18819_/CLK _18781_/D vssd1 vssd1 vccd1 vccd1 _18781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15993_ _15993_/A vssd1 vssd1 vccd1 vccd1 _19027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17732_ _17732_/A vssd1 vssd1 vccd1 vccd1 _17732_/X sky130_fd_sc_hd__clkbuf_2
X_10067_ _09690_/A _10061_/X _10063_/Y _10066_/Y _09876_/X vssd1 vssd1 vccd1 vccd1
+ _10067_/X sky130_fd_sc_hd__o221a_1
X_14944_ _12715_/A _15160_/B _14956_/S vssd1 vssd1 vccd1 vccd1 _14944_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_189_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17663_ _17662_/X _19727_/Q _17666_/S vssd1 vssd1 vccd1 vccd1 _17664_/A sky130_fd_sc_hd__mux2_1
X_14875_ _14931_/A vssd1 vssd1 vccd1 vccd1 _15117_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19402_ _19636_/CLK _19402_/D vssd1 vssd1 vccd1 vccd1 _19402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16614_ _16614_/A vssd1 vssd1 vccd1 vccd1 _19285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13826_ _17062_/A vssd1 vssd1 vccd1 vccd1 _13826_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17594_ _17594_/A vssd1 vssd1 vccd1 vccd1 _19700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19333_ _19829_/CLK _19333_/D vssd1 vssd1 vccd1 vccd1 _19333_/Q sky130_fd_sc_hd__dfxtp_1
X_16545_ _19255_/Q _13857_/X _16545_/S vssd1 vssd1 vccd1 vccd1 _16546_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12083__A1 _12082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13750__B _13750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13757_ _17738_/A _18208_/A vssd1 vssd1 vccd1 vccd1 _13839_/A sky130_fd_sc_hd__nor2_4
X_10969_ _12239_/A _12835_/B vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__or2_1
XANTENNA__12647__A _18542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19264_ _19824_/CLK _19264_/D vssd1 vssd1 vccd1 vccd1 _19264_/Q sky130_fd_sc_hd__dfxtp_1
X_12708_ _15509_/A _12708_/B vssd1 vssd1 vccd1 vccd1 _12713_/A sky130_fd_sc_hd__xnor2_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16476_ _16532_/A vssd1 vssd1 vccd1 vccd1 _16545_/S sky130_fd_sc_hd__buf_8
X_13688_ _13688_/A _13693_/C vssd1 vssd1 vccd1 vccd1 _13688_/Y sky130_fd_sc_hd__xnor2_2
X_18215_ _19947_/Q _17643_/A _18219_/S vssd1 vssd1 vccd1 vccd1 _18216_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15958__A _15966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15427_ _15071_/X _15281_/X _15426_/X vssd1 vssd1 vccd1 vccd1 _15427_/X sky130_fd_sc_hd__a21o_1
X_19195_ _19948_/CLK _19195_/D vssd1 vssd1 vccd1 vccd1 _19195_/Q sky130_fd_sc_hd__dfxtp_1
X_12639_ _12639_/A _14907_/A vssd1 vssd1 vccd1 vccd1 _12640_/B sky130_fd_sc_hd__or2_1
XFILLER_129_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13583__A1 _13582_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18146_ _18146_/A vssd1 vssd1 vccd1 vccd1 _19916_/D sky130_fd_sc_hd__clkbuf_1
X_15358_ _15282_/X _15349_/X _15357_/X _15324_/X vssd1 vssd1 vccd1 vccd1 _15358_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14309_ _18669_/Q vssd1 vssd1 vccd1 vccd1 _14316_/B sky130_fd_sc_hd__clkbuf_1
X_18077_ _18847_/Q _13621_/X _18084_/S vssd1 vssd1 vccd1 vccd1 _18077_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12382__A _15338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15289_ _15286_/X _15291_/B _15287_/X _15288_/X vssd1 vssd1 vccd1 vccd1 _15289_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17028_ _19463_/Q _17026_/X _17040_/S vssd1 vssd1 vccd1 vccd1 _17029_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13197__B _18847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11346__B1 _11181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09850_ _19381_/Q _19716_/Q _09855_/A vssd1 vssd1 vccd1 vccd1 _09851_/B sky130_fd_sc_hd__mux2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09781_ _09891_/A _09769_/X _09837_/A vssd1 vssd1 vccd1 vccd1 _09781_/X sky130_fd_sc_hd__o21a_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _19526_/CLK _18979_/D vssd1 vssd1 vccd1 vccd1 _18979_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11726__A _14159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14102__A _14102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16728__S _16736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15260__A1 _12246_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13271__B1 _12881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12557__A _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_12_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09215_ _18832_/Q _18831_/Q vssd1 vssd1 vccd1 vccd1 _09215_/X sky130_fd_sc_hd__or2_1
XFILLER_50_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13574__A1 _13573_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11585__B1 _12856_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11432__S0 _11154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09979_ _20034_/Q _19872_/Q _19281_/Q _19051_/Q _09657_/A _09637_/A vssd1 vssd1 vccd1
+ vccd1 _09979_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_190_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _18586_/Q vssd1 vssd1 vccd1 vccd1 _14034_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_162_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _11941_/A _11941_/B _11983_/S _18981_/Q vssd1 vssd1 vccd1 vccd1 _12536_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17776__A0 _17688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _14663_/A _14660_/B vssd1 vssd1 vccd1 vccd1 _14661_/A sky130_fd_sc_hd__and2_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11872_ _18477_/Q _12982_/A _14555_/B _18780_/Q _11871_/X vssd1 vssd1 vccd1 vccd1
+ _11872_/X sky130_fd_sc_hd__a221o_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _13709_/A _19007_/Q vssd1 vssd1 vccd1 vccd1 _13611_/Y sky130_fd_sc_hd__nand2_1
X_10823_ _19666_/Q _19432_/Q _18497_/Q _19762_/Q _10872_/S _10664_/A vssd1 vssd1 vccd1
+ vccd1 _10824_/B sky130_fd_sc_hd__mux4_1
XFILLER_26_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13570__B _13570_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11499__S0 _11488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14591_ _18766_/Q _13579_/X _14598_/S vssd1 vssd1 vccd1 vccd1 _14592_/B sky130_fd_sc_hd__mux2_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13062__S _13350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16330_ _16329_/X _19169_/Q _16330_/S vssd1 vssd1 vccd1 vccd1 _16331_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13542_ _18999_/Q _13542_/B vssd1 vssd1 vccd1 vccd1 _13542_/X sky130_fd_sc_hd__or2_1
X_10754_ _19334_/Q _19605_/Q _19829_/Q _19573_/Q _10750_/S _10626_/A vssd1 vssd1 vccd1
+ vccd1 _10754_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10171__S0 _10208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13014__A0 _18838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16261_ _13219_/X _19143_/Q _16269_/S vssd1 vssd1 vccd1 vccd1 _16262_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10685_ _18439_/Q _19468_/Q _19505_/Q _19079_/Q _10637_/S _10010_/A vssd1 vssd1 vccd1
+ vccd1 _10685_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15554__A2 _12807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13473_ _13473_/A _18863_/Q vssd1 vssd1 vccd1 vccd1 _13473_/X sky130_fd_sc_hd__or2_1
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18000_ _18011_/A vssd1 vssd1 vccd1 vccd1 _18009_/S sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_172_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18548_/CLK sky130_fd_sc_hd__clkbuf_16
X_15212_ _15369_/A vssd1 vssd1 vccd1 vccd1 _15212_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09776__A _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ _18772_/Q _18771_/Q _12424_/C vssd1 vssd1 vccd1 vccd1 _12483_/C sky130_fd_sc_hd__and3_2
X_16192_ _16192_/A vssd1 vssd1 vccd1 vccd1 _19113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15143_ _14858_/X _15138_/B _15489_/A _15141_/X _15142_/Y vssd1 vssd1 vccd1 vccd1
+ _15143_/X sky130_fd_sc_hd__o2111a_1
X_12355_ _12406_/C vssd1 vssd1 vccd1 vccd1 _15321_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10715__A _10836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13317__A1 _13068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11306_ _11340_/A _11305_/X _11181_/X vssd1 vssd1 vccd1 vccd1 _11306_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15711__C1 _14540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12286_ _12280_/X _12281_/Y _12284_/X _13900_/A vssd1 vssd1 vccd1 vccd1 _12287_/B
+ sky130_fd_sc_hd__o211ai_2
X_15074_ _15097_/A vssd1 vssd1 vccd1 vccd1 _15074_/X sky130_fd_sc_hd__clkbuf_2
X_19951_ _19951_/CLK _19951_/D vssd1 vssd1 vccd1 vccd1 _19951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_187_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19526_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18902_ _19488_/CLK _18902_/D vssd1 vssd1 vccd1 vccd1 _18902_/Q sky130_fd_sc_hd__dfxtp_1
X_14025_ _14026_/A _14026_/B _14024_/Y vssd1 vssd1 vccd1 vccd1 _18583_/D sky130_fd_sc_hd__o21a_1
X_11237_ _11237_/A _11237_/B vssd1 vssd1 vccd1 vccd1 _11237_/X sky130_fd_sc_hd__and2_1
XFILLER_141_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19882_ _19882_/CLK _19882_/D vssd1 vssd1 vccd1 vccd1 _19882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18833_ _18972_/CLK _18833_/D vssd1 vssd1 vccd1 vccd1 _18833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11168_ _09881_/A _11152_/X _11166_/Y _09911_/A _11167_/Y vssd1 vssd1 vccd1 vccd1
+ _12830_/B sky130_fd_sc_hd__o32a_4
XFILLER_96_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10119_ _10305_/A _10118_/X _09565_/A vssd1 vssd1 vccd1 vccd1 _10119_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_110_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _20033_/CLK sky130_fd_sc_hd__clkbuf_16
X_18764_ _19885_/CLK _18764_/D vssd1 vssd1 vccd1 vccd1 _18764_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11099_ _18431_/Q _19460_/Q _19497_/Q _19071_/Q _11186_/S _11022_/A vssd1 vssd1 vccd1
+ vccd1 _11099_/X sky130_fd_sc_hd__mux4_1
X_15976_ _15978_/A _15978_/B _15976_/C vssd1 vssd1 vccd1 vccd1 _15976_/X sky130_fd_sc_hd__and3_1
XFILLER_49_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17715_ _17715_/A vssd1 vssd1 vccd1 vccd1 _19743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15960__B _15960_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14927_ _14927_/A vssd1 vssd1 vccd1 vccd1 _14937_/S sky130_fd_sc_hd__clkbuf_2
X_18695_ _19882_/CLK _18695_/D vssd1 vssd1 vccd1 vccd1 _18695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14857__A _15183_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17646_ _17646_/A vssd1 vssd1 vccd1 vccd1 _17646_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14858_ _15068_/A vssd1 vssd1 vccd1 vccd1 _14858_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15242__A1 _18841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_125_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _18924_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13809_ _13809_/A vssd1 vssd1 vccd1 vccd1 _18501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17577_ _17577_/A vssd1 vssd1 vccd1 vccd1 _19692_/D sky130_fd_sc_hd__clkbuf_1
X_14789_ _14789_/A _14789_/B vssd1 vssd1 vccd1 vccd1 _14789_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19316_ _19973_/CLK _19316_/D vssd1 vssd1 vccd1 vccd1 _19316_/Q sky130_fd_sc_hd__dfxtp_1
X_16528_ _19247_/Q _13832_/X _16530_/S vssd1 vssd1 vccd1 vccd1 _16529_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19247_ _20032_/CLK _19247_/D vssd1 vssd1 vccd1 vccd1 _19247_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17379__S _17387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16459_ _16459_/A vssd1 vssd1 vccd1 vccd1 _16468_/S sky130_fd_sc_hd__buf_4
XANTENNA__16283__S _16291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14592__A _14595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09686__A _09686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19178_ _20027_/CLK _19178_/D vssd1 vssd1 vccd1 vccd1 _19178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18129_ _18129_/A vssd1 vssd1 vccd1 vccd1 _19910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10625__A _10625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12616__A_N _12641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13001__A _17007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09902_ _09942_/A vssd1 vssd1 vccd1 vccd1 _11558_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15627__S _15901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18003__S _18009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12840__A _12840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20022_ _20022_/CLK _20022_/D vssd1 vssd1 vccd1 vccd1 _20022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09833_ _10210_/A vssd1 vssd1 vccd1 vccd1 _09833_/X sky130_fd_sc_hd__buf_4
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _10292_/A vssd1 vssd1 vccd1 vccd1 _09765_/A sky130_fd_sc_hd__clkbuf_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09695_ _18984_/Q _18939_/Q vssd1 vssd1 vccd1 vccd1 _09696_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__13492__B1 _11733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13244__B1 _12897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17289__S _17293_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_137_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09596__A _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ _19243_/Q _19738_/Q _10470_/S vssd1 vssd1 vccd1 vccd1 _10470_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14749__D_N _09454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ _12140_/A vssd1 vssd1 vccd1 vccd1 _12140_/X sky130_fd_sc_hd__buf_4
XFILLER_151_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12071_ _18759_/Q _12071_/B _12071_/C vssd1 vssd1 vccd1 vccd1 _12071_/X sky130_fd_sc_hd__and3_1
XFILLER_104_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11022_ _11022_/A vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__buf_2
XFILLER_150_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15830_ hold4/A _15816_/X _15820_/X input36/X vssd1 vssd1 vccd1 vccd1 _15831_/B sky130_fd_sc_hd__a22o_1
XANTENNA__17752__S _17760_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _14749_/B _15752_/X _15760_/X _15756_/X vssd1 vssd1 vccd1 vccd1 _18950_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12973_ _18867_/Q _12973_/B vssd1 vssd1 vccd1 vccd1 _13015_/C sky130_fd_sc_hd__and2_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19989_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _19656_/Q vssd1 vssd1 vccd1 vccd1 _17501_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__18149__A _18206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _18807_/Q _11748_/X _14716_/S vssd1 vssd1 vccd1 vccd1 _14713_/A sky130_fd_sc_hd__mux2_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _18977_/Q vssd1 vssd1 vccd1 vccd1 _15847_/A sky130_fd_sc_hd__buf_4
XFILLER_73_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18480_ _18544_/CLK _18480_/D vssd1 vssd1 vccd1 vccd1 _18480_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _15692_/A vssd1 vssd1 vccd1 vccd1 _18922_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15224__A1 _12186_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _17103_/X _19624_/Q _17437_/S vssd1 vssd1 vccd1 vccd1 _17432_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _14646_/A _14643_/B vssd1 vssd1 vccd1 vccd1 _14644_/A sky130_fd_sc_hd__and2_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11855_ _18726_/Q _11855_/B vssd1 vssd1 vccd1 vccd1 _11855_/X sky130_fd_sc_hd__and2_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output105_A _14811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12197__A _18461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10806_ _19236_/Q _19731_/Q _11486_/S vssd1 vssd1 vccd1 vccd1 _10806_/X sky130_fd_sc_hd__mux2_1
X_17362_ _17362_/A vssd1 vssd1 vccd1 vccd1 _19593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18174__A0 _17688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19641_/CLK sky130_fd_sc_hd__clkbuf_16
X_14574_ _14577_/A _14574_/B vssd1 vssd1 vccd1 vccd1 _14575_/A sky130_fd_sc_hd__and2_1
X_11786_ _19884_/Q _12946_/A _11703_/A _18457_/Q vssd1 vssd1 vccd1 vccd1 _11786_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11797__B1 _11796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19101_ _19982_/CLK _19101_/D vssd1 vssd1 vccd1 vccd1 _19101_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17199__S _17199_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16313_ _17649_/A vssd1 vssd1 vccd1 vccd1 _16313_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13525_ _13535_/B _13524_/Y _12344_/X vssd1 vssd1 vccd1 vccd1 _13526_/B sky130_fd_sc_hd__a21o_1
X_10737_ _15943_/B vssd1 vssd1 vccd1 vccd1 _10760_/A sky130_fd_sc_hd__inv_2
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17293_ _17112_/X _19563_/Q _17293_/S vssd1 vssd1 vccd1 vccd1 _17294_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19032_ _19853_/CLK _19032_/D vssd1 vssd1 vccd1 vccd1 _19032_/Q sky130_fd_sc_hd__dfxtp_1
X_16244_ _16244_/A vssd1 vssd1 vccd1 vccd1 _19135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13456_ _18611_/Q _13120_/A _13082_/X _18743_/Q vssd1 vssd1 vccd1 vccd1 _13456_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10668_ _10668_/A _10668_/B _10668_/C vssd1 vssd1 vccd1 vccd1 _10668_/X sky130_fd_sc_hd__or3_2
XANTENNA__11549__B1 _09568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ _12459_/A _12433_/B vssd1 vssd1 vccd1 vccd1 _12408_/B sky130_fd_sc_hd__nand2_2
XFILLER_154_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16175_ _16221_/S vssd1 vssd1 vccd1 vccd1 _16184_/S sky130_fd_sc_hd__buf_2
X_10599_ _10832_/A _10599_/B vssd1 vssd1 vccd1 vccd1 _10599_/Y sky130_fd_sc_hd__nor2_1
X_13387_ _13385_/X _18449_/Q _13464_/S vssd1 vssd1 vccd1 vccd1 _13388_/A sky130_fd_sc_hd__mux2_1
Xoutput107 _12866_/B vssd1 vssd1 vccd1 vccd1 io_dbus_st_type[0] sky130_fd_sc_hd__buf_2
XFILLER_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput118 _12849_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[18] sky130_fd_sc_hd__buf_2
X_15126_ _15093_/X _15109_/X _15125_/X _15048_/X _12046_/Y vssd1 vssd1 vccd1 vccd1
+ _15126_/X sky130_fd_sc_hd__a32o_1
XFILLER_115_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12338_ _12338_/A vssd1 vssd1 vccd1 vccd1 _12338_/X sky130_fd_sc_hd__buf_2
Xoutput129 _12862_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[28] sky130_fd_sc_hd__buf_2
XFILLER_141_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19934_ _19998_/CLK _19934_/D vssd1 vssd1 vccd1 vccd1 _19934_/Q sky130_fd_sc_hd__dfxtp_1
X_15057_ _14938_/X _14926_/X _15114_/S vssd1 vssd1 vccd1 vccd1 _15057_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12269_ _12299_/A _12298_/A vssd1 vssd1 vccd1 vccd1 _12272_/A sky130_fd_sc_hd__xor2_4
X_14008_ _14044_/A _14008_/B _14013_/C vssd1 vssd1 vccd1 vccd1 _18577_/D sky130_fd_sc_hd__nor3_1
X_19865_ _19865_/CLK _19865_/D vssd1 vssd1 vccd1 vccd1 _19865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18816_ _19910_/CLK _18816_/D vssd1 vssd1 vccd1 vccd1 _18816_/Q sky130_fd_sc_hd__dfxtp_1
X_19796_ _19796_/CLK _19796_/D vssd1 vssd1 vccd1 vccd1 _19796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15959_ _19013_/Q _15951_/X _15958_/X vssd1 vssd1 vccd1 vccd1 _19013_/D sky130_fd_sc_hd__a21o_1
X_18747_ _19063_/CLK _18747_/D vssd1 vssd1 vccd1 vccd1 _18747_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16278__S _16280_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10288__B1 _09807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09480_ _09480_/A _11951_/A _14756_/B vssd1 vssd1 vccd1 vccd1 _09496_/A sky130_fd_sc_hd__nor3_1
X_18678_ _18687_/CLK _18678_/D vssd1 vssd1 vccd1 vccd1 _18678_/Q sky130_fd_sc_hd__dfxtp_1
X_17629_ _17629_/A vssd1 vssd1 vccd1 vccd1 _19716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15910__S _15946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17837__S _17843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16741__S _16747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15865__B _16839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17138__A _17675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16977__A _16977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20005_ _20005_/CLK _20005_/D vssd1 vssd1 vccd1 vccd1 _20005_/Q sky130_fd_sc_hd__dfxtp_1
X_09816_ _09816_/A vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_63_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ _09747_/A vssd1 vssd1 vccd1 vccd1 _09940_/A sky130_fd_sc_hd__buf_2
XFILLER_36_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09678_ _19158_/Q _19419_/Q _19318_/Q _19653_/Q _09920_/S _10057_/A vssd1 vssd1 vccd1
+ vccd1 _09679_/B sky130_fd_sc_hd__mux4_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10374__S0 _10279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16916__S _16918_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11125__S _11125_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A _11640_/B vssd1 vssd1 vccd1 vccd1 _11642_/A sky130_fd_sc_hd__or2_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10249__B _12856_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ _19159_/Q _19420_/Q _19319_/Q _19654_/Q _11566_/S _11554_/A vssd1 vssd1 vccd1
+ vccd1 _11572_/B sky130_fd_sc_hd__mux4_1
XANTENNA__16706__A1 _13774_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13310_ _19902_/Q _13451_/B vssd1 vssd1 vccd1 vccd1 _13310_/X sky130_fd_sc_hd__and2_1
X_10522_ _10522_/A vssd1 vssd1 vccd1 vccd1 _10522_/X sky130_fd_sc_hd__buf_2
XFILLER_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12991__A2 _11682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14290_ _18663_/Q _18662_/Q _18661_/Q _14290_/D vssd1 vssd1 vccd1 vccd1 _14300_/D
+ sky130_fd_sc_hd__and4_1
X_10453_ _10458_/A _10453_/B vssd1 vssd1 vccd1 vccd1 _10453_/X sky130_fd_sc_hd__or2_1
X_13241_ input9/X _13231_/X _13234_/X vssd1 vssd1 vccd1 vccd1 _13248_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__17747__S _17749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09476__D _14766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input66_A io_ibus_valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ _10375_/X _10378_/X _10380_/X _10383_/X _09807_/A vssd1 vssd1 vccd1 vccd1
+ _10384_/X sky130_fd_sc_hd__a221o_4
X_13172_ _18846_/Q _13609_/B _13349_/S vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ _12215_/A _12215_/B _12092_/A vssd1 vssd1 vccd1 vccd1 _12124_/B sky130_fd_sc_hd__a21o_2
X_17980_ _17980_/A vssd1 vssd1 vccd1 vccd1 _19857_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12480__A _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12054_ _15633_/C _12153_/B _12153_/C _12054_/D vssd1 vssd1 vccd1 vccd1 _12054_/X
+ sky130_fd_sc_hd__and4_1
X_16931_ _16313_/X _19425_/Q _16931_/S vssd1 vssd1 vccd1 vccd1 _16932_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11005_ _19200_/Q _19791_/Q _19953_/Q _19168_/Q _11048_/S _10978_/A vssd1 vssd1 vccd1
+ vccd1 _11006_/B sky130_fd_sc_hd__mux4_1
XANTENNA__15791__A _15833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19650_ _19972_/CLK _19650_/D vssd1 vssd1 vccd1 vccd1 _19650_/Q sky130_fd_sc_hd__dfxtp_1
X_16862_ _16316_/X _19394_/Q _16870_/S vssd1 vssd1 vccd1 vccd1 _16863_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14248__A2 _14279_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18601_ _19941_/CLK _18601_/D vssd1 vssd1 vccd1 vccd1 _18601_/Q sky130_fd_sc_hd__dfxtp_1
X_15813_ _15813_/A _15813_/B vssd1 vssd1 vccd1 vccd1 _15814_/A sky130_fd_sc_hd__and2_1
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19581_ _19581_/CLK _19581_/D vssd1 vssd1 vccd1 vccd1 _19581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16793_ _16339_/X _19364_/Q _16797_/S vssd1 vssd1 vccd1 vccd1 _16794_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16098__S _16100_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13456__B1 _13082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18532_ _18868_/CLK _18532_/D vssd1 vssd1 vccd1 vccd1 _18532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15744_ _09522_/A _15734_/X _15742_/X _15743_/X vssd1 vssd1 vccd1 vccd1 _18943_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12956_ _12956_/A _12956_/B vssd1 vssd1 vccd1 vccd1 _12956_/Y sky130_fd_sc_hd__nor2_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12639__B _14907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11543__B _11543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18463_ _18526_/CLK _18463_/D vssd1 vssd1 vccd1 vccd1 _18463_/Q sky130_fd_sc_hd__dfxtp_1
X_11907_ _09305_/X _11905_/X _09342_/X _12317_/A _12536_/A vssd1 vssd1 vccd1 vccd1
+ _14771_/A sky130_fd_sc_hd__o2111a_4
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _18915_/Q _12501_/B _15677_/S vssd1 vssd1 vccd1 vccd1 _15676_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16826__S _16830_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12887_ _12887_/A vssd1 vssd1 vccd1 vccd1 _12887_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _19617_/Q _17078_/X _17420_/S vssd1 vssd1 vccd1 vccd1 _17415_/A sky130_fd_sc_hd__mux2_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14956__A0 _12738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14629_/A _14626_/B vssd1 vssd1 vccd1 vccd1 _14627_/A sky130_fd_sc_hd__and2_1
XFILLER_159_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18394_ _17694_/X _20027_/Q _18396_/S vssd1 vssd1 vccd1 vccd1 _18395_/A sky130_fd_sc_hd__mux2_1
X_11838_ _13879_/A _18712_/Q _14534_/S vssd1 vssd1 vccd1 vccd1 _11838_/X sky130_fd_sc_hd__or3_1
XFILLER_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17345_ _17345_/A vssd1 vssd1 vccd1 vccd1 _19586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _18757_/Q _14554_/X _14601_/A vssd1 vssd1 vccd1 vccd1 _14558_/B sky130_fd_sc_hd__mux2_1
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11769_ _18746_/Q _13926_/A vssd1 vssd1 vccd1 vccd1 _11774_/A sky130_fd_sc_hd__or2_1
XFILLER_147_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10442__B1 _09913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13508_ _13508_/A _13508_/B vssd1 vssd1 vccd1 vccd1 _16069_/B sky130_fd_sc_hd__nand2_2
XFILLER_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17276_ _17192_/X _19556_/Q _17276_/S vssd1 vssd1 vccd1 vccd1 _17277_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14488_ _14488_/A vssd1 vssd1 vccd1 vccd1 _14493_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_19015_ _19023_/CLK _19015_/D vssd1 vssd1 vccd1 vccd1 _19015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16227_ _16295_/S vssd1 vssd1 vccd1 vccd1 _16236_/S sky130_fd_sc_hd__buf_2
XANTENNA__17657__S _17666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13439_ _13439_/A _13725_/B vssd1 vssd1 vccd1 vccd1 _13439_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15966__A _15966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16561__S _16569_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09964__A _10493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16158_ _12963_/X _19098_/Q _16162_/S vssd1 vssd1 vccd1 vccd1 _16159_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15109_ _14977_/X _15098_/X _15108_/X _15005_/X vssd1 vssd1 vccd1 vccd1 _15109_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16089_ _13002_/X _19068_/Q _16089_/S vssd1 vssd1 vccd1 vccd1 _16090_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12390__A _12390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16881__A0 _16345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15684__A1 _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19917_ _19981_/CLK _19917_/D vssd1 vssd1 vccd1 vccd1 _19917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17392__S _17398_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19848_ _19946_/CLK _19848_/D vssd1 vssd1 vccd1 vccd1 _19848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11170__A1 _15925_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09601_ _10996_/A vssd1 vssd1 vccd1 vccd1 _11050_/A sky130_fd_sc_hd__buf_2
XFILLER_95_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19779_ _19973_/CLK _19779_/D vssd1 vssd1 vccd1 vccd1 _19779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11734__A _11734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ _09532_/A vssd1 vssd1 vccd1 vccd1 _09532_/X sky130_fd_sc_hd__buf_2
XFILLER_25_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09204__A _11956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09463_ _18992_/Q vssd1 vssd1 vccd1 vccd1 _12316_/A sky130_fd_sc_hd__buf_4
XANTENNA__16736__S _16736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15739__A2 _15738_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14947__A0 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09394_ _09394_/A _09401_/A vssd1 vssd1 vccd1 vccd1 _11703_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10659__S1 _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17567__S _17573_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09874__A _09874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09324__B_N _09468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10736__A1 _09546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10831__S1 _10820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15675__A1 _12501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ _15531_/A _12758_/B _15542_/A _14990_/A vssd1 vssd1 vccd1 vccd1 _12811_/B
+ sky130_fd_sc_hd__o31a_1
X_13790_ _17026_/A vssd1 vssd1 vccd1 vccd1 _13790_/X sky130_fd_sc_hd__buf_2
XFILLER_90_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12741_ _12741_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _12742_/B sky130_fd_sc_hd__nor2_2
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16646__S _16652_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10672__B1 _09563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15460_ _15506_/A _15463_/A vssd1 vssd1 vccd1 vccd1 _15460_/X sky130_fd_sc_hd__or2_1
XFILLER_31_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12672_ _18543_/Q vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__buf_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _18699_/Q _18698_/Q _14411_/C _14411_/D vssd1 vssd1 vccd1 vccd1 _14422_/D
+ sky130_fd_sc_hd__and4_1
X_11623_ _11595_/X _11596_/Y _11622_/X vssd1 vssd1 vccd1 vccd1 _11628_/B sky130_fd_sc_hd__o21ai_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15391_ _18850_/Q _15363_/X _15390_/X vssd1 vssd1 vccd1 vccd1 _18850_/D sky130_fd_sc_hd__o21a_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17130_ _17130_/A vssd1 vssd1 vccd1 vccd1 _19499_/D sky130_fd_sc_hd__clkbuf_1
X_14342_ _14345_/B _14364_/A _14332_/X vssd1 vssd1 vccd1 vccd1 _14342_/Y sky130_fd_sc_hd__a21oi_1
X_11554_ _11554_/A vssd1 vssd1 vccd1 vccd1 _11565_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17061_ _17061_/A vssd1 vssd1 vccd1 vccd1 _19473_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17477__S _17481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10505_ _18442_/Q _19471_/Q _19508_/Q _19082_/Q _09653_/A _10542_/A vssd1 vssd1 vccd1
+ vccd1 _10505_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14273_ _14288_/A _14273_/B vssd1 vssd1 vccd1 vccd1 _14273_/Y sky130_fd_sc_hd__nor2_1
X_11485_ _09848_/A _11475_/X _11484_/X _09538_/A _18846_/Q vssd1 vssd1 vccd1 vccd1
+ _15940_/C sky130_fd_sc_hd__a32o_4
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16012_ _13137_/X _19036_/Q _16020_/S vssd1 vssd1 vccd1 vccd1 _16013_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09784__A _10094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13224_ _18880_/Q _18881_/Q _13224_/C vssd1 vssd1 vccd1 vccd1 _13256_/C sky130_fd_sc_hd__and3_1
XFILLER_155_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10436_ _10484_/A _10435_/X _09779_/A vssd1 vssd1 vccd1 vccd1 _10436_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09342__C_N _09341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output172_A _12235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13155_ _18877_/Q vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__clkbuf_2
X_10367_ _10064_/A _10366_/X _09566_/A vssd1 vssd1 vccd1 vccd1 _10367_/X sky130_fd_sc_hd__o21a_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15666__A1 _12416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12106_ _16069_/A _12134_/B vssd1 vssd1 vccd1 vccd1 _12107_/B sky130_fd_sc_hd__or2b_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10298_ _10282_/X _10288_/X _10297_/X _09823_/A vssd1 vssd1 vccd1 vccd1 _10298_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17963_ _19850_/Q _17004_/X _17965_/S vssd1 vssd1 vccd1 vccd1 _17964_/A sky130_fd_sc_hd__mux2_1
X_13086_ _18873_/Q vssd1 vssd1 vccd1 vccd1 _13580_/A sky130_fd_sc_hd__buf_2
X_19702_ _19960_/CLK _19702_/D vssd1 vssd1 vccd1 vccd1 _19702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16914_ _16393_/X _19418_/Q _16914_/S vssd1 vssd1 vccd1 vccd1 _16915_/A sky130_fd_sc_hd__mux2_1
X_12037_ _12078_/D vssd1 vssd1 vccd1 vccd1 _15103_/B sky130_fd_sc_hd__buf_2
XANTENNA__15952__C _15952_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17894_ _17894_/A vssd1 vssd1 vccd1 vccd1 _19819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19633_ _19633_/CLK _19633_/D vssd1 vssd1 vccd1 vccd1 _19633_/Q sky130_fd_sc_hd__dfxtp_1
X_16845_ _16845_/A vssd1 vssd1 vccd1 vccd1 _19388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11554__A _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17940__S _17948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16776_ _16776_/A vssd1 vssd1 vccd1 vccd1 _19356_/D sky130_fd_sc_hd__clkbuf_1
X_19564_ _19951_/CLK _19564_/D vssd1 vssd1 vccd1 vccd1 _19564_/Q sky130_fd_sc_hd__dfxtp_1
X_13988_ _18570_/Q _13990_/C _13987_/Y vssd1 vssd1 vccd1 vccd1 _18570_/D sky130_fd_sc_hd__o21a_1
XFILLER_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18515_ _19842_/CLK _18515_/D vssd1 vssd1 vccd1 vccd1 _18515_/Q sky130_fd_sc_hd__dfxtp_1
X_15727_ hold2/X _15720_/X _15726_/Y _15713_/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__o211a_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _17640_/A vssd1 vssd1 vccd1 vccd1 _12939_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16556__S _16558_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19495_ _19982_/CLK _19495_/D vssd1 vssd1 vccd1 vccd1 _19495_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18337__A _18337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14865__A _14865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18446_ _19999_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_1
X_15658_ _18907_/Q _18528_/Q _15666_/S vssd1 vssd1 vccd1 vccd1 _15659_/A sky130_fd_sc_hd__mux2_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14609_ _14612_/A _14609_/B vssd1 vssd1 vccd1 vccd1 _14610_/A sky130_fd_sc_hd__and2_1
X_18377_ _17668_/X _20019_/Q _18385_/S vssd1 vssd1 vccd1 vccd1 _18378_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12404__A1 _09458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15589_ _13174_/A _18909_/Q _15589_/S vssd1 vssd1 vccd1 vccd1 _15590_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12385__A _12385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17328_ _17339_/A vssd1 vssd1 vccd1 vccd1 _17337_/S sky130_fd_sc_hd__buf_4
XFILLER_30_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_11_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__B1 _09279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__A1 _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17387__S _17387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17259_ _17167_/X _19548_/Q _17265_/S vssd1 vssd1 vccd1 vccd1 _17260_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16291__S _16291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12168__A0 _18763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11066__S1 _11065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11143__A1 _09848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16320__A _17656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11143__B2 _18839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11694__A2 _11683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17850__S _17854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09515_ _12004_/C _09513_/X _09514_/X vssd1 vssd1 vccd1 vccd1 _14765_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__16466__S _16468_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12994__S _13215_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _15856_/A _13518_/A vssd1 vssd1 vccd1 vccd1 _14771_/B sky130_fd_sc_hd__nor2_2
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13199__A2 _13091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ _15775_/A _18955_/Q _18954_/Q _18953_/Q vssd1 vssd1 vccd1 vccd1 _14227_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA__12295__A _15936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14714__S _14716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12159__B1 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15896__A1 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11270_ _19355_/Q _19690_/Q _11270_/S vssd1 vssd1 vccd1 vccd1 _11270_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10221_ _10392_/A _10207_/Y _10210_/Y _10220_/Y vssd1 vssd1 vccd1 vccd1 _10221_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _10208_/A vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13854__A _17090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10083_ _19937_/Q _19551_/Q _20001_/Q _19120_/Q _09939_/A _10278_/A vssd1 vssd1 vccd1
+ vccd1 _10084_/B sky130_fd_sc_hd__mux4_1
X_14960_ _15082_/B _14958_/X _15169_/A vssd1 vssd1 vccd1 vccd1 _14960_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10568__S0 _10529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13911_ _18549_/Q _12820_/A _12816_/X _12820_/Y _14792_/A vssd1 vssd1 vccd1 vccd1
+ _18549_/D sky130_fd_sc_hd__o221a_1
XFILLER_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input29_A io_dbus_rdata[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__S _10691_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ _14882_/X _14888_/X _15118_/S vssd1 vssd1 vccd1 vccd1 _14891_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17760__S _17760_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16630_ _16313_/X _19292_/Q _16630_/S vssd1 vssd1 vccd1 vccd1 _16631_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13842_ _17078_/A vssd1 vssd1 vccd1 vccd1 _13842_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16561_ _19261_/Q _13774_/X _16569_/S vssd1 vssd1 vccd1 vccd1 _16562_/A sky130_fd_sc_hd__mux2_1
X_13773_ _13773_/A vssd1 vssd1 vccd1 vccd1 _18490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14685__A _14742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ _11328_/A vssd1 vssd1 vccd1 vccd1 _11212_/A sky130_fd_sc_hd__buf_2
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18300_ _17662_/X _19985_/Q _18302_/S vssd1 vssd1 vccd1 vccd1 _18301_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15512_ _14977_/X _15135_/X _15511_/X _15400_/X vssd1 vssd1 vccd1 vccd1 _15512_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09779__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19280_ _20033_/CLK _19280_/D vssd1 vssd1 vccd1 vccd1 _19280_/Q sky130_fd_sc_hd__dfxtp_1
X_12724_ _18784_/Q vssd1 vssd1 vccd1 vccd1 _12750_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16492_ _16492_/A vssd1 vssd1 vccd1 vccd1 _19230_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10740__S0 _10750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12917__B _16474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18231_ _18231_/A vssd1 vssd1 vccd1 vccd1 _19954_/D sky130_fd_sc_hd__clkbuf_1
X_15443_ _15443_/A vssd1 vssd1 vccd1 vccd1 _18854_/D sky130_fd_sc_hd__clkbuf_1
X_12655_ _12347_/X _12653_/Y _12654_/X _12350_/X vssd1 vssd1 vccd1 vccd1 _12655_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18162_ _18162_/A vssd1 vssd1 vccd1 vccd1 _19923_/D sky130_fd_sc_hd__clkbuf_1
X_11606_ _11606_/A _11606_/B _11606_/C vssd1 vssd1 vccd1 vccd1 _11606_/Y sky130_fd_sc_hd__nand3_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15374_ _15305_/X _15367_/Y _15373_/Y vssd1 vssd1 vccd1 vccd1 _15375_/C sky130_fd_sc_hd__a21oi_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12586_ _12513_/A _12515_/B _12540_/A _15436_/A _12515_/A vssd1 vssd1 vccd1 vccd1
+ _12591_/A sky130_fd_sc_hd__o41a_1
X_17113_ _17112_/X _19494_/Q _17113_/S vssd1 vssd1 vccd1 vccd1 _17114_/A sky130_fd_sc_hd__mux2_1
X_14325_ _18673_/Q _18672_/Q _18671_/Q _14325_/D vssd1 vssd1 vccd1 vccd1 _14336_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_117_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11537_ _19159_/Q _19420_/Q _19319_/Q _19654_/Q _09635_/X _09639_/X vssd1 vssd1 vccd1
+ vccd1 _11538_/B sky130_fd_sc_hd__mux4_2
XFILLER_8_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18093_ _18093_/A vssd1 vssd1 vccd1 vccd1 _19899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15947__C _15947_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15887__A1 _09471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17044_ _19468_/Q _17042_/X _17056_/S vssd1 vssd1 vccd1 vccd1 _17045_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15887__B2 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output97_A _12094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14256_ _18651_/Q _18650_/Q _14256_/C _14256_/D vssd1 vssd1 vccd1 vccd1 _14264_/D
+ sky130_fd_sc_hd__and4_2
XFILLER_172_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11468_ _19237_/Q _19732_/Q _11468_/S vssd1 vssd1 vccd1 vccd1 _11468_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17935__S _17937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ _13207_/A _13224_/C vssd1 vssd1 vccd1 vccd1 _13207_/Y sky130_fd_sc_hd__nand2_1
X_10419_ _18853_/Q vssd1 vssd1 vccd1 vccd1 _10419_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10453__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14187_ _18634_/Q _14188_/C _18635_/Q vssd1 vssd1 vccd1 vccd1 _14189_/B sky130_fd_sc_hd__a21oi_1
XFILLER_48_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11373__A1 _11206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _11440_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11399_/X sky130_fd_sc_hd__or2_1
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13138_ _13502_/S vssd1 vssd1 vccd1 vccd1 _13203_/S sky130_fd_sc_hd__buf_2
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _18997_/CLK _18995_/D vssd1 vssd1 vccd1 vccd1 _18995_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _19843_/Q _17084_/X _17948_/S vssd1 vssd1 vccd1 vccd1 _17947_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _18558_/Q vssd1 vssd1 vccd1 vccd1 _13956_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10333__C1 _10162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17877_ _17877_/A vssd1 vssd1 vccd1 vccd1 _19812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17670__S _17682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19616_ _20033_/CLK _19616_/D vssd1 vssd1 vccd1 vccd1 _19616_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10884__B1 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16828_ _16390_/X _19380_/Q _16830_/S vssd1 vssd1 vccd1 vccd1 _16829_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19547_ _19997_/CLK _19547_/D vssd1 vssd1 vccd1 vccd1 _19547_/Q sky130_fd_sc_hd__dfxtp_1
X_16759_ _16759_/A vssd1 vssd1 vccd1 vccd1 _19349_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14595__A _14595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09300_ _16846_/B _09465_/C _18976_/Q vssd1 vssd1 vccd1 vccd1 _09542_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__09689__A _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19478_ _20033_/CLK _19478_/D vssd1 vssd1 vccd1 vccd1 _19478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09231_ _09480_/A _11951_/A _09456_/A vssd1 vssd1 vccd1 vccd1 _11939_/C sky130_fd_sc_hd__or3_1
X_18429_ _19693_/CLK _18429_/D vssd1 vssd1 vccd1 vccd1 _18429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10939__A1 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12843__A _12843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11364__A1 _11292_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10798__S0 _10797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09995_ _09995_/A vssd1 vssd1 vccd1 vccd1 _10356_/S sky130_fd_sc_hd__buf_4
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13105__A2 _13081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10324__C1 _09876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17580__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10770_ _10936_/A _10770_/B vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__or2_1
XFILLER_71_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10722__S0 _10764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09429_ _15633_/A _12918_/B vssd1 vssd1 vccd1 vccd1 _15719_/A sky130_fd_sc_hd__nand2_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12440_ _12411_/A _14877_/A _12439_/X vssd1 vssd1 vccd1 vccd1 _12440_/X sky130_fd_sc_hd__o21a_1
XFILLER_139_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12371_ _12479_/S _12369_/X _12370_/X _12056_/X vssd1 vssd1 vccd1 vccd1 _12371_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12753__A _12753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14110_ _13924_/B _14108_/B _14102_/X vssd1 vssd1 vccd1 vccd1 _14110_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_125_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11322_ _11322_/A vssd1 vssd1 vccd1 vccd1 _11322_/X sky130_fd_sc_hd__buf_2
XFILLER_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15090_ _14830_/X _15069_/X _15088_/X _15089_/X vssd1 vssd1 vccd1 vccd1 _15090_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14541__A1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041_ _14042_/A _14042_/C _14040_/Y vssd1 vssd1 vccd1 vccd1 _18589_/D sky130_fd_sc_hd__o21a_1
X_11253_ _18429_/Q _19458_/Q _19495_/Q _19069_/Q _11212_/X _11045_/X vssd1 vssd1 vccd1
+ vccd1 _11253_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10789__S0 _10787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09643__S1 _09851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ _09849_/A _10194_/X _10203_/X _09540_/A _18859_/Q vssd1 vssd1 vccd1 vccd1
+ _15972_/C sky130_fd_sc_hd__a32o_4
X_11184_ _19659_/Q _19425_/Q _18490_/Q _19755_/Q _11171_/X _11172_/X vssd1 vssd1 vccd1
+ vccd1 _11185_/B sky130_fd_sc_hd__mux4_1
XFILLER_122_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17800_ _17723_/X _19778_/Q _17804_/S vssd1 vssd1 vccd1 vccd1 _17801_/A sky130_fd_sc_hd__mux2_1
X_10135_ _10553_/A _10135_/B vssd1 vssd1 vccd1 vccd1 _10135_/X sky130_fd_sc_hd__or2_1
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15992_ _12939_/X _19027_/Q _15998_/S vssd1 vssd1 vccd1 vccd1 _15993_/A sky130_fd_sc_hd__mux2_1
X_18780_ _19900_/CLK _18780_/D vssd1 vssd1 vccd1 vccd1 _18780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10066_ _10064_/X _10065_/X _09980_/X vssd1 vssd1 vccd1 vccd1 _10066_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17731_ _17731_/A vssd1 vssd1 vccd1 vccd1 _19748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14943_ _12713_/B _15138_/B _14956_/S vssd1 vssd1 vccd1 vccd1 _14943_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output135_A _12827_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17243__A0 _17144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17490__S _17492_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14874_ _14870_/X _14872_/X _15032_/S vssd1 vssd1 vccd1 vccd1 _14874_/X sky130_fd_sc_hd__mux2_1
X_17662_ _17662_/A vssd1 vssd1 vccd1 vccd1 _17662_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19401_ _19989_/CLK _19401_/D vssd1 vssd1 vccd1 vccd1 _19401_/Q sky130_fd_sc_hd__dfxtp_1
X_13825_ _13825_/A vssd1 vssd1 vccd1 vccd1 _18506_/D sky130_fd_sc_hd__clkbuf_1
X_16613_ _19285_/Q _13851_/X _16613_/S vssd1 vssd1 vccd1 vccd1 _16614_/A sky130_fd_sc_hd__mux2_1
X_17593_ _17141_/X _19700_/Q _17595_/S vssd1 vssd1 vccd1 vccd1 _17594_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19332_ _20025_/CLK _19332_/D vssd1 vssd1 vccd1 vccd1 _19332_/Q sky130_fd_sc_hd__dfxtp_1
X_16544_ _16544_/A vssd1 vssd1 vccd1 vccd1 _19254_/D sky130_fd_sc_hd__clkbuf_1
X_13756_ _18280_/A vssd1 vssd1 vccd1 vccd1 _18208_/A sky130_fd_sc_hd__buf_2
X_10968_ _12239_/A _12835_/B vssd1 vssd1 vccd1 vccd1 _11604_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13280__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _12756_/A _15498_/A _12686_/B vssd1 vssd1 vccd1 vccd1 _12708_/B sky130_fd_sc_hd__a21oi_1
XFILLER_149_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16475_ _16692_/A _17635_/A vssd1 vssd1 vccd1 vccd1 _16532_/A sky130_fd_sc_hd__nor2_4
X_19263_ _19949_/CLK _19263_/D vssd1 vssd1 vccd1 vccd1 _19263_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10448__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16834__S _16834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13687_ _18476_/Q _13517_/X _13682_/Y _13686_/X vssd1 vssd1 vccd1 vccd1 _18476_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10899_ _19202_/Q _19793_/Q _19955_/Q _19170_/Q _10892_/X _10893_/X vssd1 vssd1 vccd1
+ vccd1 _10900_/B sky130_fd_sc_hd__mux4_1
X_18214_ _18214_/A vssd1 vssd1 vccd1 vccd1 _19946_/D sky130_fd_sc_hd__clkbuf_1
X_15426_ _15236_/A _15423_/X _15425_/Y _15413_/X vssd1 vssd1 vccd1 vccd1 _15426_/X
+ sky130_fd_sc_hd__a31o_1
X_19194_ _19485_/CLK _19194_/D vssd1 vssd1 vccd1 vccd1 _19194_/Q sky130_fd_sc_hd__dfxtp_1
X_12638_ _12639_/A _14907_/A vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15958__B _15966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18145_ _17646_/X _19916_/Q _18147_/S vssd1 vssd1 vccd1 vccd1 _18146_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13759__A _13858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15357_ _15399_/A _15357_/B _15357_/C vssd1 vssd1 vccd1 vccd1 _15357_/X sky130_fd_sc_hd__and3_1
X_12569_ _15962_/C _18918_/Q _12687_/A vssd1 vssd1 vccd1 vccd1 _14863_/A sky130_fd_sc_hd__mux2_2
XFILLER_8_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16135__A _16135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14308_ _18668_/Q _14304_/B _14307_/Y vssd1 vssd1 vccd1 vccd1 _18668_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18076_ _18076_/A vssd1 vssd1 vccd1 vccd1 _19894_/D sky130_fd_sc_hd__clkbuf_1
X_15288_ _15302_/A _15291_/A vssd1 vssd1 vccd1 vccd1 _15288_/X sky130_fd_sc_hd__or2_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17027_ _17094_/S vssd1 vssd1 vccd1 vccd1 _17040_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__15974__A _15982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14239_ _14239_/A _14241_/B vssd1 vssd1 vccd1 vccd1 _14239_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09780_ _09780_/A vssd1 vssd1 vccd1 vccd1 _09837_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _18992_/CLK _18978_/D vssd1 vssd1 vccd1 vccd1 _18978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _19835_/Q _17058_/X _17937_/S vssd1 vssd1 vccd1 vccd1 _17930_/A sky130_fd_sc_hd__mux2_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12838__A _12838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13271__A1 _18473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09212__A input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09214_ _18828_/Q _09354_/B vssd1 vssd1 vccd1 vccd1 _09342_/B sky130_fd_sc_hd__or2_1
XFILLER_14_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11337__A1 _09559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09882__A _09882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11432__S1 _11107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_opt_1_0_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09978_ _10365_/A vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_133_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11940_ _11948_/A _11948_/B _11940_/C _11940_/D vssd1 vssd1 vccd1 vccd1 _11940_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _19904_/Q _13164_/B _11706_/A _18813_/Q vssd1 vssd1 vccd1 vccd1 _11871_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _14552_/A vssd1 vssd1 vccd1 vccd1 _13709_/A sky130_fd_sc_hd__clkbuf_2
X_10822_ _10822_/A _10822_/B vssd1 vssd1 vccd1 vccd1 _10822_/Y sky130_fd_sc_hd__nand2_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14590_/A vssd1 vssd1 vccd1 vccd1 _18765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11499__S1 _10856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13541_ _13541_/A vssd1 vssd1 vccd1 vccd1 _18458_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_1_clock clkbuf_1_1_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_10753_ _19142_/Q _19403_/Q _19302_/Q _19637_/Q _09725_/A _10638_/A vssd1 vssd1 vccd1
+ vccd1 _10753_/X sky130_fd_sc_hd__mux4_2
XFILLER_41_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15003__A2 _14996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10171__S1 _10153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16260_ _16282_/A vssd1 vssd1 vccd1 vccd1 _16269_/S sky130_fd_sc_hd__buf_4
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13014__A1 _13542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13472_ _18580_/Q _13189_/X _13469_/X _13470_/X _13471_/X vssd1 vssd1 vccd1 vccd1
+ _13472_/X sky130_fd_sc_hd__a2111o_4
X_10684_ _10695_/A _10684_/B vssd1 vssd1 vccd1 vccd1 _10684_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15211_ _15286_/A vssd1 vssd1 vccd1 vccd1 _15211_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12423_ _12399_/A _12424_/C _18772_/Q vssd1 vssd1 vccd1 vccd1 _12423_/Y sky130_fd_sc_hd__a21oi_2
X_16191_ _13250_/X _19113_/Q _16195_/S vssd1 vssd1 vccd1 vccd1 _16192_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14762__A1 _12866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12483__A _18774_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15142_ _15142_/A _15142_/B vssd1 vssd1 vccd1 vccd1 _15142_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12354_ _11904_/A _12842_/A _12353_/Y vssd1 vssd1 vccd1 vccd1 _12406_/C sky130_fd_sc_hd__a21oi_1
XFILLER_5_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15794__A _15879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ _18427_/Q _19456_/Q _19493_/Q _19067_/Q _10618_/A _11086_/A vssd1 vssd1 vccd1
+ vccd1 _11305_/X sky130_fd_sc_hd__mux4_1
X_19950_ _19950_/CLK _19950_/D vssd1 vssd1 vccd1 vccd1 _19950_/Q sky130_fd_sc_hd__dfxtp_1
X_15073_ _14923_/X _15072_/X _14984_/X vssd1 vssd1 vccd1 vccd1 _15073_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12285_ _12285_/A vssd1 vssd1 vccd1 vccd1 _13900_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18901_ _18997_/CLK _18901_/D vssd1 vssd1 vccd1 vccd1 _18901_/Q sky130_fd_sc_hd__dfxtp_2
X_14024_ _14026_/A _14026_/B _14019_/X vssd1 vssd1 vccd1 vccd1 _14024_/Y sky130_fd_sc_hd__a21oi_1
X_11236_ _19229_/Q _19724_/Q _11295_/S vssd1 vssd1 vccd1 vccd1 _11237_/B sky130_fd_sc_hd__mux2_1
XFILLER_171_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19881_ _19882_/CLK _19881_/D vssd1 vssd1 vccd1 vccd1 _19881_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10536__C1 _09806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17464__A0 _17151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold7_A hold7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10000__B2 _18858_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18832_ _18960_/CLK _18832_/D vssd1 vssd1 vccd1 vccd1 _18832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11167_ _18839_/Q vssd1 vssd1 vccd1 vccd1 _11167_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14203__A _14427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10118_ _18451_/Q _19480_/Q _19517_/Q _19091_/Q _09595_/A _10109_/X vssd1 vssd1 vccd1
+ vccd1 _10118_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18763_ _19062_/CLK _18763_/D vssd1 vssd1 vccd1 vccd1 _18763_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15975_ _19021_/Q _15954_/X _15955_/X _15974_/Y vssd1 vssd1 vccd1 vccd1 _19021_/D
+ sky130_fd_sc_hd__a22o_1
X_11098_ _11242_/A _11098_/B vssd1 vssd1 vccd1 vccd1 _11098_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17714_ _17713_/X _19743_/Q _17714_/S vssd1 vssd1 vccd1 vccd1 _17715_/A sky130_fd_sc_hd__mux2_1
X_10049_ _10049_/A vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__buf_2
X_14926_ _14924_/X _14925_/X _14938_/S vssd1 vssd1 vccd1 vccd1 _14926_/X sky130_fd_sc_hd__mux2_1
X_18694_ _19888_/CLK _18694_/D vssd1 vssd1 vccd1 vccd1 _18694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17645_ _17645_/A vssd1 vssd1 vccd1 vccd1 _19721_/D sky130_fd_sc_hd__clkbuf_1
X_14857_ _15183_/A vssd1 vssd1 vccd1 vccd1 _15068_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15242__A2 _09433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13808_ _18501_/Q _13806_/X _13820_/S vssd1 vssd1 vccd1 vccd1 _13809_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13253__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14788_ _14788_/A vssd1 vssd1 vccd1 vccd1 _18828_/D sky130_fd_sc_hd__clkbuf_1
X_17576_ _17115_/X _19692_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17577_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19315_ _19972_/CLK _19315_/D vssd1 vssd1 vccd1 vccd1 _19315_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11264__B1 _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16527_ _16527_/A vssd1 vssd1 vccd1 vccd1 _19246_/D sky130_fd_sc_hd__clkbuf_1
X_13739_ _13746_/B _13739_/B vssd1 vssd1 vccd1 vccd1 _13739_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19246_ _20031_/CLK _19246_/D vssd1 vssd1 vccd1 vccd1 _19246_/Q sky130_fd_sc_hd__dfxtp_1
X_16458_ _16458_/A vssd1 vssd1 vccd1 vccd1 _19216_/D sky130_fd_sc_hd__clkbuf_1
X_15409_ _15099_/X _15406_/Y _15408_/X _15105_/X vssd1 vssd1 vccd1 vccd1 _15412_/B
+ sky130_fd_sc_hd__a211o_1
X_19177_ _19963_/CLK _19177_/D vssd1 vssd1 vccd1 vccd1 _19177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16389_ _16389_/A vssd1 vssd1 vccd1 vccd1 _19187_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12393__A _12393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11567__A1 _09833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18128_ _18127_/X _19910_/Q _18128_/S vssd1 vssd1 vccd1 vccd1 _18129_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18059_ _18059_/A vssd1 vssd1 vccd1 vccd1 _19889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09901_ _09897_/X _09899_/X _09900_/X _09750_/A _09837_/X vssd1 vssd1 vccd1 vccd1
+ _09908_/B sky130_fd_sc_hd__o221a_1
XFILLER_99_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17455__A0 _17138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20021_ _20021_/CLK _20021_/D vssd1 vssd1 vccd1 vccd1 _20021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09832_ _10424_/A vssd1 vssd1 vccd1 vccd1 _10210_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _10438_/A vssd1 vssd1 vccd1 vccd1 _10292_/A sky130_fd_sc_hd__clkbuf_2
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12819__A1 _18788_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16739__S _16747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11178__S0 _11171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09694_ _18863_/Q _09540_/X _09547_/X _09693_/X vssd1 vssd1 vccd1 vccd1 _15980_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15879__A _15879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10816__A _15938_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16497__A1 _13787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12070_ _12020_/X _12071_/B _12071_/C vssd1 vssd1 vccd1 vccd1 _12070_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11021_ _11021_/A vssd1 vssd1 vccd1 vccd1 _11022_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10551__A _10668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14023__A _14447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15472__A2 _15474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15760_ _15760_/A _15760_/B vssd1 vssd1 vccd1 vccd1 _15760_/X sky130_fd_sc_hd__or2_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12972_ _18868_/Q vssd1 vssd1 vccd1 vccd1 _12973_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_A io_dbus_rdata[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14711_ _14711_/A vssd1 vssd1 vccd1 vccd1 _18806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11923_ _11950_/A _09316_/A _11920_/D _11921_/X _11922_/X vssd1 vssd1 vccd1 vccd1
+ _12085_/A sky130_fd_sc_hd__o311a_2
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09782__S0 _09733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15691_ _18922_/Q _12674_/A _15699_/S vssd1 vssd1 vccd1 vccd1 _15692_/A sky130_fd_sc_hd__mux2_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17430_ _17430_/A vssd1 vssd1 vccd1 vccd1 _19623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14642_ _12679_/B _11898_/X _14649_/S vssd1 vssd1 vccd1 vccd1 _14643_/B sky130_fd_sc_hd__mux2_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ _12876_/A vssd1 vssd1 vccd1 vccd1 _13189_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _19364_/Q _19699_/Q _10859_/S vssd1 vssd1 vccd1 vccd1 _10805_/X sky130_fd_sc_hd__mux2_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11246__B1 _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15789__A _15789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14573_ _12134_/B hold7/A _14581_/S vssd1 vssd1 vccd1 vccd1 _14574_/B sky130_fd_sc_hd__mux2_1
X_17361_ _19593_/Q _17001_/X _17365_/S vssd1 vssd1 vccd1 vccd1 _17362_/A sky130_fd_sc_hd__mux2_1
X_11785_ _11785_/A _11790_/B vssd1 vssd1 vccd1 vccd1 _11819_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13801__S _13804_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12994__A0 _18837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19100_ _19981_/CLK _19100_/D vssd1 vssd1 vccd1 vccd1 _19100_/Q sky130_fd_sc_hd__dfxtp_1
X_16312_ _16312_/A vssd1 vssd1 vccd1 vccd1 _19163_/D sky130_fd_sc_hd__clkbuf_1
X_13524_ _13504_/A _13523_/C _12973_/B vssd1 vssd1 vccd1 vccd1 _13524_/Y sky130_fd_sc_hd__o21ai_1
X_10736_ _09546_/A _10721_/X _10734_/X _10078_/X _10735_/Y vssd1 vssd1 vccd1 vccd1
+ _15943_/B sky130_fd_sc_hd__o32a_4
X_17292_ _17292_/A vssd1 vssd1 vccd1 vccd1 _19562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19031_ _19755_/CLK _19031_/D vssd1 vssd1 vccd1 vccd1 _19031_/Q sky130_fd_sc_hd__dfxtp_1
X_16243_ _13065_/X _19135_/Q _16247_/S vssd1 vssd1 vccd1 vccd1 _16244_/A sky130_fd_sc_hd__mux2_1
X_13455_ _14336_/B _13081_/X _11687_/X _18643_/Q vssd1 vssd1 vccd1 vccd1 _13455_/X
+ sky130_fd_sc_hd__a22o_1
X_10667_ _10674_/A _10661_/X _10666_/X _09686_/A vssd1 vssd1 vccd1 vccd1 _10668_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12406_ _12406_/A _12406_/B _12406_/C _15338_/A vssd1 vssd1 vccd1 vccd1 _12433_/B
+ sky130_fd_sc_hd__or4_2
X_16174_ _16174_/A vssd1 vssd1 vccd1 vccd1 _19105_/D sky130_fd_sc_hd__clkbuf_1
X_13386_ _13386_/A vssd1 vssd1 vccd1 vccd1 _13464_/S sky130_fd_sc_hd__buf_4
X_10598_ _19144_/Q _19405_/Q _19304_/Q _19639_/Q _10724_/S _10654_/A vssd1 vssd1 vccd1
+ vccd1 _10599_/B sky130_fd_sc_hd__mux4_1
XFILLER_154_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15125_ _15419_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15125_/X sky130_fd_sc_hd__or2_1
Xoutput108 _14813_/A vssd1 vssd1 vccd1 vccd1 io_dbus_st_type[1] sky130_fd_sc_hd__buf_2
X_12337_ _12372_/B vssd1 vssd1 vccd1 vccd1 _12338_/A sky130_fd_sc_hd__buf_2
XFILLER_56_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput119 _12850_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[19] sky130_fd_sc_hd__buf_2
XFILLER_154_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19933_ _19997_/CLK _19933_/D vssd1 vssd1 vccd1 vccd1 _19933_/Q sky130_fd_sc_hd__dfxtp_1
X_15056_ _15054_/X _15055_/X _15082_/B vssd1 vssd1 vccd1 vccd1 _15056_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12268_ _12266_/Y _18907_/Q _12409_/A vssd1 vssd1 vccd1 vccd1 _12298_/A sky130_fd_sc_hd__mux2_4
XFILLER_123_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17437__A0 _17112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13171__B1 _13166_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ _18577_/Q _18576_/Q _14007_/C vssd1 vssd1 vccd1 vccd1 _14013_/C sky130_fd_sc_hd__and3_1
X_11219_ _19196_/Q _19787_/Q _19949_/Q _19164_/Q _11063_/X _11073_/X vssd1 vssd1 vccd1
+ vccd1 _11219_/X sky130_fd_sc_hd__mux4_1
X_19864_ _19864_/CLK _19864_/D vssd1 vssd1 vccd1 vccd1 _19864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12199_ _12162_/A _12198_/X _18764_/Q _12059_/A vssd1 vssd1 vccd1 vccd1 _12255_/C
+ sky130_fd_sc_hd__o211a_2
Xoutput90 _12717_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[27] sky130_fd_sc_hd__buf_2
XFILLER_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18815_ _19910_/CLK _18815_/D vssd1 vssd1 vccd1 vccd1 _18815_/Q sky130_fd_sc_hd__dfxtp_1
X_19795_ _19976_/CLK _19795_/D vssd1 vssd1 vccd1 vccd1 _19795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18746_ _18762_/CLK _18746_/D vssd1 vssd1 vccd1 vccd1 _18746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15958_ _15966_/A _15966_/B _15958_/C vssd1 vssd1 vccd1 vccd1 _15958_/X sky130_fd_sc_hd__and3_1
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14909_ _14909_/A vssd1 vssd1 vccd1 vccd1 _15177_/B sky130_fd_sc_hd__buf_2
X_18677_ _18677_/CLK _18677_/D vssd1 vssd1 vccd1 vccd1 _18677_/Q sky130_fd_sc_hd__dfxtp_1
X_15889_ _15889_/A vssd1 vssd1 vccd1 vccd1 _18989_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15215__A2 _15219_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17628_ _17192_/X _19716_/Q _17628_/S vssd1 vssd1 vccd1 vccd1 _17629_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17559_ _17559_/A vssd1 vssd1 vccd1 vccd1 _19685_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13711__S _16066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09697__A _18827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12835__B _12835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19229_ _19726_/CLK _19229_/D vssd1 vssd1 vccd1 vccd1 _19229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12737__A0 _15976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12851__A _12851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18014__S _18020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17979__A1 _17026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20004_ _20036_/CLK _20004_/D vssd1 vssd1 vccd1 vccd1 _20004_/Q sky130_fd_sc_hd__dfxtp_1
X_09815_ _19388_/Q vssd1 vssd1 vccd1 vccd1 _09816_/A sky130_fd_sc_hd__buf_2
XANTENNA_input3_A io_dbus_rdata[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09746_ _10207_/A vssd1 vssd1 vccd1 vccd1 _09747_/A sky130_fd_sc_hd__buf_2
XFILLER_101_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09669__B1 _10073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_171_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _18773_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _19350_/Q _19621_/Q _19845_/Q _19589_/Q _09855_/A _09642_/A vssd1 vssd1 vccd1
+ vccd1 _09677_/X sky130_fd_sc_hd__mux4_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12298__A _12298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17600__A0 _17151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11571__S0 _11566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_186_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _18992_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11323__S0 _09586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13232__A4 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11570_ _19351_/Q _19622_/Q _19846_/Q _19590_/Q _11553_/X _11565_/A vssd1 vssd1 vccd1
+ vccd1 _11570_/X sky130_fd_sc_hd__mux4_2
XFILLER_156_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10521_ _10521_/A vssd1 vssd1 vccd1 vccd1 _10521_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10451__A1 _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15914__A0 hold6/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13240_ _13240_/A vssd1 vssd1 vccd1 vccd1 _18440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10452_ _19147_/Q _19408_/Q _19307_/Q _19642_/Q _10180_/S _09610_/A vssd1 vssd1 vccd1
+ vccd1 _10453_/B sky130_fd_sc_hd__mux4_1
XFILLER_136_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14193__A2 _14197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15390__A1 _12470_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13857__A _17093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ _18563_/Q _13070_/X _13166_/X _13168_/X _13170_/X vssd1 vssd1 vccd1 vccd1
+ _13609_/B sky130_fd_sc_hd__a2111o_2
X_10383_ _10484_/A _10381_/X _10382_/X vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__o21a_1
XFILLER_151_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12122_ _12120_/X _12122_/B vssd1 vssd1 vccd1 vccd1 _12215_/C sky130_fd_sc_hd__and2b_2
XFILLER_123_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input59_A io_ibus_inst[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_124_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _18923_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17763__S _17771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12053_ _12128_/C _12053_/B vssd1 vssd1 vccd1 vccd1 _12054_/D sky130_fd_sc_hd__nor2_1
X_16930_ _16930_/A vssd1 vssd1 vccd1 vccd1 _19424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ _11006_/A _11002_/X _11003_/X vssd1 vssd1 vccd1 vccd1 _11004_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__18092__A0 _18091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10062__S0 _09918_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16861_ _16918_/S vssd1 vssd1 vccd1 vccd1 _16870_/S sky130_fd_sc_hd__buf_2
XFILLER_120_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18600_ _20037_/CLK _18600_/D vssd1 vssd1 vccd1 vccd1 _18600_/Q sky130_fd_sc_hd__dfxtp_1
X_15812_ _11925_/B _11860_/A _15798_/X input62/X vssd1 vssd1 vccd1 vccd1 _15813_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_139_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18660_/CLK sky130_fd_sc_hd__clkbuf_16
X_19580_ _19644_/CLK _19580_/D vssd1 vssd1 vccd1 vccd1 _19580_/Q sky130_fd_sc_hd__dfxtp_1
X_16792_ _16792_/A vssd1 vssd1 vccd1 vccd1 _19363_/D sky130_fd_sc_hd__clkbuf_1
X_18531_ _19880_/CLK _18531_/D vssd1 vssd1 vccd1 vccd1 _18531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15743_ _15769_/A vssd1 vssd1 vccd1 vccd1 _15743_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12955_ _13936_/B _12877_/X _12951_/X _12953_/X _12954_/X vssd1 vssd1 vccd1 vccd1
+ _13505_/B sky130_fd_sc_hd__a2111o_4
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _11941_/B vssd1 vssd1 vccd1 vccd1 _12317_/A sky130_fd_sc_hd__clkinv_2
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _19885_/CLK _18462_/D vssd1 vssd1 vccd1 vccd1 _18462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _15674_/A vssd1 vssd1 vccd1 vccd1 _18914_/D sky130_fd_sc_hd__clkbuf_1
X_12886_ _19059_/Q _12878_/X _12879_/X _18757_/Q _12885_/X vssd1 vssd1 vccd1 vccd1
+ _12886_/X sky130_fd_sc_hd__a221o_2
XFILLER_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14405__B1 _14366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17413_/A vssd1 vssd1 vccd1 vccd1 _19616_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _11773_/A _11860_/C _15789_/A vssd1 vssd1 vccd1 vccd1 _14534_/S sky130_fd_sc_hd__o21a_1
X_14625_ _18776_/Q _13661_/X _14632_/S vssd1 vssd1 vccd1 vccd1 _14626_/B sky130_fd_sc_hd__mux2_1
XANTENNA__14956__A1 _15100_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18393_ _18393_/A vssd1 vssd1 vccd1 vccd1 _20026_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11840__A _15875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _17186_/X _19586_/Q _17348_/S vssd1 vssd1 vccd1 vccd1 _17345_/A sky130_fd_sc_hd__mux2_1
X_14556_ _14652_/A vssd1 vssd1 vccd1 vccd1 _14601_/A sky130_fd_sc_hd__buf_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _15875_/A vssd1 vssd1 vccd1 vccd1 _14544_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10442__A1 _09884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10719_ _10719_/A vssd1 vssd1 vccd1 vccd1 _10719_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14708__A1 _13629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15905__A0 _18995_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13507_ _11813_/X _13505_/X _13506_/Y _11831_/X _18996_/Q vssd1 vssd1 vccd1 vccd1
+ _13508_/B sky130_fd_sc_hd__a32o_4
X_17275_ _17275_/A vssd1 vssd1 vccd1 vccd1 _19555_/D sky130_fd_sc_hd__clkbuf_1
X_14487_ _14495_/A _14487_/B _14487_/C vssd1 vssd1 vccd1 vccd1 _18728_/D sky130_fd_sc_hd__nor3_1
XFILLER_174_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11699_ _11699_/A vssd1 vssd1 vccd1 vccd1 _15758_/A sky130_fd_sc_hd__buf_2
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19014_ _19055_/CLK _19014_/D vssd1 vssd1 vccd1 vccd1 _19014_/Q sky130_fd_sc_hd__dfxtp_1
X_16226_ _16282_/A vssd1 vssd1 vccd1 vccd1 _16295_/S sky130_fd_sc_hd__buf_6
X_13438_ _18578_/Q _12877_/X _13433_/X _13435_/X _13437_/X vssd1 vssd1 vccd1 vccd1
+ _13725_/B sky130_fd_sc_hd__a2111o_2
XFILLER_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15966__B _15966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16157_ _16157_/A vssd1 vssd1 vccd1 vccd1 _19097_/D sky130_fd_sc_hd__clkbuf_1
X_13369_ input18/X _13318_/X _13368_/X vssd1 vssd1 vccd1 vccd1 _13369_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12671__A _15482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ _14923_/X _15100_/B _15438_/A _15106_/X _15107_/Y vssd1 vssd1 vccd1 vccd1
+ _15108_/X sky130_fd_sc_hd__o2111a_1
XFILLER_170_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16088_ _16088_/A vssd1 vssd1 vccd1 vccd1 _19067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13144__A0 _18844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17673__S _17682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19916_ _19980_/CLK _19916_/D vssd1 vssd1 vccd1 vccd1 _19916_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15982__A _15982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15039_ _14899_/X _14902_/X _15039_/S vssd1 vssd1 vccd1 vccd1 _15039_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09899__B1 _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09980__A _09980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19847_ _19946_/CLK _19847_/D vssd1 vssd1 vccd1 vccd1 _19847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16289__S _16291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09600_ _10972_/A vssd1 vssd1 vccd1 vccd1 _10996_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19778_ _19972_/CLK _19778_/D vssd1 vssd1 vccd1 vccd1 _19778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09531_ _19487_/Q vssd1 vssd1 vccd1 vccd1 _09532_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18729_ _18731_/CLK _18729_/D vssd1 vssd1 vccd1 vccd1 _18729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09462_ _18985_/Q vssd1 vssd1 vccd1 vccd1 _09466_/A sky130_fd_sc_hd__buf_6
XFILLER_58_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14947__A1 _15177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09393_ _09401_/A _11777_/C _11707_/A vssd1 vssd1 vccd1 vccd1 _09410_/A sky130_fd_sc_hd__o21ba_2
XANTENNA__18009__S _18009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12846__A _12863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__S0 _10618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17848__S _17854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16752__S _16758_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_41_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _20022_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10736__A2 _10721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _20024_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__18074__A0 _18846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09729_ _09729_/A vssd1 vssd1 vccd1 vccd1 _10166_/S sky130_fd_sc_hd__buf_4
XANTENNA__16927__S _16931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12110__A1 _12134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11544__S0 _11534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ _12740_/A _15520_/B vssd1 vssd1 vccd1 vccd1 _12741_/B sky130_fd_sc_hd__nor2_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _15482_/A vssd1 vssd1 vccd1 vccd1 _12671_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12949__B1 _12944_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14452_/A _14410_/B _14410_/C vssd1 vssd1 vccd1 vccd1 _18698_/D sky130_fd_sc_hd__nor3_1
X_11622_ _11600_/Y _11614_/X _11622_/C _11622_/D vssd1 vssd1 vccd1 vccd1 _11622_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _12470_/Y _15364_/X _15389_/X _15360_/X vssd1 vssd1 vccd1 vccd1 _15390_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14341_ _18677_/Q _14369_/B _14340_/Y vssd1 vssd1 vccd1 vccd1 _18677_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17758__S _17760_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _11553_/A vssd1 vssd1 vccd1 vccd1 _11553_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_156_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17060_ _19473_/Q _17058_/X _17072_/S vssd1 vssd1 vccd1 vccd1 _17061_/A sky130_fd_sc_hd__mux2_1
X_10504_ _10508_/A _10504_/B vssd1 vssd1 vccd1 vccd1 _10504_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14272_ _18658_/Q _14280_/A _14275_/D vssd1 vssd1 vccd1 vccd1 _14273_/B sky130_fd_sc_hd__and3_1
XFILLER_144_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11484_ _11477_/X _11479_/X _11481_/X _11483_/X _09874_/A vssd1 vssd1 vccd1 vccd1
+ _11484_/X sky130_fd_sc_hd__a221o_2
XFILLER_7_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16011_ _16057_/S vssd1 vssd1 vccd1 vccd1 _16020_/S sky130_fd_sc_hd__buf_2
X_13223_ _13223_/A vssd1 vssd1 vccd1 vccd1 _13223_/X sky130_fd_sc_hd__buf_4
XANTENNA__13374__B1 _12944_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10435_ _18444_/Q _19473_/Q _19510_/Q _19084_/Q _10469_/S _10163_/X vssd1 vssd1 vccd1
+ vccd1 _10435_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17059__A _17075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13587__A _13656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13154_ _13245_/A _11857_/B _11857_/C _11857_/D _13153_/X vssd1 vssd1 vccd1 vccd1
+ _13154_/X sky130_fd_sc_hd__o41a_1
X_10366_ _18445_/Q _19474_/Q _19511_/Q _19085_/Q _10058_/A _10054_/A vssd1 vssd1 vccd1
+ vccd1 _10366_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output165_A _12801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12105_ _18761_/Q vssd1 vssd1 vccd1 vccd1 _12134_/B sky130_fd_sc_hd__clkbuf_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17962_ _17962_/A vssd1 vssd1 vccd1 vccd1 _19849_/D sky130_fd_sc_hd__clkbuf_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _18841_/Q _13570_/B _13360_/A vssd1 vssd1 vccd1 vccd1 _13085_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10297_ _09780_/A _10290_/Y _10292_/Y _10294_/Y _10296_/Y vssd1 vssd1 vccd1 vccd1
+ _10297_/X sky130_fd_sc_hd__o32a_1
XFILLER_111_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19701_ _19959_/CLK _19701_/D vssd1 vssd1 vccd1 vccd1 _19701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16913_ _16913_/A vssd1 vssd1 vccd1 vccd1 _19417_/D sky130_fd_sc_hd__clkbuf_1
X_12036_ _12085_/A _09495_/A _12034_/X _12035_/Y vssd1 vssd1 vccd1 vccd1 _12078_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17893_ _19819_/Q _17007_/X _17893_/S vssd1 vssd1 vccd1 vccd1 _17894_/A sky130_fd_sc_hd__mux2_1
X_19632_ _19986_/CLK _19632_/D vssd1 vssd1 vccd1 vccd1 _19632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16844_ _17201_/A _16844_/B vssd1 vssd1 vccd1 vccd1 _16845_/A sky130_fd_sc_hd__and2_1
XFILLER_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19563_ _19948_/CLK _19563_/D vssd1 vssd1 vccd1 vccd1 _19563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16775_ _16313_/X _19356_/Q _16775_/S vssd1 vssd1 vccd1 vccd1 _16776_/A sky130_fd_sc_hd__mux2_1
X_13987_ _18570_/Q _13990_/C _13969_/X vssd1 vssd1 vccd1 vccd1 _13987_/Y sky130_fd_sc_hd__a21oi_1
X_18514_ _19973_/CLK _18514_/D vssd1 vssd1 vccd1 vccd1 _18514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ _17098_/A _15732_/B vssd1 vssd1 vccd1 vccd1 _15726_/Y sky130_fd_sc_hd__nand2_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _16998_/A vssd1 vssd1 vccd1 vccd1 _17640_/A sky130_fd_sc_hd__clkbuf_2
X_19494_ _20013_/CLK _19494_/D vssd1 vssd1 vccd1 vccd1 _19494_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17040__A1 _17039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18445_ _19998_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ _15703_/S vssd1 vssd1 vccd1 vccd1 _15666_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12869_ _14938_/S vssd1 vssd1 vccd1 vccd1 _14957_/S sky130_fd_sc_hd__buf_2
XANTENNA__15042__A _15094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14608_ _12399_/A _13621_/X _14615_/S vssd1 vssd1 vccd1 vccd1 _14609_/B sky130_fd_sc_hd__mux2_1
X_18376_ _18422_/S vssd1 vssd1 vccd1 vccd1 _18385_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_159_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15588_ _15588_/A vssd1 vssd1 vccd1 vccd1 _18876_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17327_ _17327_/A vssd1 vssd1 vccd1 vccd1 _19578_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09900__S0 _11553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16572__S _16580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14539_ _16836_/A vssd1 vssd1 vccd1 vccd1 _17208_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18353__A _18409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09975__A _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17258_ _17258_/A vssd1 vssd1 vccd1 vccd1 _19547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16209_ _13385_/X _19121_/Q _16217_/S vssd1 vssd1 vccd1 vccd1 _16210_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17189_ _17726_/A vssd1 vssd1 vccd1 vccd1 _17189_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10125__S _10125_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11128__C1 _11003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12891__A2 _12889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16747__S _16747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09514_ _09514_/A _09514_/B _09514_/C _09514_/D vssd1 vssd1 vccd1 vccd1 _09514_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_83_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10103__B1 _09913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17031__A1 _17030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09445_ _15786_/B vssd1 vssd1 vccd1 vccd1 _13518_/A sky130_fd_sc_hd__clkbuf_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09376_ _18956_/Q vssd1 vssd1 vccd1 vccd1 _15775_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17578__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14791__A _14791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16482__S _16486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09885__A _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15345__A1 _18847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12159__A1 _18460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14553__C1 _11717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__A _10824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10220_ _10480_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _10220_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10265__S0 _09657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13108__A0 _18842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10151_ _10574_/S vssd1 vssd1 vccd1 vccd1 _10208_/A sky130_fd_sc_hd__buf_2
XFILLER_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10035__S _10037_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18202__S _18202_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _10082_/A vssd1 vssd1 vccd1 vccd1 _10278_/A sky130_fd_sc_hd__buf_2
XFILLER_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10568__S1 _10011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ _13910_/A vssd1 vssd1 vccd1 vccd1 _14792_/A sky130_fd_sc_hd__buf_6
XFILLER_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14890_ _15020_/A vssd1 vssd1 vccd1 vccd1 _15118_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13841_ _13841_/A vssd1 vssd1 vccd1 vccd1 _18511_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16657__S _16663_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14966__A _14966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13870__A _14529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13772_ _18490_/Q _13771_/X _13772_/S vssd1 vssd1 vccd1 vccd1 _13773_/A sky130_fd_sc_hd__mux2_1
X_16560_ _16617_/S vssd1 vssd1 vccd1 vccd1 _16569_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_28_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10984_ _10775_/A _10979_/Y _10982_/Y _10983_/X vssd1 vssd1 vccd1 vccd1 _10984_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15511_ _15522_/A _15511_/B _15511_/C vssd1 vssd1 vccd1 vccd1 _15511_/X sky130_fd_sc_hd__and3_1
X_12723_ _12522_/A _12721_/X _12722_/X _12480_/X vssd1 vssd1 vccd1 vccd1 _12723_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16491_ _19230_/Q _13778_/X _16497_/S vssd1 vssd1 vccd1 vccd1 _16492_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10740__S1 _10626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12917__C _16150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18230_ _19954_/Q _17665_/A _18230_/S vssd1 vssd1 vccd1 vccd1 _18231_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12654_ _12679_/B _12679_/C vssd1 vssd1 vccd1 vccd1 _12654_/X sky130_fd_sc_hd__or2_1
X_15442_ _18854_/Q _15441_/X _15480_/S vssd1 vssd1 vccd1 vccd1 _15443_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17488__S _17492_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11605_ _11605_/A _11605_/B vssd1 vssd1 vccd1 vccd1 _11614_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18161_ _17668_/X _19923_/Q _18169_/S vssd1 vssd1 vccd1 vccd1 _18162_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12585_ _18539_/Q _12553_/X _12580_/X _12584_/Y vssd1 vssd1 vccd1 vccd1 _12585_/X
+ sky130_fd_sc_hd__o22a_4
X_15373_ _15373_/A _15373_/B vssd1 vssd1 vccd1 vccd1 _15373_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_128_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17112_ _17649_/A vssd1 vssd1 vccd1 vccd1 _17112_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11536_ _11547_/A _11531_/X _11533_/Y _11535_/Y vssd1 vssd1 vccd1 vccd1 _11536_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_14324_ _14327_/B _14327_/C _18673_/Q vssd1 vssd1 vccd1 vccd1 _14326_/B sky130_fd_sc_hd__a21oi_1
XFILLER_157_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18092_ _18091_/X _19899_/Q _18095_/S vssd1 vssd1 vccd1 vccd1 _18093_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17043_ _17075_/A vssd1 vssd1 vccd1 vccd1 _17056_/S sky130_fd_sc_hd__buf_2
X_14255_ _18653_/Q _18652_/Q vssd1 vssd1 vccd1 vccd1 _14256_/D sky130_fd_sc_hd__and2_1
XFILLER_156_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11467_ _19365_/Q _19700_/Q _11467_/S vssd1 vssd1 vccd1 vccd1 _11467_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13898__A1 _18539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13206_ _18880_/Q vssd1 vssd1 vccd1 vccd1 _13207_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10418_ _10411_/Y _10413_/Y _10415_/Y _10417_/Y _10502_/A vssd1 vssd1 vccd1 vccd1
+ _10418_/X sky130_fd_sc_hd__o221a_1
XANTENNA__10256__S0 _09967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14186_ _18634_/Q _14188_/C _14185_/Y vssd1 vssd1 vccd1 vccd1 _18634_/D sky130_fd_sc_hd__o21a_1
X_11398_ _19914_/Q _19528_/Q _19978_/Q _19097_/Q _11356_/X _11357_/X vssd1 vssd1 vccd1
+ vccd1 _11399_/B sky130_fd_sc_hd__mux4_1
XFILLER_98_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13137_ _17668_/A vssd1 vssd1 vccd1 vccd1 _13137_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10349_ _18855_/Q _09843_/X _09884_/A _10348_/X vssd1 vssd1 vccd1 vccd1 _12854_/B
+ sky130_fd_sc_hd__o2bb2a_4
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18994_ _18994_/CLK _18994_/D vssd1 vssd1 vccd1 vccd1 _18994_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18038__A0 _18037_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _17945_/A vssd1 vssd1 vccd1 vccd1 _19842_/D sky130_fd_sc_hd__clkbuf_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14311__A2 _14317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13068_ _13145_/A vssd1 vssd1 vccd1 vccd1 _13068_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12019_ _12059_/A vssd1 vssd1 vccd1 vccd1 _12168_/S sky130_fd_sc_hd__buf_2
XFILLER_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17876_ _19812_/Q _17087_/X _17876_/S vssd1 vssd1 vccd1 vccd1 _17877_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19615_ _19839_/CLK _19615_/D vssd1 vssd1 vccd1 vccd1 _19615_/Q sky130_fd_sc_hd__dfxtp_1
X_16827_ _16827_/A vssd1 vssd1 vccd1 vccd1 _19379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18993__D input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16567__S _16569_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19546_ _19706_/CLK _19546_/D vssd1 vssd1 vccd1 vccd1 _19546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16758_ _19349_/Q _13851_/X _16758_/S vssd1 vssd1 vccd1 vccd1 _16759_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10636__A1 _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15709_ _18930_/Q _15705_/X _15708_/X vssd1 vssd1 vccd1 vccd1 _18930_/D sky130_fd_sc_hd__a21o_1
XFILLER_62_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19477_ _19839_/CLK _19477_/D vssd1 vssd1 vccd1 vccd1 _19477_/Q sky130_fd_sc_hd__dfxtp_1
X_16689_ _16399_/X _19319_/Q _16689_/S vssd1 vssd1 vccd1 vccd1 _16690_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12396__A _16066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09230_ _09230_/A _09283_/A _11919_/A vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__or3_1
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18428_ _20013_/CLK _18428_/D vssd1 vssd1 vccd1 vccd1 _18428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17398__S _17398_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18359_ _17643_/X _20011_/Q _18363_/S vssd1 vssd1 vccd1 vccd1 _18360_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15327__A1 _12364_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10495__S0 _09653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12843__B _12844_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13889__A1 _12416_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11459__B _12834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17427__A _17483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09994_ _10129_/S vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__buf_4
XANTENNA__18022__S _18024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10349__A1_N _18855_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17861__S _17865_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10875__A1 _09664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15802__A2 _11860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09428_ _09444_/A _12064_/B _09443_/B vssd1 vssd1 vccd1 vccd1 _12918_/B sky130_fd_sc_hd__and3_4
XFILLER_13_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10538__B _12849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ _12061_/A _12066_/A vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17101__S _17113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12370_ _12279_/A _12279_/B _12279_/C _12364_/Y vssd1 vssd1 vccd1 vccd1 _12370_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12753__B _12863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11321_ _11199_/A _11318_/X _11320_/X _11332_/A vssd1 vssd1 vccd1 vccd1 _11321_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16940__S _16942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14040_ _14042_/A _14042_/C _14019_/X vssd1 vssd1 vccd1 vccd1 _14040_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11252_ _11252_/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11252_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10203_ _10196_/X _10198_/X _10200_/X _10202_/X _09876_/A vssd1 vssd1 vccd1 vccd1
+ _10203_/X sky130_fd_sc_hd__a221o_1
XANTENNA__10789__S1 _10788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11183_ _11174_/Y _11176_/Y _11179_/Y _11182_/Y _09817_/A vssd1 vssd1 vccd1 vccd1
+ _11183_/X sky130_fd_sc_hd__o221a_1
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10134_ _19155_/Q _19416_/Q _19315_/Q _19650_/Q _09653_/A _10542_/A vssd1 vssd1 vccd1
+ vccd1 _10135_/B sky130_fd_sc_hd__mux4_1
XANTENNA_input41_A io_ibus_inst[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15991_ _15991_/A vssd1 vssd1 vccd1 vccd1 _19026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17771__S _17771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17730_ _17729_/X _19748_/Q _17730_/S vssd1 vssd1 vccd1 vccd1 _17731_/A sky130_fd_sc_hd__mux2_1
X_10065_ _19344_/Q _19615_/Q _19839_/Q _19583_/Q _09597_/A _10054_/X vssd1 vssd1 vccd1
+ vccd1 _10065_/X sky130_fd_sc_hd__mux4_1
X_14942_ _15094_/A vssd1 vssd1 vccd1 vccd1 _15165_/S sky130_fd_sc_hd__buf_2
XFILLER_48_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_54_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10866__A1 _10843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10410__S0 _09995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17661_ _17661_/A vssd1 vssd1 vccd1 vccd1 _19726_/D sky130_fd_sc_hd__clkbuf_1
X_14873_ _15029_/A vssd1 vssd1 vccd1 vccd1 _15032_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__14696__A _14742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19400_ _20020_/CLK _19400_/D vssd1 vssd1 vccd1 vccd1 _19400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13804__S _13804_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16612_ _16612_/A vssd1 vssd1 vccd1 vccd1 _19284_/D sky130_fd_sc_hd__clkbuf_1
X_13824_ _18506_/Q _13822_/X _13836_/S vssd1 vssd1 vccd1 vccd1 _13825_/A sky130_fd_sc_hd__mux2_1
X_17592_ _17592_/A vssd1 vssd1 vccd1 vccd1 _19699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19331_ _19732_/CLK _19331_/D vssd1 vssd1 vccd1 vccd1 _19331_/Q sky130_fd_sc_hd__dfxtp_1
X_16543_ _19254_/Q _13854_/X _16545_/S vssd1 vssd1 vccd1 vccd1 _16544_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13755_ _17098_/A _17098_/B _16846_/C vssd1 vssd1 vccd1 vccd1 _18280_/A sky130_fd_sc_hd__or3_1
X_10967_ _09702_/A _10950_/X _10966_/X _09842_/A _18842_/Q vssd1 vssd1 vccd1 vccd1
+ _12835_/B sky130_fd_sc_hd__a32o_4
XFILLER_16_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11507__A2_N _09843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09302__B _18938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12706_ _12706_/A vssd1 vssd1 vccd1 vccd1 _15509_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19262_ _19853_/CLK _19262_/D vssd1 vssd1 vccd1 vccd1 _19262_/Q sky130_fd_sc_hd__dfxtp_1
X_16474_ _16691_/A _16474_/B _16298_/C vssd1 vssd1 vccd1 vccd1 _17635_/A sky130_fd_sc_hd__or3b_2
XFILLER_31_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10898_ _10900_/A _10897_/X _09774_/A vssd1 vssd1 vccd1 vccd1 _10898_/X sky130_fd_sc_hd__o21a_1
X_13686_ _13650_/X _13685_/X _13517_/A vssd1 vssd1 vccd1 vccd1 _13686_/X sky130_fd_sc_hd__a21bo_1
XFILLER_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13568__A0 _18461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18213_ _19946_/Q _17640_/A _18219_/S vssd1 vssd1 vccd1 vccd1 _18214_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15425_ _15142_/A _15420_/Y _15424_/Y vssd1 vssd1 vccd1 vccd1 _15425_/Y sky130_fd_sc_hd__a21oi_1
X_19193_ _19946_/CLK _19193_/D vssd1 vssd1 vccd1 vccd1 _19193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12637_ _10104_/A _18921_/Q _12805_/S vssd1 vssd1 vccd1 vccd1 _14907_/A sky130_fd_sc_hd__mux2_4
XANTENNA__15958__C _15958_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18144_ _18144_/A vssd1 vssd1 vccd1 vccd1 _19915_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12240__A0 _12239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15356_ _15305_/X _15350_/Y _15355_/Y vssd1 vssd1 vccd1 vccd1 _15357_/C sky130_fd_sc_hd__a21oi_1
X_12568_ _12568_/A _15436_/A vssd1 vssd1 vccd1 vccd1 _12571_/A sky130_fd_sc_hd__xnor2_1
XFILLER_102_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17946__S _17948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11519_ _15962_/C _12853_/B vssd1 vssd1 vccd1 vccd1 _11519_/X sky130_fd_sc_hd__and2_1
X_14307_ _14319_/A _14317_/D vssd1 vssd1 vccd1 vccd1 _14307_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18075_ _18074_/X _19894_/Q _18078_/S vssd1 vssd1 vccd1 vccd1 _18076_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12499_ _18536_/Q vssd1 vssd1 vccd1 vccd1 _12501_/B sky130_fd_sc_hd__buf_2
X_15287_ _15369_/A vssd1 vssd1 vccd1 vccd1 _15287_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17026_ _17026_/A vssd1 vssd1 vccd1 vccd1 _17026_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15974__B _15974_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14238_ _18648_/Q _14242_/C _14242_/D vssd1 vssd1 vccd1 vccd1 _14241_/B sky130_fd_sc_hd__and3_1
XFILLER_171_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13775__A _13858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14169_ _18628_/Q _14172_/C _14160_/X vssd1 vssd1 vccd1 vccd1 _14169_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _19523_/CLK _18977_/D vssd1 vssd1 vccd1 vccd1 _18977_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17928_ _17939_/A vssd1 vssd1 vccd1 vccd1 _17937_/S sky130_fd_sc_hd__buf_4
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17859_ _19804_/Q _17062_/X _17865_/S vssd1 vssd1 vccd1 vccd1 _17860_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19529_ _19979_/CLK _19529_/D vssd1 vssd1 vccd1 vccd1 _19529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13271__A2 _11755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ _18830_/Q _18829_/Q vssd1 vssd1 vccd1 vccd1 _09354_/B sky130_fd_sc_hd__or2_1
XFILLER_14_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12854__A _12857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16326__A _17662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16760__S _16762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12534__A1 _18537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ _10411_/A vssd1 vssd1 vccd1 vccd1 _10365_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17591__S _17595_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11409__S _11409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_5_0_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_clock clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11870_ _11870_/A vssd1 vssd1 vccd1 vccd1 _12982_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10821_ _19235_/Q _19730_/Q _10821_/S vssd1 vssd1 vccd1 vccd1 _10822_/B sky130_fd_sc_hd__mux2_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10752_ _10638_/X _10749_/X _10751_/X vssd1 vssd1 vccd1 vccd1 _10752_/Y sky130_fd_sc_hd__a21oi_1
X_13540_ _18458_/Q _13538_/X _13575_/S vssd1 vssd1 vccd1 vccd1 _13541_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13471_ _18612_/Q _13120_/X _11776_/X _18744_/Q vssd1 vssd1 vccd1 vccd1 _13471_/X
+ sky130_fd_sc_hd__a22o_1
X_10683_ _19928_/Q _19542_/Q _19992_/Q _19111_/Q _10521_/A _10638_/X vssd1 vssd1 vccd1
+ vccd1 _10684_/B sky130_fd_sc_hd__mux4_1
XFILLER_139_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12422_ _13508_/A vssd1 vssd1 vccd1 vccd1 _12422_/X sky130_fd_sc_hd__clkbuf_4
X_15210_ _15219_/A _15219_/B vssd1 vssd1 vccd1 vccd1 _15210_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10459__S0 _09995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16190_ _16190_/A vssd1 vssd1 vccd1 vccd1 _19112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12353_ _12859_/A _12428_/A _12318_/Y vssd1 vssd1 vccd1 vccd1 _12353_/Y sky130_fd_sc_hd__a21oi_1
X_15141_ _15077_/X _15142_/B _15140_/X _14855_/A vssd1 vssd1 vccd1 vccd1 _15141_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__16670__S _16674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11304_ _19916_/Q _19530_/Q _19980_/Q _19099_/Q _11158_/S _11108_/X vssd1 vssd1 vccd1
+ vccd1 _11304_/X sky130_fd_sc_hd__mux4_1
X_15072_ _14979_/X _15041_/X _15132_/S vssd1 vssd1 vccd1 vccd1 _15072_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12284_ _12283_/A _12309_/C _12283_/Y _12344_/A vssd1 vssd1 vccd1 vccd1 _12284_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_154_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18900_ _18997_/CLK _18900_/D vssd1 vssd1 vccd1 vccd1 _18900_/Q sky130_fd_sc_hd__dfxtp_1
X_14023_ _14447_/B _14026_/A vssd1 vssd1 vccd1 vccd1 _18582_/D sky130_fd_sc_hd__nor2_1
X_11235_ _19660_/Q _19426_/Q _18491_/Q _19756_/Q _11156_/S _11172_/X vssd1 vssd1 vccd1
+ vccd1 _11235_/X sky130_fd_sc_hd__mux4_1
X_19880_ _19880_/CLK _19880_/D vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18831_ _18960_/CLK _18831_/D vssd1 vssd1 vccd1 vccd1 _18831_/Q sky130_fd_sc_hd__dfxtp_1
X_11166_ _11166_/A _11166_/B _11166_/C vssd1 vssd1 vccd1 vccd1 _11166_/Y sky130_fd_sc_hd__nor3_1
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10117_ _10312_/A _10117_/B vssd1 vssd1 vccd1 vccd1 _10117_/Y sky130_fd_sc_hd__nor2_1
X_18762_ _18762_/CLK _18762_/D vssd1 vssd1 vccd1 vccd1 _18762_/Q sky130_fd_sc_hd__dfxtp_1
X_15974_ _15982_/A _15974_/B vssd1 vssd1 vccd1 vccd1 _15974_/Y sky130_fd_sc_hd__nor2_1
X_11097_ _19920_/Q _19534_/Q _19984_/Q _19103_/Q _11023_/S _11296_/A vssd1 vssd1 vccd1
+ vccd1 _11098_/B sky130_fd_sc_hd__mux4_1
XFILLER_76_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17713_ _17713_/A vssd1 vssd1 vccd1 vccd1 _17713_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10048_ _10048_/A vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__buf_2
X_14925_ _12519_/A _15321_/B _14933_/S vssd1 vssd1 vccd1 vccd1 _14925_/X sky130_fd_sc_hd__mux2_1
X_18693_ _18693_/CLK _18693_/D vssd1 vssd1 vccd1 vccd1 _18693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17644_ _17643_/X _19721_/Q _17650_/S vssd1 vssd1 vccd1 vccd1 _17645_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15778__A1 _09471_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14856_ _14835_/Y _15346_/A _15489_/A _14847_/X _14855_/Y vssd1 vssd1 vccd1 vccd1
+ _14856_/X sky130_fd_sc_hd__o32a_1
XFILLER_91_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ _13839_/A vssd1 vssd1 vccd1 vccd1 _13820_/S sky130_fd_sc_hd__buf_4
XFILLER_63_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17575_ _17632_/S vssd1 vssd1 vccd1 vccd1 _17584_/S sky130_fd_sc_hd__buf_2
X_14787_ _14800_/A _14787_/B vssd1 vssd1 vccd1 vccd1 _14788_/A sky130_fd_sc_hd__and2_1
XFILLER_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _11999_/A vssd1 vssd1 vccd1 vccd1 _12279_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_19314_ _19942_/CLK _19314_/D vssd1 vssd1 vccd1 vccd1 _19314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16526_ _19246_/Q _13829_/X _16530_/S vssd1 vssd1 vccd1 vccd1 _16527_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13738_ _13737_/A _13737_/C _18895_/Q vssd1 vssd1 vccd1 vccd1 _13739_/B sky130_fd_sc_hd__o21ai_1
XFILLER_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19245_ _19836_/CLK _19245_/D vssd1 vssd1 vccd1 vccd1 _19245_/Q sky130_fd_sc_hd__dfxtp_1
X_16457_ _19216_/Q _13835_/X _16457_/S vssd1 vssd1 vccd1 vccd1 _16458_/A sky130_fd_sc_hd__mux2_1
X_13669_ _13664_/Y _13667_/X _18130_/S vssd1 vssd1 vccd1 vccd1 _13669_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15408_ _15155_/X _15410_/B _15102_/X _15407_/X vssd1 vssd1 vccd1 vccd1 _15408_/X
+ sky130_fd_sc_hd__o211a_1
X_19176_ _20025_/CLK _19176_/D vssd1 vssd1 vccd1 vccd1 _19176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16388_ _16387_/X _19187_/Q _16394_/S vssd1 vssd1 vccd1 vccd1 _16389_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15950__A1 _19010_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17676__S _17682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13961__B1 _11884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18127_ _18862_/Q _13733_/X _18130_/S vssd1 vssd1 vccd1 vccd1 _18127_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17152__A0 _17151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15339_ _15305_/X _15334_/Y _15338_/Y vssd1 vssd1 vccd1 vccd1 _15340_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__16580__S _16580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__A _10194_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18058_ _18057_/X _19889_/Q _18061_/S vssd1 vssd1 vccd1 vccd1 _18059_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10870__S0 _10919_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09900_ _19684_/Q _19450_/Q _18515_/Q _19780_/Q _11553_/A _09826_/A vssd1 vssd1 vccd1
+ vccd1 _09900_/X sky130_fd_sc_hd__mux4_1
X_17009_ _17009_/A vssd1 vssd1 vccd1 vccd1 _19457_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15196__S _15480_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20020_ _20020_/CLK _20020_/D vssd1 vssd1 vccd1 vccd1 _20020_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09396__D_N _18950_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ _10690_/A vssd1 vssd1 vccd1 vccd1 _10424_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09762_ _10001_/A vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__buf_2
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18300__S _18302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11178__S1 _11172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09693_ _09862_/A _09645_/X _09692_/X vssd1 vssd1 vccd1 vccd1 _09693_/X sky130_fd_sc_hd__a21bo_1
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12849__A _12851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13492__A2 _11683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13444__S _13464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13229__C1 _13307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12568__B _15436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10369__A _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11255__A1 _11003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15941__A1 _19007_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13401__C1 _13399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10816__B _12841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10832__A _10832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10518__B1 _10162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14304__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _11388_/A vssd1 vssd1 vccd1 vccd1 _11021_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _13360_/A _18836_/Q _11796_/X _12970_/X vssd1 vssd1 vccd1 vccd1 _12971_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _18806_/Q _11724_/X _14716_/S vssd1 vssd1 vccd1 vccd1 _14711_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11961_/A _11919_/C _09276_/X _14819_/A _11931_/C vssd1 vssd1 vccd1 vccd1
+ _11922_/X sky130_fd_sc_hd__o311a_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09782__S1 _09768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15690_ _15690_/A vssd1 vssd1 vccd1 vccd1 _15699_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _14641_/A vssd1 vssd1 vccd1 vccd1 _18780_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11853_ _18594_/Q _11851_/X _11852_/X _18626_/Q vssd1 vssd1 vccd1 vccd1 _11857_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10279__A _10279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10804_ _10858_/A _10804_/B vssd1 vssd1 vccd1 vccd1 _10804_/Y sky130_fd_sc_hd__nor2_1
X_17360_ _17360_/A vssd1 vssd1 vccd1 vccd1 _19592_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11246__A1 _09702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ _13048_/B vssd1 vssd1 vccd1 vccd1 _13269_/A sky130_fd_sc_hd__clkbuf_2
X_14572_ _14572_/A vssd1 vssd1 vccd1 vccd1 _18760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11246__B2 _18838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11341__S1 _11108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16311_ _16310_/X _19163_/Q _16314_/S vssd1 vssd1 vccd1 vccd1 _16312_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11797__A2 _11776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12994__A1 _13529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13523_ _18867_/Q _18868_/Q _13523_/C vssd1 vssd1 vccd1 vccd1 _13535_/B sky130_fd_sc_hd__or3_1
XFILLER_158_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ _18847_/Q vssd1 vssd1 vccd1 vccd1 _10735_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17291_ _17109_/X _19562_/Q _17293_/S vssd1 vssd1 vccd1 vccd1 _17292_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19030_ _20013_/CLK _19030_/D vssd1 vssd1 vccd1 vccd1 _19030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16242_ _16242_/A vssd1 vssd1 vccd1 vccd1 _19134_/D sky130_fd_sc_hd__clkbuf_1
X_10666_ _10832_/A _10666_/B vssd1 vssd1 vccd1 vccd1 _10666_/X sky130_fd_sc_hd__or2_1
X_13454_ _18675_/Q vssd1 vssd1 vccd1 vccd1 _14336_/B sky130_fd_sc_hd__buf_2
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11549__A2 _11548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17496__S _17496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ _11904_/X _12844_/A _12404_/Y vssd1 vssd1 vccd1 vccd1 _15355_/A sky130_fd_sc_hd__a21oi_4
X_13385_ _17716_/A vssd1 vssd1 vccd1 vccd1 _13385_/X sky130_fd_sc_hd__clkbuf_2
X_16173_ _13115_/X _19105_/Q _16173_/S vssd1 vssd1 vccd1 vccd1 _16174_/A sky130_fd_sc_hd__mux2_1
X_10597_ _10597_/A vssd1 vssd1 vccd1 vccd1 _10654_/A sky130_fd_sc_hd__buf_2
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15124_ _15116_/X _15123_/X _15171_/S vssd1 vssd1 vccd1 vccd1 _15125_/B sky130_fd_sc_hd__mux2_2
Xoutput109 _12822_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[0] sky130_fd_sc_hd__buf_2
XFILLER_115_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12336_ _18530_/Q vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_127_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19932_ _19996_/CLK _19932_/D vssd1 vssd1 vccd1 vccd1 _19932_/Q sky130_fd_sc_hd__dfxtp_1
X_12267_ _12358_/S vssd1 vssd1 vccd1 vccd1 _12409_/A sky130_fd_sc_hd__buf_2
X_15055_ _14957_/X _14946_/X _15055_/S vssd1 vssd1 vccd1 vccd1 _15055_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output72_A _12273_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ _11257_/A _11218_/B vssd1 vssd1 vccd1 vccd1 _11218_/Y sky130_fd_sc_hd__nor2_1
X_14006_ _18576_/Q _14007_/C _18577_/Q vssd1 vssd1 vccd1 vccd1 _14008_/B sky130_fd_sc_hd__a21oi_1
X_19863_ _19976_/CLK _19863_/D vssd1 vssd1 vccd1 vccd1 _19863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12198_ _12135_/X _12164_/X _12165_/X _12167_/A vssd1 vssd1 vccd1 vccd1 _12198_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput80 _12498_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[18] sky130_fd_sc_hd__buf_2
XANTENNA__11182__B1 _11181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput91 _12743_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[28] sky130_fd_sc_hd__buf_2
XANTENNA__11049__S _11049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18814_ _19912_/CLK _18814_/D vssd1 vssd1 vccd1 vccd1 _18814_/Q sky130_fd_sc_hd__dfxtp_1
X_11149_ _11149_/A _11149_/B vssd1 vssd1 vccd1 vccd1 _11149_/Y sky130_fd_sc_hd__nor2_1
X_19794_ _20020_/CLK _19794_/D vssd1 vssd1 vccd1 vccd1 _19794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13459__C1 _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18745_ _18745_/CLK _18745_/D vssd1 vssd1 vccd1 vccd1 _18745_/Q sky130_fd_sc_hd__dfxtp_1
X_15957_ _19012_/Q _15954_/X _15955_/X _15956_/Y vssd1 vssd1 vccd1 vccd1 _19012_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13474__A2 _13472_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__A1 _09848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ _15219_/B _15474_/B _14908_/S vssd1 vssd1 vccd1 vccd1 _14908_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11485__B2 _18846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18676_ _18677_/CLK _18676_/D vssd1 vssd1 vccd1 vccd1 _18676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15888_ _15897_/A _15888_/B vssd1 vssd1 vccd1 vccd1 _15889_/A sky130_fd_sc_hd__and2_1
XFILLER_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17627_ _17627_/A vssd1 vssd1 vccd1 vccd1 _19715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14839_ _14993_/C vssd1 vssd1 vccd1 vccd1 _14990_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17558_ _19685_/Q vssd1 vssd1 vccd1 vccd1 _17559_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_149_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16509_ _16509_/A vssd1 vssd1 vccd1 vccd1 _19238_/D sky130_fd_sc_hd__clkbuf_1
X_17489_ _17489_/A vssd1 vssd1 vccd1 vccd1 _19650_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10917__A _15934_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19228_ _19949_/CLK _19228_/D vssd1 vssd1 vccd1 vccd1 _19228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_176_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19159_ _19856_/CLK _19159_/D vssd1 vssd1 vccd1 vccd1 _19159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12851__B _12851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20003_ _20003_/CLK _20003_/D vssd1 vssd1 vccd1 vccd1 _20003_/Q sky130_fd_sc_hd__dfxtp_1
X_09814_ _09957_/A _09814_/B vssd1 vssd1 vccd1 vccd1 _09814_/X sky130_fd_sc_hd__or2_1
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09745_ _09745_/A vssd1 vssd1 vccd1 vccd1 _10207_/A sky130_fd_sc_hd__buf_4
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09669__A1 _11533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14662__A1 _13742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _10073_/A vssd1 vssd1 vccd1 vccd1 _11543_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11571__S1 _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11323__S1 _11322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12976__B2 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10827__A _10832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10520_ _10520_/A _10520_/B vssd1 vssd1 vccd1 vccd1 _10520_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10451_ _10458_/A _10446_/X _10448_/X _10450_/X vssd1 vssd1 vccd1 vccd1 _10451_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11087__S0 _11023_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13170_ _18659_/Q _13081_/X _13194_/A _14485_/A vssd1 vssd1 vccd1 vccd1 _13170_/X
+ sky130_fd_sc_hd__a22o_1
X_10382_ _10382_/A vssd1 vssd1 vccd1 vccd1 _10382_/X sky130_fd_sc_hd__buf_2
XFILLER_108_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ _12121_/A _14912_/A vssd1 vssd1 vccd1 vccd1 _12122_/B sky130_fd_sc_hd__or2_1
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09357__B1 _09347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ _18521_/Q _12052_/B vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14969__A _15553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ _11003_/A vssd1 vssd1 vccd1 vccd1 _11003_/X sky130_fd_sc_hd__buf_2
XFILLER_132_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10062__S1 _09646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16860_ _16860_/A vssd1 vssd1 vccd1 vccd1 _19393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15811_ _15811_/A vssd1 vssd1 vccd1 vccd1 _18966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16791_ _16336_/X _19363_/Q _16797_/S vssd1 vssd1 vccd1 vccd1 _16792_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18530_ _18867_/CLK _18530_/D vssd1 vssd1 vccd1 vccd1 _18530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15742_ _18943_/Q _15745_/B vssd1 vssd1 vccd1 vccd1 _15742_/X sky130_fd_sc_hd__or2_1
XFILLER_58_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _18648_/Q _11889_/X _12890_/X _18716_/Q vssd1 vssd1 vccd1 vccd1 _12954_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _18993_/CLK _18461_/D vssd1 vssd1 vccd1 vccd1 _18461_/Q sky130_fd_sc_hd__dfxtp_1
X_11905_ _14821_/A _11904_/X _09338_/X _14758_/A vssd1 vssd1 vccd1 vccd1 _11905_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15673_ _18914_/Q _12501_/A _15677_/S vssd1 vssd1 vccd1 vccd1 _15674_/A sky130_fd_sc_hd__mux2_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ _18790_/Q _12880_/X _12881_/X _14345_/B _12884_/X vssd1 vssd1 vccd1 vccd1
+ _12885_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17412_ _19616_/Q _17074_/X _17420_/S vssd1 vssd1 vccd1 vccd1 _17413_/A sky130_fd_sc_hd__mux2_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09798__A _09798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14624_ _14624_/A vssd1 vssd1 vccd1 vccd1 _18775_/D sky130_fd_sc_hd__clkbuf_1
X_18392_ _17691_/X _20026_/Q _18396_/S vssd1 vssd1 vccd1 vccd1 _18393_/A sky130_fd_sc_hd__mux2_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _11915_/B vssd1 vssd1 vccd1 vccd1 _15789_/A sky130_fd_sc_hd__buf_2
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17343_/A vssd1 vssd1 vccd1 vccd1 _19585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14555_ _14672_/B _14555_/B vssd1 vssd1 vccd1 vccd1 _14652_/A sky130_fd_sc_hd__and2_2
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10737__A _15943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ _15856_/A vssd1 vssd1 vccd1 vccd1 _15875_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _13726_/A _18996_/Q vssd1 vssd1 vccd1 vccd1 _13506_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14169__B1 _14160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10718_ _20023_/Q _19861_/Q _19270_/Q _19040_/Q _10764_/S _09606_/A vssd1 vssd1 vccd1
+ vccd1 _10718_/X sky130_fd_sc_hd__mux4_1
X_17274_ _17189_/X _19555_/Q _17276_/S vssd1 vssd1 vccd1 vccd1 _17275_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14486_ _14485_/A _14485_/C _18728_/Q vssd1 vssd1 vccd1 vccd1 _14487_/C sky130_fd_sc_hd__a21oi_1
X_11698_ _11785_/A _11712_/B vssd1 vssd1 vccd1 vccd1 _11698_/Y sky130_fd_sc_hd__nor2_1
X_19013_ _19023_/CLK _19013_/D vssd1 vssd1 vccd1 vccd1 _19013_/Q sky130_fd_sc_hd__dfxtp_1
X_16225_ _16692_/A _17426_/B vssd1 vssd1 vccd1 vccd1 _16282_/A sky130_fd_sc_hd__or2_4
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13437_ _18674_/Q _11889_/X _13194_/X _14526_/B vssd1 vssd1 vccd1 vccd1 _13437_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11078__S0 _11121_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10649_ _09820_/A _10636_/X _10648_/X vssd1 vssd1 vccd1 vccd1 _10649_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15966__C _15966_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16156_ _12939_/X _19097_/Q _16162_/S vssd1 vssd1 vccd1 vccd1 _16157_/A sky130_fd_sc_hd__mux2_1
X_13368_ _13368_/A vssd1 vssd1 vccd1 vccd1 _13368_/X sky130_fd_sc_hd__buf_2
XFILLER_114_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15107_ _15181_/A _15107_/B vssd1 vssd1 vccd1 vccd1 _15107_/Y sky130_fd_sc_hd__nand2_1
X_12319_ _11667_/A _12428_/A _12318_/Y vssd1 vssd1 vccd1 vccd1 _12319_/Y sky130_fd_sc_hd__a21oi_1
X_16087_ _12978_/X _19067_/Q _16089_/S vssd1 vssd1 vccd1 vccd1 _16088_/A sky130_fd_sc_hd__mux2_1
X_13299_ input13/X _13231_/X _13234_/X vssd1 vssd1 vccd1 vccd1 _13299_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_114_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13144__A1 _11828_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19915_ _19979_/CLK _19915_/D vssd1 vssd1 vccd1 vccd1 _19915_/Q sky130_fd_sc_hd__dfxtp_1
X_15038_ _15036_/X _15037_/X _15041_/S vssd1 vssd1 vccd1 vccd1 _15038_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15982__B _15982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09899__A1 _09833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14892__A1 _12753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19846_ _19846_/CLK _19846_/D vssd1 vssd1 vccd1 vccd1 _19846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19777_ _19939_/CLK _19777_/D vssd1 vssd1 vccd1 vccd1 _19777_/Q sky130_fd_sc_hd__dfxtp_1
X_16989_ _16989_/A vssd1 vssd1 vccd1 vccd1 _19451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09530_ _09530_/A vssd1 vssd1 vccd1 vccd1 _19485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18728_ _18731_/CLK _18728_/D vssd1 vssd1 vccd1 vccd1 _18728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09461_ _12003_/A _14761_/C _09514_/B vssd1 vssd1 vccd1 vccd1 _12055_/B sky130_fd_sc_hd__or3_2
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18659_ _18660_/CLK _18659_/D vssd1 vssd1 vccd1 vccd1 _18659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09392_ _09406_/C _11699_/A _09394_/A _11783_/C vssd1 vssd1 vccd1 vccd1 _11707_/A
+ sky130_fd_sc_hd__nor4b_1
XANTENNA__12958__A1 _12875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10418__C1 _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__S1 _11086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17346__A0 _17189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11750__B _13910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12862__A _12863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13383__A1 _13223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10736__A3 _10734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10382__A _10382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13686__A2 _13685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18074__A1 _13612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11241__S0 _11156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11449__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ _10573_/S vssd1 vssd1 vccd1 vccd1 _09729_/A sky130_fd_sc_hd__buf_2
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11544__S1 _09660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09659_ _19382_/Q _19717_/Q _09659_/S vssd1 vssd1 vccd1 vccd1 _09660_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__A3 _15474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17104__S _17113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12670_ _12670_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _15482_/A sky130_fd_sc_hd__xnor2_4
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09411__A _18711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12949__A1 _18456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11621_/A _11621_/B vssd1 vssd1 vccd1 vccd1 _11622_/D sky130_fd_sc_hd__nand2_1
XANTENNA__12949__B2 _14350_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10557__A _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14340_ _14413_/A _14364_/A vssd1 vssd1 vccd1 vccd1 _14340_/Y sky130_fd_sc_hd__nor2_1
X_11552_ _18864_/Q _09540_/X _11541_/X _11551_/X vssd1 vssd1 vccd1 vccd1 _15982_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10503_ _19931_/Q _19545_/Q _19995_/Q _19114_/Q _10125_/S _10497_/X vssd1 vssd1 vccd1
+ vccd1 _10504_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11483_ _11477_/A _11482_/X _10719_/X vssd1 vssd1 vccd1 vccd1 _11483_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14271_ _14280_/A _14275_/D _14270_/Y vssd1 vssd1 vccd1 vccd1 _18657_/D sky130_fd_sc_hd__o21a_1
XFILLER_109_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ _16010_/A vssd1 vssd1 vccd1 vccd1 _19035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10434_ _10434_/A _10434_/B vssd1 vssd1 vccd1 vccd1 _10434_/Y sky130_fd_sc_hd__nor2_1
X_13222_ _13222_/A vssd1 vssd1 vccd1 vccd1 _18439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09673__S0 _09855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17774__S _17782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10365_ _10365_/A _10365_/B vssd1 vssd1 vccd1 vccd1 _10365_/X sky130_fd_sc_hd__or2_1
X_13153_ _13226_/A _18845_/Q vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__or2_1
XFILLER_88_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12104_ _18761_/Q _16069_/A vssd1 vssd1 vccd1 vccd1 _12107_/A sky130_fd_sc_hd__or2b_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17961_ _19849_/Q _17001_/X _17965_/S vssd1 vssd1 vccd1 vccd1 _17962_/A sky130_fd_sc_hd__mux2_1
X_13084_ _13956_/B _13070_/X _13077_/X _13079_/X _13083_/X vssd1 vssd1 vccd1 vccd1
+ _13570_/B sky130_fd_sc_hd__a2111o_2
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10296_ _10292_/A _10295_/X _09780_/A vssd1 vssd1 vccd1 vccd1 _10296_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_111_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output158_A _12656_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19700_ _19764_/CLK _19700_/D vssd1 vssd1 vccd1 vccd1 _19700_/Q sky130_fd_sc_hd__dfxtp_1
X_16912_ _16390_/X _19417_/Q _16914_/S vssd1 vssd1 vccd1 vccd1 _16913_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12035_ _12085_/A _12826_/B vssd1 vssd1 vccd1 vccd1 _12035_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17075__A _17075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12885__B1 _12881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17892_ _17892_/A vssd1 vssd1 vccd1 vccd1 _19818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19631_ _19985_/CLK _19631_/D vssd1 vssd1 vccd1 vccd1 _19631_/Q sky130_fd_sc_hd__dfxtp_1
X_16843_ _17203_/A _16843_/B vssd1 vssd1 vccd1 vccd1 _19387_/D sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_124_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19562_ _19562_/CLK _19562_/D vssd1 vssd1 vccd1 vccd1 _19562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16774_ _16774_/A vssd1 vssd1 vccd1 vccd1 _19355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13986_ _18569_/Q _13984_/B _13985_/Y vssd1 vssd1 vccd1 vccd1 _18569_/D sky130_fd_sc_hd__o21a_1
XFILLER_19_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18513_ _19972_/CLK _18513_/D vssd1 vssd1 vccd1 vccd1 _18513_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15725_ _12003_/A _15720_/X _15724_/Y _15713_/X vssd1 vssd1 vccd1 vccd1 _18936_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19493_ _20012_/CLK _19493_/D vssd1 vssd1 vccd1 vccd1 _19493_/Q sky130_fd_sc_hd__dfxtp_1
X_12937_ _12874_/X _12935_/X _12936_/X input12/X _12906_/X vssd1 vssd1 vccd1 vccd1
+ _16998_/A sky130_fd_sc_hd__a32o_4
XANTENNA__17576__A0 _17115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18444_ _19581_/CLK _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15656_ _15656_/A vssd1 vssd1 vccd1 vccd1 _18906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12868_ _14865_/A vssd1 vssd1 vccd1 vccd1 _14938_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14607_ _14607_/A vssd1 vssd1 vccd1 vccd1 _18770_/D sky130_fd_sc_hd__clkbuf_1
X_18375_ _18375_/A vssd1 vssd1 vccd1 vccd1 _20018_/D sky130_fd_sc_hd__clkbuf_1
X_11819_ _11819_/A vssd1 vssd1 vccd1 vccd1 _12881_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16853__S _16859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15587_ _13603_/A _18908_/Q _15589_/S vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__mux2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12799_ _12799_/A _12799_/B vssd1 vssd1 vccd1 vccd1 _12799_/Y sky130_fd_sc_hd__nand2_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17326_ _17160_/X _19578_/Q _17326_/S vssd1 vssd1 vccd1 vccd1 _17327_/A sky130_fd_sc_hd__mux2_1
X_14538_ input67/X _14544_/B vssd1 vssd1 vccd1 vccd1 _14538_/X sky130_fd_sc_hd__or2_1
XANTENNA__11612__A1 _11462_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17257_ _17163_/X _19547_/Q _17265_/S vssd1 vssd1 vccd1 vccd1 _17258_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13778__A _17014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14469_ _14468_/A _14468_/C _18722_/Q vssd1 vssd1 vccd1 vccd1 _14470_/C sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_49_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16208_ _16208_/A vssd1 vssd1 vccd1 vccd1 _16217_/S sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_170_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _18994_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17188_ _17188_/A vssd1 vssd1 vccd1 vccd1 _19517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16139_ _16139_/A vssd1 vssd1 vccd1 vccd1 _19090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11471__S0 _10821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_185_clock clkbuf_opt_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _18967_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14402__A _14413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19829_ _19829_/CLK _19829_/D vssd1 vssd1 vccd1 vccd1 _19829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09513_ _12003_/C _12004_/A _12004_/B _09514_/D vssd1 vssd1 vccd1 vccd1 _09513_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__17567__A0 _17103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10103__A1 _09884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12857__A _12857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _09444_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _15786_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_123_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19055_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12576__B _18539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17859__S _17865_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09375_ _18952_/Q _18951_/Q vssd1 vssd1 vccd1 vccd1 _11777_/B sky130_fd_sc_hd__or2b_1
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12800__B1 _12234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14791__B _15740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_138_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18731_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_165_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12159__A2 _12556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13108__A1 _13577_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ _10376_/A vssd1 vssd1 vccd1 vccd1 _10335_/A sky130_fd_sc_hd__buf_2
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _15968_/B vssd1 vssd1 vccd1 vccd1 _10104_/A sky130_fd_sc_hd__inv_2
XFILLER_0_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10840__A _18844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16003__S _16009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12331__A2 _12298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14608__A1 _13621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16938__S _16942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13840_ _18511_/Q _13838_/X _13852_/S vssd1 vssd1 vccd1 vccd1 _13841_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13771_ _17007_/A vssd1 vssd1 vccd1 vccd1 _13771_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13292__B1 _12984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10983_ _10996_/A vssd1 vssd1 vccd1 vccd1 _10983_/X sky130_fd_sc_hd__buf_4
XANTENNA__11671__A _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15510_ _15159_/X _15505_/Y _15509_/Y vssd1 vssd1 vccd1 vccd1 _15511_/C sky130_fd_sc_hd__a21oi_1
XFILLER_128_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12722_ _18481_/Q _12722_/B vssd1 vssd1 vccd1 vccd1 _12722_/X sky130_fd_sc_hd__or2_1
X_16490_ _16490_/A vssd1 vssd1 vccd1 vccd1 _19229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17769__S _17771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15441_ _15405_/X _15439_/X _15440_/X _14826_/A _12574_/X vssd1 vssd1 vccd1 vccd1
+ _15441_/X sky130_fd_sc_hd__a32o_1
X_12653_ _12679_/B _12679_/C vssd1 vssd1 vccd1 vccd1 _12653_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18160_ _18206_/S vssd1 vssd1 vccd1 vccd1 _18169_/S sky130_fd_sc_hd__clkbuf_4
X_11604_ _11604_/A _11604_/B vssd1 vssd1 vccd1 vccd1 _11605_/B sky130_fd_sc_hd__nand2_1
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15372_ _15366_/X _15367_/Y _15371_/X _15353_/X vssd1 vssd1 vccd1 vccd1 _15375_/B
+ sky130_fd_sc_hd__a211o_1
X_12584_ _12530_/X _12581_/Y _12628_/C _12583_/X vssd1 vssd1 vccd1 vccd1 _12584_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_129_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17111_ _17111_/A vssd1 vssd1 vccd1 vccd1 _19493_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10802__C1 _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14323_ _14407_/A vssd1 vssd1 vccd1 vccd1 _14356_/A sky130_fd_sc_hd__clkbuf_2
X_11535_ _09639_/X _11534_/X _11543_/A vssd1 vssd1 vccd1 vccd1 _11535_/Y sky130_fd_sc_hd__a21oi_1
X_18091_ _18851_/Q _11764_/X _18101_/S vssd1 vssd1 vccd1 vccd1 _18091_/X sky130_fd_sc_hd__mux2_2
XANTENNA_clkbuf_leaf_50_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17042_ _17042_/A vssd1 vssd1 vccd1 vccd1 _17042_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14254_ _14278_/B _14250_/B _18653_/Q vssd1 vssd1 vccd1 vccd1 _14257_/B sky130_fd_sc_hd__a21oi_1
X_11466_ _11477_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11466_/X sky130_fd_sc_hd__or2_1
XFILLER_139_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13205_ input7/X _13091_/A _13094_/A vssd1 vssd1 vccd1 vccd1 _13217_/A sky130_fd_sc_hd__a21o_1
X_10417_ _10458_/A _10416_/X _10192_/A vssd1 vssd1 vccd1 vccd1 _10417_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10256__S1 _09612_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14185_ _18634_/Q _14188_/C _14160_/X vssd1 vssd1 vccd1 vccd1 _14185_/Y sky130_fd_sc_hd__a21oi_1
X_11397_ _11181_/X _11392_/X _11396_/X _09816_/A vssd1 vssd1 vccd1 vccd1 _11397_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09971__B1 _09566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ _17026_/A vssd1 vssd1 vccd1 vccd1 _17668_/A sky130_fd_sc_hd__buf_2
XFILLER_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10348_ _10333_/X _10338_/X _09823_/A _10347_/X vssd1 vssd1 vccd1 vccd1 _10348_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_135_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18993_ _18993_/CLK input70/X vssd1 vssd1 vccd1 vccd1 _18993_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10279_ _10279_/A vssd1 vssd1 vccd1 vccd1 _10279_/X sky130_fd_sc_hd__clkbuf_4
X_17944_ _19842_/Q _17081_/X _17948_/S vssd1 vssd1 vccd1 vccd1 _17945_/A sky130_fd_sc_hd__mux2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13067_/A vssd1 vssd1 vccd1 vccd1 _18431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12018_ _18757_/Q _16075_/A vssd1 vssd1 vccd1 vccd1 _12059_/A sky130_fd_sc_hd__and2_1
X_17875_ _17875_/A vssd1 vssd1 vccd1 vccd1 _19811_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15786__C_N _15690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19614_ _19868_/CLK _19614_/D vssd1 vssd1 vccd1 vccd1 _19614_/Q sky130_fd_sc_hd__dfxtp_1
X_16826_ _16387_/X _19379_/Q _16830_/S vssd1 vssd1 vccd1 vccd1 _16827_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19545_ _19995_/CLK _19545_/D vssd1 vssd1 vccd1 vccd1 _19545_/Q sky130_fd_sc_hd__dfxtp_1
X_16757_ _16757_/A vssd1 vssd1 vccd1 vccd1 _19348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19764_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13969_ _14102_/A vssd1 vssd1 vccd1 vccd1 _13969_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15708_ _09481_/C _11865_/A _13700_/X _14529_/A vssd1 vssd1 vccd1 vccd1 _15708_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__15053__A _15978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11294__C1 _11015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19476_ _20030_/CLK _19476_/D vssd1 vssd1 vccd1 vccd1 _19476_/Q sky130_fd_sc_hd__dfxtp_1
X_16688_ _16688_/A vssd1 vssd1 vccd1 vccd1 _19318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_0_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__17679__S _17682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15988__A _16044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18427_ _20012_/CLK _18427_/D vssd1 vssd1 vccd1 vccd1 _18427_/Q sky130_fd_sc_hd__dfxtp_1
X_15639_ _15639_/A vssd1 vssd1 vccd1 vccd1 _18898_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16583__S _16591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19993_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__14783__B1 _14782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18358_ _18358_/A vssd1 vssd1 vccd1 vccd1 _20010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17309_ _17135_/X _19570_/Q _17315_/S vssd1 vssd1 vccd1 vccd1 _17310_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10495__S1 _10587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18289_ _17646_/X _19980_/Q _18291_/S vssd1 vssd1 vccd1 vccd1 _18290_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13301__A _17058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09962__B1 _09913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09993_ _19345_/Q _19616_/Q _19840_/Q _19584_/Q _09967_/X _09637_/A vssd1 vssd1 vccd1
+ vccd1 _09993_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16758__S _16758_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13274__B1 _11733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12587__A _12587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17589__S _17595_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09427_ _09423_/B _09415_/X _09420_/X _09426_/X vssd1 vssd1 vccd1 vccd1 _09443_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__16493__S _16497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ _13091_/A _09358_/B vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__and2_1
XFILLER_166_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15410__B _15410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09289_ _09289_/A _09289_/B _09289_/C _11931_/C vssd1 vssd1 vccd1 vccd1 _09292_/C
+ sky130_fd_sc_hd__or4b_1
XANTENNA__12526__S _12814_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14307__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11320_ _11320_/A _11320_/B vssd1 vssd1 vccd1 vccd1 _11320_/X sky130_fd_sc_hd__and2_1
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_clock clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_147_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11251_ _19918_/Q _19532_/Q _19982_/Q _19101_/Q _10977_/S _10983_/X vssd1 vssd1 vccd1
+ vccd1 _11252_/B sky130_fd_sc_hd__mux4_1
XFILLER_118_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18213__S _18219_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10202_ _10369_/A _10201_/X _09980_/A vssd1 vssd1 vccd1 vccd1 _10202_/X sky130_fd_sc_hd__o21a_1
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11182_ _11227_/A _11180_/X _11181_/X vssd1 vssd1 vccd1 vccd1 _11182_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11760__B1 _11759_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ _19347_/Q _19618_/Q _19842_/Q _19586_/Q _10449_/S _10185_/A vssd1 vssd1 vccd1
+ vccd1 _10133_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15990_ _12909_/X _19026_/Q _15998_/S vssd1 vssd1 vccd1 vccd1 _15991_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10064_ _10064_/A vssd1 vssd1 vccd1 vccd1 _10064_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input34_A io_ibus_inst[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14941_ _14941_/A vssd1 vssd1 vccd1 vccd1 _14941_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10315__A1 _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16668__S _16674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17660_ _17659_/X _19726_/Q _17666_/S vssd1 vssd1 vccd1 vccd1 _17661_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10410__S1 _10400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14872_ _15234_/B _15463_/B _14908_/S vssd1 vssd1 vccd1 vccd1 _14872_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16611_ _19284_/Q _13848_/X _16613_/S vssd1 vssd1 vccd1 vccd1 _16612_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13823_ _13839_/A vssd1 vssd1 vccd1 vccd1 _13836_/S sky130_fd_sc_hd__clkbuf_8
X_17591_ _17138_/X _19699_/Q _17595_/S vssd1 vssd1 vccd1 vccd1 _17592_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16542_ _16542_/A vssd1 vssd1 vccd1 vccd1 _19253_/D sky130_fd_sc_hd__clkbuf_1
X_19330_ _19957_/CLK _19330_/D vssd1 vssd1 vccd1 vccd1 _19330_/Q sky130_fd_sc_hd__dfxtp_1
X_13754_ _16992_/A vssd1 vssd1 vccd1 vccd1 _13754_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10966_ _09775_/A _10952_/X _10956_/X _10965_/X _11166_/A vssd1 vssd1 vccd1 vccd1
+ _10966_/X sky130_fd_sc_hd__a311o_1
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _12778_/A _12705_/B vssd1 vssd1 vccd1 vccd1 _12706_/A sky130_fd_sc_hd__or2_1
X_19261_ _19949_/CLK _19261_/D vssd1 vssd1 vccd1 vccd1 _19261_/Q sky130_fd_sc_hd__dfxtp_1
X_16473_ _16473_/A vssd1 vssd1 vccd1 vccd1 _19223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13685_ _13656_/X _13683_/X _13684_/Y _13660_/X _19016_/Q vssd1 vssd1 vccd1 vccd1
+ _13685_/X sky130_fd_sc_hd__a32o_2
X_10897_ _18434_/Q _19463_/Q _19500_/Q _19074_/Q _10787_/A _10856_/A vssd1 vssd1 vccd1
+ vccd1 _10897_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13820__S _13820_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18212_ _18212_/A vssd1 vssd1 vccd1 vccd1 _19945_/D sky130_fd_sc_hd__clkbuf_1
X_15424_ _15424_/A _15424_/B vssd1 vssd1 vccd1 vccd1 _15424_/Y sky130_fd_sc_hd__nor2_1
X_19192_ _19947_/CLK _19192_/D vssd1 vssd1 vccd1 vccd1 _19192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12636_ _12636_/A _15474_/A vssd1 vssd1 vccd1 vccd1 _12639_/A sky130_fd_sc_hd__xnor2_1
XFILLER_129_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09867__S0 _09598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18143_ _17643_/X _19915_/Q _18147_/S vssd1 vssd1 vccd1 vccd1 _18144_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12240__A1 _18906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15355_ _15355_/A _15355_/B vssd1 vssd1 vccd1 vccd1 _15355_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12567_ _09468_/A _12587_/A _12588_/A _12566_/Y vssd1 vssd1 vccd1 vccd1 _15436_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_79_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14306_ _18668_/Q _18667_/Q _18666_/Q _14306_/D vssd1 vssd1 vccd1 vccd1 _14317_/D
+ sky130_fd_sc_hd__and4_4
X_11518_ _11592_/A _11624_/A _11592_/C _10540_/A _11517_/X vssd1 vssd1 vccd1 vccd1
+ _11589_/C sky130_fd_sc_hd__a311o_2
X_18074_ _18846_/Q _13612_/X _18084_/S vssd1 vssd1 vccd1 vccd1 _18074_/X sky130_fd_sc_hd__mux2_1
X_15286_ _15286_/A vssd1 vssd1 vccd1 vccd1 _15286_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12498_ _12498_/A vssd1 vssd1 vccd1 vccd1 _12498_/Y sky130_fd_sc_hd__inv_6
XFILLER_156_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17025_ _17025_/A vssd1 vssd1 vccd1 vccd1 _19462_/D sky130_fd_sc_hd__clkbuf_1
X_14237_ _18647_/Q _18646_/Q vssd1 vssd1 vccd1 vccd1 _14242_/D sky130_fd_sc_hd__and2_1
X_11449_ _09772_/A _11440_/X _11444_/X _11448_/X _09816_/A vssd1 vssd1 vccd1 vccd1
+ _11449_/X sky130_fd_sc_hd__a311o_4
XANTENNA__11426__S0 _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09944__B1 _09809_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14168_ _18627_/Q _14166_/B _14167_/Y vssd1 vssd1 vccd1 vccd1 _18627_/D sky130_fd_sc_hd__o21a_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11576__A _15982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _18592_/Q vssd1 vssd1 vccd1 vccd1 _14051_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10480__A _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18976_ _19526_/CLK _18976_/D vssd1 vssd1 vccd1 vccd1 _18976_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _14099_/A vssd1 vssd1 vccd1 vccd1 _14105_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15493__A1 _18858_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17927_ _17927_/A vssd1 vssd1 vccd1 vccd1 _19834_/D sky130_fd_sc_hd__clkbuf_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16578__S _16580_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13791__A _13858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17858_ _17858_/A vssd1 vssd1 vccd1 vccd1 _19803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16809_ _16809_/A vssd1 vssd1 vccd1 vccd1 _19371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17789_ _17707_/X _19773_/Q _17793_/S vssd1 vssd1 vccd1 vccd1 _17790_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19528_ _19978_/CLK _19528_/D vssd1 vssd1 vccd1 vccd1 _19528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19459_ _19855_/CLK _19459_/D vssd1 vssd1 vccd1 vccd1 _19459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ input70/X vssd1 vssd1 vccd1 vccd1 _13926_/A sky130_fd_sc_hd__buf_2
XANTENNA__09858__S0 _11532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12854__B _12854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15230__B _15234_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14508__B1 _14507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17872__S _17876_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09976_ _10191_/A vssd1 vssd1 vccd1 vccd1 _10411_/A sky130_fd_sc_hd__buf_2
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13495__B1 _13490_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10820_ _10820_/A _10820_/B vssd1 vssd1 vccd1 vccd1 _10820_/Y sky130_fd_sc_hd__nand2_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09403__B _11869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10156__S0 _10141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10751_ _10690_/A _10750_/X _09759_/A vssd1 vssd1 vccd1 vccd1 _10751_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14747__B1 _15732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15421__A _15553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13470_ _18676_/Q _11889_/X _11852_/X _18644_/Q vssd1 vssd1 vccd1 vccd1 _13470_/X
+ sky130_fd_sc_hd__a22o_1
X_10682_ _10695_/A _10681_/X _10579_/X vssd1 vssd1 vccd1 vccd1 _10682_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ _12418_/X _12419_/Y _12420_/Y vssd1 vssd1 vccd1 vccd1 _12421_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10459__S1 _10400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16951__S _16953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10233__B1 _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15140_ _15082_/A _15138_/B _15081_/X _15139_/X vssd1 vssd1 vccd1 vccd1 _15140_/X
+ sky130_fd_sc_hd__o211a_1
X_12352_ _12340_/B _11997_/X _12346_/Y _12351_/X vssd1 vssd1 vccd1 vccd1 _12352_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11981__B1 _09911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13876__A _15715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ _11225_/A _11300_/X _11302_/X vssd1 vssd1 vccd1 vccd1 _11303_/Y sky130_fd_sc_hd__o21ai_1
X_15071_ _15365_/A vssd1 vssd1 vccd1 vccd1 _15071_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12283_ _12283_/A _12309_/C vssd1 vssd1 vccd1 vccd1 _12283_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14022_ _18582_/Q vssd1 vssd1 vccd1 vccd1 _14026_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11234_ _09773_/A _11225_/X _11227_/X _09803_/A _11233_/X vssd1 vssd1 vccd1 vccd1
+ _11234_/X sky130_fd_sc_hd__a311o_1
XFILLER_84_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10536__A1 _10382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17782__S _17782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18830_ _19880_/CLK _18830_/D vssd1 vssd1 vccd1 vccd1 _18830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ _11088_/A _11162_/X _11164_/X _11095_/X vssd1 vssd1 vccd1 vccd1 _11166_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16672__A0 _16374_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10116_ _19940_/Q _19554_/Q _20004_/Q _19123_/Q _09595_/A _10260_/A vssd1 vssd1 vccd1
+ vccd1 _10117_/B sky130_fd_sc_hd__mux4_1
XANTENNA_output140_A _12836_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18761_ _18762_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 _18761_/Q sky130_fd_sc_hd__dfxtp_1
X_11096_ _11242_/A _11094_/X _11095_/X vssd1 vssd1 vccd1 vccd1 _11096_/Y sky130_fd_sc_hd__o21ai_1
X_15973_ _19020_/Q _14803_/X _15972_/X vssd1 vssd1 vccd1 vccd1 _19020_/D sky130_fd_sc_hd__a21o_1
XFILLER_121_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17712_ _17712_/A vssd1 vssd1 vccd1 vccd1 _19742_/D sky130_fd_sc_hd__clkbuf_1
X_10047_ _15970_/C _12857_/B vssd1 vssd1 vccd1 vccd1 _10047_/Y sky130_fd_sc_hd__nand2_1
X_14924_ _15410_/B _15306_/B _14933_/S vssd1 vssd1 vccd1 vccd1 _14924_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18692_ _18693_/CLK _18692_/D vssd1 vssd1 vccd1 vccd1 _18692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17643_ _17643_/A vssd1 vssd1 vccd1 vccd1 _17643_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14855_ _14855_/A _14855_/B vssd1 vssd1 vccd1 vccd1 _14855_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13806_ _17042_/A vssd1 vssd1 vccd1 vccd1 _13806_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17811__A _17867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17574_ _17574_/A vssd1 vssd1 vccd1 vccd1 _19691_/D sky130_fd_sc_hd__clkbuf_1
X_14786_ _09188_/Y _14748_/X _14789_/B _18828_/Q vssd1 vssd1 vccd1 vccd1 _14787_/B
+ sky130_fd_sc_hd__a22o_1
X_11998_ _12503_/A vssd1 vssd1 vccd1 vccd1 _12448_/S sky130_fd_sc_hd__buf_2
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16525_ _16525_/A vssd1 vssd1 vccd1 vccd1 _19245_/D sky130_fd_sc_hd__clkbuf_1
X_19313_ _19873_/CLK _19313_/D vssd1 vssd1 vccd1 vccd1 _19313_/Q sky130_fd_sc_hd__dfxtp_1
X_13737_ _13737_/A _18895_/Q _13737_/C vssd1 vssd1 vccd1 vccd1 _13746_/B sky130_fd_sc_hd__or3_1
X_10949_ _10905_/A _10948_/X _09792_/A vssd1 vssd1 vccd1 vccd1 _10949_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16456_ _16456_/A vssd1 vssd1 vccd1 vccd1 _19215_/D sky130_fd_sc_hd__clkbuf_1
X_19244_ _19771_/CLK _19244_/D vssd1 vssd1 vccd1 vccd1 _19244_/Q sky130_fd_sc_hd__dfxtp_1
X_13668_ _18104_/A vssd1 vssd1 vccd1 vccd1 _18130_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15407_ _15539_/A _15410_/A vssd1 vssd1 vccd1 vccd1 _15407_/X sky130_fd_sc_hd__or2_1
X_19175_ _19960_/CLK _19175_/D vssd1 vssd1 vccd1 vccd1 _19175_/Q sky130_fd_sc_hd__dfxtp_1
X_12619_ _12619_/A _15449_/B vssd1 vssd1 vccd1 vccd1 _12619_/X sky130_fd_sc_hd__or2b_1
XANTENNA__17957__S _17965_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16387_ _17723_/A vssd1 vssd1 vccd1 vccd1 _16387_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13599_ _13603_/A _13603_/C vssd1 vssd1 vccd1 vccd1 _13599_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_129_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18126_ _18126_/A vssd1 vssd1 vccd1 vccd1 _19909_/D sky130_fd_sc_hd__clkbuf_1
X_15338_ _15338_/A _15338_/B vssd1 vssd1 vccd1 vccd1 _15338_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18057_ _18841_/Q _13572_/X _18067_/S vssd1 vssd1 vccd1 vccd1 _18057_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15269_ _15209_/X _15265_/Y _15267_/X _15268_/X vssd1 vssd1 vccd1 vccd1 _15272_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10870__S1 _10596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17008_ _19457_/Q _17007_/X _17008_/S vssd1 vssd1 vccd1 vccd1 _17009_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14910__A0 _15177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18101__A0 _18854_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17692__S _17698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09830_ _09830_/A vssd1 vssd1 vccd1 vccd1 _10690_/A sky130_fd_sc_hd__buf_2
XFILLER_140_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _10567_/A vssd1 vssd1 vccd1 vccd1 _10001_/A sky130_fd_sc_hd__buf_2
XFILLER_112_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18959_ _18960_/CLK _18959_/D vssd1 vssd1 vccd1 vccd1 _18959_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09692_ _09862_/A _09692_/B _09692_/C vssd1 vssd1 vccd1 vccd1 _09692_/X sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_172_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12849__B _12849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12865__A _12865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16771__S _16775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15941__A2 _15921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10766__A1 _09664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09959_ _09765_/A _09958_/X _09809_/A vssd1 vssd1 vccd1 vccd1 _09959_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17107__S _17113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ _18717_/Q _11776_/X _13245_/A vssd1 vssd1 vccd1 vccd1 _12970_/X sky130_fd_sc_hd__a21o_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10377__S0 _10209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _11961_/A _11919_/C _09246_/X _11932_/A _11920_/X vssd1 vssd1 vccd1 vccd1
+ _11921_/X sky130_fd_sc_hd__o311a_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14640_ _14646_/A _14640_/B vssd1 vssd1 vccd1 vccd1 _14641_/A sky130_fd_sc_hd__and2_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _12887_/A vssd1 vssd1 vccd1 vccd1 _11852_/X sky130_fd_sc_hd__buf_2
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10803_ _19667_/Q _19433_/Q _18498_/Q _19763_/Q _10787_/X _10788_/X vssd1 vssd1 vccd1
+ vccd1 _10804_/B sky130_fd_sc_hd__mux4_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _15833_/A _14571_/B vssd1 vssd1 vccd1 vccd1 _14572_/A sky130_fd_sc_hd__or2_1
XANTENNA__13640__A0 _18470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _15760_/A _11705_/A _11783_/C _15758_/A vssd1 vssd1 vccd1 vccd1 _13048_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16310_ _17646_/A vssd1 vssd1 vccd1 vccd1 _16310_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13522_ _19879_/Q vssd1 vssd1 vccd1 vccd1 _13523_/C sky130_fd_sc_hd__inv_2
XFILLER_159_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10734_ _09686_/A _10723_/Y _10729_/Y _10733_/Y _09874_/A vssd1 vssd1 vccd1 vccd1
+ _10734_/X sky130_fd_sc_hd__o311a_2
X_17290_ _17290_/A vssd1 vssd1 vccd1 vccd1 _19561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16241_ _13042_/X _19134_/Q _16247_/S vssd1 vssd1 vccd1 vccd1 _16242_/A sky130_fd_sc_hd__mux2_1
X_13453_ _18819_/Q _13071_/X _12984_/X _18786_/Q _13452_/X vssd1 vssd1 vccd1 vccd1
+ _13453_/X sky130_fd_sc_hd__a221o_1
X_10665_ _19143_/Q _19404_/Q _19303_/Q _19638_/Q _10724_/S _10820_/A vssd1 vssd1 vccd1
+ vccd1 _10666_/B sky130_fd_sc_hd__mux4_1
XANTENNA__16681__S _16685_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12404_ _09458_/A _12428_/A _12318_/Y vssd1 vssd1 vccd1 vccd1 _12404_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_167_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16172_ _16172_/A vssd1 vssd1 vccd1 vccd1 _19104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13384_ _17074_/A vssd1 vssd1 vccd1 vccd1 _17716_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10596_ _10596_/A vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__buf_2
XFILLER_126_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15123_ _15119_/X _15122_/X _15190_/S vssd1 vssd1 vccd1 vccd1 _15123_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17078__A _17078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12335_ _12335_/A vssd1 vssd1 vccd1 vccd1 _12335_/Y sky130_fd_sc_hd__inv_6
XFILLER_127_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19931_ _19995_/CLK _19931_/D vssd1 vssd1 vccd1 vccd1 _19931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15054_ _14949_/X _14935_/X _15121_/S vssd1 vssd1 vccd1 vccd1 _15054_/X sky130_fd_sc_hd__mux2_1
X_12266_ _15934_/B vssd1 vssd1 vccd1 vccd1 _12266_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14005_ _18576_/Q _14007_/C _14004_/Y vssd1 vssd1 vccd1 vccd1 _18576_/D sky130_fd_sc_hd__o21a_1
X_11217_ _20013_/Q _19851_/Q _19260_/Q _19030_/Q _11212_/X _11208_/X vssd1 vssd1 vccd1
+ vccd1 _11218_/B sky130_fd_sc_hd__mux4_1
X_19862_ _19976_/CLK _19862_/D vssd1 vssd1 vccd1 vccd1 _19862_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09308__B _12831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18401__S _18407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__A _18754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12197_ _18461_/Q _12372_/B vssd1 vssd1 vccd1 vccd1 _12197_/X sky130_fd_sc_hd__or2_1
XANTENNA__11182__A1 _11227_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput81 _12521_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[19] sky130_fd_sc_hd__buf_2
Xoutput92 _12766_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[29] sky130_fd_sc_hd__buf_2
XFILLER_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18813_ _19900_/CLK _18813_/D vssd1 vssd1 vccd1 vccd1 _18813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11148_ _20015_/Q _19853_/Q _19262_/Q _19032_/Q _11017_/A _11015_/X vssd1 vssd1 vccd1
+ vccd1 _11149_/B sky130_fd_sc_hd__mux4_1
X_19793_ _19856_/CLK _19793_/D vssd1 vssd1 vccd1 vccd1 _19793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11854__A _12876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18744_ _18744_/CLK _18744_/D vssd1 vssd1 vccd1 vccd1 _18744_/Q sky130_fd_sc_hd__dfxtp_1
X_15956_ _15964_/A _15956_/B vssd1 vssd1 vccd1 vccd1 _15956_/Y sky130_fd_sc_hd__nor2_2
X_11079_ _11070_/X _11078_/X _09682_/A vssd1 vssd1 vccd1 vccd1 _11079_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09324__A _18937_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ _14907_/A vssd1 vssd1 vccd1 vccd1 _15474_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__11485__A2 _11475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18675_ _18677_/CLK _18675_/D vssd1 vssd1 vccd1 vccd1 _18675_/Q sky130_fd_sc_hd__dfxtp_1
X_15887_ _09471_/C _15875_/X _15879_/X input54/X vssd1 vssd1 vccd1 vccd1 _15888_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17626_ _17189_/X _19715_/Q _17628_/S vssd1 vssd1 vccd1 vccd1 _17627_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14838_ _14948_/S _15004_/B vssd1 vssd1 vccd1 vccd1 _14993_/C sky130_fd_sc_hd__or2b_1
XFILLER_91_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17557_ _17557_/A vssd1 vssd1 vccd1 vccd1 _19684_/D sky130_fd_sc_hd__clkbuf_1
X_14769_ _14769_/A vssd1 vssd1 vccd1 vccd1 _18823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16508_ _19238_/Q _13803_/X _16508_/S vssd1 vssd1 vccd1 vccd1 _16509_/A sky130_fd_sc_hd__mux2_1
X_17488_ _17186_/X _19650_/Q _17492_/S vssd1 vssd1 vccd1 vccd1 _17489_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10917__B _12837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19227_ _19948_/CLK _19227_/D vssd1 vssd1 vccd1 vccd1 _19227_/Q sky130_fd_sc_hd__dfxtp_1
X_16439_ _16439_/A vssd1 vssd1 vccd1 vccd1 _19207_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16591__S _16591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_119_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19158_ _19622_/CLK _19158_/D vssd1 vssd1 vccd1 vccd1 _19158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18109_ _18108_/X _19904_/Q _18112_/S vssd1 vssd1 vccd1 vccd1 _18110_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19089_ _20033_/CLK _19089_/D vssd1 vssd1 vccd1 vccd1 _19089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10652__B _12847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18311__S _18313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20002_ _20002_/CLK _20002_/D vssd1 vssd1 vccd1 vccd1 _20002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12370__B1 _12364_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09813_ _19158_/Q _19419_/Q _19318_/Q _19653_/Q _09898_/S _09895_/A vssd1 vssd1 vccd1
+ vccd1 _09814_/B sky130_fd_sc_hd__mux4_1
XFILLER_115_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09744_ _10473_/A vssd1 vssd1 vccd1 vccd1 _09745_/A sky130_fd_sc_hd__buf_2
XFILLER_101_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10359__S0 _10356_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09234__A _18990_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09675_ _09660_/X _09669_/X _09673_/X _11547_/A _09568_/A vssd1 vssd1 vccd1 vccd1
+ _09692_/B sky130_fd_sc_hd__o221a_1
XFILLER_54_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10436__B1 _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18282__A _18350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10450_ _10109_/X _10449_/X _10112_/A vssd1 vssd1 vccd1 vccd1 _10450_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11087__S1 _11296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15127__A0 _18836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _19213_/Q _19804_/Q _19966_/Q _19181_/Q _10469_/S _10163_/X vssd1 vssd1 vccd1
+ vccd1 _10381_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10843__A _10843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12120_ _12121_/A _14912_/A vssd1 vssd1 vccd1 vccd1 _12120_/X sky130_fd_sc_hd__and2_1
XFILLER_123_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13689__A0 _11879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09357__A1 _09425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ _18520_/Q _18521_/Q _15633_/D vssd1 vssd1 vccd1 vccd1 _12128_/C sky130_fd_sc_hd__and3_1
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10598__S0 _10724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ _18432_/Q _19461_/Q _19498_/Q _19072_/Q _10995_/X _10996_/X vssd1 vssd1 vccd1
+ vccd1 _11002_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10372__C1 _09876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11674__A _15719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15810_ _15813_/A _15810_/B vssd1 vssd1 vccd1 vccd1 _15811_/A sky130_fd_sc_hd__and2_1
XANTENNA__15146__A _15458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16790_ _16790_/A vssd1 vssd1 vccd1 vccd1 _19362_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14050__A _14094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15850__A1 _11982_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15741_ _18942_/Q _15738_/B _15740_/Y _15730_/X vssd1 vssd1 vccd1 vccd1 _18942_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15850__B2 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _18584_/Q _11732_/X _12887_/X _14133_/B vssd1 vssd1 vccd1 vccd1 _12953_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11904_ _11904_/A vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__buf_4
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ _19885_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_1
X_15672_ _15672_/A vssd1 vssd1 vccd1 vccd1 _18913_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _19881_/Q _13431_/B vssd1 vssd1 vccd1 vccd1 _12884_/X sky130_fd_sc_hd__and2_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17411_ _17411_/A vssd1 vssd1 vccd1 vccd1 _17420_/S sky130_fd_sc_hd__buf_4
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14623_ _14629_/A _14623_/B vssd1 vssd1 vccd1 vccd1 _14624_/A sky130_fd_sc_hd__and2_1
X_18391_ _18391_/A vssd1 vssd1 vccd1 vccd1 _20025_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _15633_/A vssd1 vssd1 vccd1 vccd1 _11915_/B sky130_fd_sc_hd__buf_2
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output103_A _09188_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _17183_/X _19585_/Q _17348_/S vssd1 vssd1 vccd1 vccd1 _17343_/A sky130_fd_sc_hd__mux2_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _13531_/A _18994_/Q _09341_/X _14553_/X vssd1 vssd1 vccd1 vccd1 _14554_/X
+ sky130_fd_sc_hd__a31o_4
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _11728_/C _11764_/X _11765_/X vssd1 vssd1 vccd1 vccd1 _18747_/D sky130_fd_sc_hd__a21o_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _18996_/Q _13505_/B vssd1 vssd1 vccd1 vccd1 _13505_/X sky130_fd_sc_hd__or2_1
X_10717_ _10936_/A vssd1 vssd1 vccd1 vccd1 _11477_/A sky130_fd_sc_hd__clkbuf_2
X_17273_ _17273_/A vssd1 vssd1 vccd1 vccd1 _19554_/D sky130_fd_sc_hd__clkbuf_1
X_14485_ _14485_/A _18728_/Q _14485_/C vssd1 vssd1 vccd1 vccd1 _14487_/B sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_120_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11697_ _11697_/A _11697_/B _11697_/C _15775_/A vssd1 vssd1 vccd1 vccd1 _11712_/B
+ sky130_fd_sc_hd__or4b_4
XANTENNA__16705__A _16762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16224_ _16691_/A _16691_/B _16298_/C vssd1 vssd1 vccd1 vccd1 _17426_/B sky130_fd_sc_hd__or3_1
X_19012_ _19973_/CLK _19012_/D vssd1 vssd1 vccd1 vccd1 _19012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13436_ _18742_/Q vssd1 vssd1 vccd1 vccd1 _14526_/B sky130_fd_sc_hd__clkbuf_1
X_10648_ _10579_/X _10641_/Y _10643_/Y _10647_/Y _09805_/A vssd1 vssd1 vccd1 vccd1
+ _10648_/X sky130_fd_sc_hd__o311a_1
XFILLER_127_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11078__S1 _11077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16155_ _16155_/A vssd1 vssd1 vccd1 vccd1 _19096_/D sky130_fd_sc_hd__clkbuf_1
X_13367_ _13367_/A vssd1 vssd1 vccd1 vccd1 _18448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10579_ _10579_/A vssd1 vssd1 vccd1 vccd1 _10579_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15669__A1 _12416_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15106_ _15099_/X _15107_/B _15104_/X _15105_/X vssd1 vssd1 vccd1 vccd1 _15106_/X
+ sky130_fd_sc_hd__a211o_1
X_12318_ _12658_/A _12318_/B vssd1 vssd1 vccd1 vccd1 _12318_/Y sky130_fd_sc_hd__nand2_4
X_16086_ _16086_/A vssd1 vssd1 vccd1 vccd1 _19066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13298_ _13068_/X _13296_/X _13460_/A vssd1 vssd1 vccd1 vccd1 _13298_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19914_ _19978_/CLK _19914_/D vssd1 vssd1 vccd1 vccd1 _19914_/Q sky130_fd_sc_hd__dfxtp_1
X_15037_ _14915_/X _14897_/X _15039_/S vssd1 vssd1 vccd1 vccd1 _15037_/X sky130_fd_sc_hd__mux2_1
X_12249_ _12277_/B _12249_/B vssd1 vssd1 vccd1 vccd1 _12249_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19845_ _19975_/CLK _19845_/D vssd1 vssd1 vccd1 vccd1 _19845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10363__C1 _09555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17970__S _17976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19776_ _19971_/CLK _19776_/D vssd1 vssd1 vccd1 vccd1 _19776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16988_ _16396_/X _19451_/Q _16990_/S vssd1 vssd1 vccd1 vccd1 _16989_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18727_ _18741_/CLK _18727_/D vssd1 vssd1 vccd1 vccd1 _18727_/Q sky130_fd_sc_hd__dfxtp_1
X_15939_ _19006_/Q _15921_/X _15938_/X vssd1 vssd1 vccd1 vccd1 _19006_/D sky130_fd_sc_hd__a21o_1
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09460_ _14756_/B _12004_/B vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__or2_1
X_18658_ _18660_/CLK _18658_/D vssd1 vssd1 vccd1 vccd1 _18658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17609_ _17163_/X _19707_/Q _17617_/S vssd1 vssd1 vccd1 vccd1 _17610_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09391_ _18950_/Q vssd1 vssd1 vccd1 vccd1 _09406_/C sky130_fd_sc_hd__inv_2
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09808__C1 _09807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18589_ _18724_/CLK _18589_/D vssd1 vssd1 vccd1 vccd1 _18589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12958__A2 _13505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12862__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15839__A1_N input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10663__A _10663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13974__A _13991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18041__S _18044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11241__S1 _11108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17880__S _17880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09727_ _10574_/S vssd1 vssd1 vccd1 vccd1 _10573_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09658_ _09918_/S vssd1 vssd1 vccd1 vccd1 _09659_/S sky130_fd_sc_hd__buf_4
XFILLER_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _10921_/S vssd1 vssd1 vccd1 vccd1 _11468_/S sky130_fd_sc_hd__buf_2
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11617_/B _11617_/C _11617_/A vssd1 vssd1 vccd1 vccd1 _11621_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12949__A2 _12943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11082__B1 _09537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11551_ _09862_/A _11550_/X _09547_/X vssd1 vssd1 vccd1 vccd1 _11551_/X sky130_fd_sc_hd__a21o_1
XFILLER_156_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17120__S _17129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10502_ _10502_/A _10502_/B _10502_/C vssd1 vssd1 vccd1 vccd1 _10502_/Y sky130_fd_sc_hd__nor3_1
XFILLER_11_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14270_ _14288_/A _14270_/B vssd1 vssd1 vccd1 vccd1 _14270_/Y sky130_fd_sc_hd__nor2_1
X_11482_ _20022_/Q _19860_/Q _19269_/Q _19039_/Q _10708_/X _10710_/X vssd1 vssd1 vccd1
+ vccd1 _11482_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13221_ _13219_/X _18439_/Q _13284_/S vssd1 vssd1 vccd1 vccd1 _13222_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10433_ _19933_/Q _19547_/Q _19997_/Q _19116_/Q _10328_/S _10027_/A vssd1 vssd1 vccd1
+ vccd1 _10434_/B sky130_fd_sc_hd__mux4_1
XFILLER_155_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13374__A2 _12943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09673__S1 _09642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input64_A io_ibus_inst[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13152_ _13152_/A vssd1 vssd1 vccd1 vccd1 _18435_/D sky130_fd_sc_hd__clkbuf_1
X_10364_ _19934_/Q _19548_/Q _19998_/Q _19117_/Q _10356_/S _10261_/A vssd1 vssd1 vccd1
+ vccd1 _10365_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12103_ _09444_/A _16075_/A _12066_/B _12102_/X vssd1 vssd1 vccd1 vccd1 _16069_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_152_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17356__A _17424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13884__A _16836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17960_ _17960_/A vssd1 vssd1 vccd1 vccd1 _19848_/D sky130_fd_sc_hd__clkbuf_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _14279_/B _13081_/X _13082_/X _18722_/Q vssd1 vssd1 vccd1 vccd1 _13083_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10295_ _18447_/Q _19476_/Q _19513_/Q _19087_/Q _10037_/S _10329_/A vssd1 vssd1 vccd1
+ vccd1 _10295_/X sky130_fd_sc_hd__mux4_1
XANTENNA__16260__A _16282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16911_ _16911_/A vssd1 vssd1 vccd1 vccd1 _19416_/D sky130_fd_sc_hd__clkbuf_1
X_12034_ _18971_/Q _12033_/X _12084_/S vssd1 vssd1 vccd1 vccd1 _12034_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17891_ _19818_/Q _17004_/X _17893_/S vssd1 vssd1 vccd1 vccd1 _17892_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19630_ _19726_/CLK _19630_/D vssd1 vssd1 vccd1 vccd1 _19630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16842_ _16842_/A vssd1 vssd1 vccd1 vccd1 _19386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19561_ _19562_/CLK _19561_/D vssd1 vssd1 vccd1 vccd1 _19561_/Q sky130_fd_sc_hd__dfxtp_1
X_13985_ _14010_/A _13990_/C vssd1 vssd1 vccd1 vccd1 _13985_/Y sky130_fd_sc_hd__nor2_1
X_16773_ _16310_/X _19355_/Q _16775_/S vssd1 vssd1 vccd1 vccd1 _16774_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18512_ _19940_/CLK _18512_/D vssd1 vssd1 vccd1 vccd1 _18512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15724_ _16846_/B _15732_/B vssd1 vssd1 vccd1 vccd1 _15724_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12936_ _12936_/A _18866_/Q vssd1 vssd1 vccd1 vccd1 _12936_/X sky130_fd_sc_hd__or2_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ _20012_/CLK _19492_/D vssd1 vssd1 vccd1 vccd1 _19492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09602__A _11050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ _20028_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _12867_/A vssd1 vssd1 vccd1 vccd1 _12867_/X sky130_fd_sc_hd__clkbuf_1
X_15655_ _18906_/Q _12277_/B _15655_/S vssd1 vssd1 vccd1 vccd1 _15656_/A sky130_fd_sc_hd__mux2_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _12946_/A vssd1 vssd1 vccd1 vccd1 _13290_/B sky130_fd_sc_hd__clkbuf_2
X_14606_ _14612_/A _14606_/B vssd1 vssd1 vccd1 vccd1 _14607_/A sky130_fd_sc_hd__and2_1
X_18374_ _17665_/X _20018_/Q _18374_/S vssd1 vssd1 vccd1 vccd1 _18375_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15586_ _15586_/A vssd1 vssd1 vccd1 vccd1 _18875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12798_ _12799_/A _12799_/B vssd1 vssd1 vccd1 vccd1 _12798_/X sky130_fd_sc_hd__or2_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _17325_/A vssd1 vssd1 vccd1 vccd1 _19577_/D sky130_fd_sc_hd__clkbuf_1
X_14537_ _14537_/A vssd1 vssd1 vccd1 vccd1 _18751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11749_ _14665_/A vssd1 vssd1 vccd1 vccd1 _13910_/A sky130_fd_sc_hd__buf_2
X_17256_ _17267_/A vssd1 vssd1 vccd1 vccd1 _17265_/S sky130_fd_sc_hd__buf_4
XFILLER_147_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14468_ _14468_/A _18722_/Q _14468_/C vssd1 vssd1 vccd1 vccd1 _14470_/B sky130_fd_sc_hd__and3_1
XFILLER_88_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16207_ _16207_/A vssd1 vssd1 vccd1 vccd1 _19120_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14562__A1 _13531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17965__S _17965_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13419_ _13439_/A _13717_/B vssd1 vssd1 vccd1 vccd1 _13419_/Y sky130_fd_sc_hd__nand2_1
X_17187_ _17186_/X _19517_/Q _17193_/S vssd1 vssd1 vccd1 vccd1 _17188_/A sky130_fd_sc_hd__mux2_1
X_14399_ _14399_/A _14399_/B _14399_/C vssd1 vssd1 vccd1 vccd1 _18695_/D sky130_fd_sc_hd__nor3_1
X_16138_ _13406_/X _19090_/Q _16144_/S vssd1 vssd1 vccd1 vccd1 _16139_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13794__A _17030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16069_ _16069_/A _16069_/B vssd1 vssd1 vccd1 vccd1 _16069_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15201__A_N _12031_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19828_ _19828_/CLK _19828_/D vssd1 vssd1 vccd1 vccd1 _19828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19759_ _19985_/CLK _19759_/D vssd1 vssd1 vccd1 vccd1 _19759_/Q sky130_fd_sc_hd__dfxtp_1
X_09512_ _12003_/A _12003_/B _09482_/B vssd1 vssd1 vccd1 vccd1 _09514_/D sky130_fd_sc_hd__or3b_1
XFILLER_37_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12857__B _12857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _12064_/B _09443_/B vssd1 vssd1 vccd1 vccd1 _09444_/B sky130_fd_sc_hd__and2_1
XANTENNA__11761__B _13257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09374_ _18950_/Q vssd1 vssd1 vccd1 vccd1 _15760_/A sky130_fd_sc_hd__buf_2
XFILLER_40_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13969__A _14102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14564__S _14581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12800__A1 _12170_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16345__A _17681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16080__A _16148_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10080_ _09547_/X _10067_/X _10076_/X _10078_/X _10079_/Y vssd1 vssd1 vccd1 vccd1
+ _15968_/B sky130_fd_sc_hd__o32a_2
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10878__B1 _10719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13643__S _13689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13770_ _13770_/A vssd1 vssd1 vccd1 vccd1 _18489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10982_ _11258_/S _19232_/Q vssd1 vssd1 vccd1 vccd1 _10982_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12721_ _12717_/X _12720_/Y _12814_/S vssd1 vssd1 vccd1 vccd1 _12721_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15440_ _15478_/A _15440_/B vssd1 vssd1 vccd1 vccd1 _15440_/X sky130_fd_sc_hd__or2_1
X_12652_ _18781_/Q vssd1 vssd1 vccd1 vccd1 _12679_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_71_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11603_ _11601_/Y _11463_/Y _11602_/X vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__o21a_1
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15371_ _15368_/X _15373_/B _15369_/X _15370_/X vssd1 vssd1 vccd1 vccd1 _15371_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12583_ _12583_/A vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__buf_2
XFILLER_156_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12783__A _12783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11150__S0 _09721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14322_ _14327_/B _14327_/C _14321_/Y vssd1 vssd1 vccd1 vccd1 _18672_/D sky130_fd_sc_hd__o21a_1
X_17110_ _17109_/X _19493_/Q _17113_/S vssd1 vssd1 vccd1 vccd1 _17111_/A sky130_fd_sc_hd__mux2_1
X_11534_ _19383_/Q _19718_/Q _11534_/S vssd1 vssd1 vccd1 vccd1 _11534_/X sky130_fd_sc_hd__mux2_1
X_18090_ _18090_/A vssd1 vssd1 vccd1 vccd1 _19898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17785__S _17793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17041_ _17041_/A vssd1 vssd1 vccd1 vccd1 _19467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14253_ _14278_/B _14250_/B _14252_/Y vssd1 vssd1 vccd1 vccd1 _18652_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11465_ _19668_/Q _19434_/Q _18499_/Q _19764_/Q _10821_/S _10597_/A vssd1 vssd1 vccd1
+ vccd1 _11466_/B sky130_fd_sc_hd__mux4_1
XFILLER_171_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12555__A0 _12551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13204_ _13204_/A vssd1 vssd1 vccd1 vccd1 _18438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10416_ _20029_/Q _19867_/Q _19276_/Q _19046_/Q _10319_/X _10320_/X vssd1 vssd1 vccd1
+ vccd1 _10416_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14184_ _18633_/Q _14182_/B _14183_/Y vssd1 vssd1 vccd1 vccd1 _18633_/D sky130_fd_sc_hd__o21a_1
XANTENNA_output170_A _12173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11396_ _11435_/A _11393_/X _11395_/X _09788_/A vssd1 vssd1 vccd1 vccd1 _11396_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13135_ _09532_/X _13133_/X _13134_/X vssd1 vssd1 vccd1 vccd1 _17026_/A sky130_fd_sc_hd__o21a_4
X_10347_ _10162_/X _10340_/Y _10342_/Y _10344_/Y _10346_/Y vssd1 vssd1 vccd1 vccd1
+ _10347_/X sky130_fd_sc_hd__o32a_1
XFILLER_125_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ _18992_/CLK _18992_/D vssd1 vssd1 vccd1 vccd1 _18992_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14503__A _14528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17943_ _17943_/A vssd1 vssd1 vccd1 vccd1 _19841_/D sky130_fd_sc_hd__clkbuf_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13066_ _13065_/X _18431_/Q _13116_/S vssd1 vssd1 vccd1 vccd1 _13067_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10278_ _10278_/A _10278_/B vssd1 vssd1 vccd1 vccd1 _10278_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17246__A0 _17147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ _12062_/A vssd1 vssd1 vccd1 vccd1 _16075_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17874_ _19811_/Q _17084_/X _17876_/S vssd1 vssd1 vccd1 vccd1 _17875_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19613_ _19999_/CLK _19613_/D vssd1 vssd1 vccd1 vccd1 _19613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16825_ _16825_/A vssd1 vssd1 vccd1 vccd1 _19378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19544_ _20024_/CLK _19544_/D vssd1 vssd1 vccd1 vccd1 _19544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15334__A _15338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16756_ _19348_/Q _13848_/X _16758_/S vssd1 vssd1 vccd1 vccd1 _16757_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12086__A2 _09495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13968_ _18563_/Q _13966_/B _13967_/Y vssd1 vssd1 vccd1 vccd1 _18563_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10097__A1 _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15707_ _18929_/Q _15705_/X _15706_/X vssd1 vssd1 vccd1 vccd1 _18929_/D sky130_fd_sc_hd__a21o_1
X_19475_ _19999_/CLK _19475_/D vssd1 vssd1 vccd1 vccd1 _19475_/Q sky130_fd_sc_hd__dfxtp_1
X_12919_ _18352_/A _17738_/A _16846_/C vssd1 vssd1 vccd1 vccd1 _18352_/B sky130_fd_sc_hd__o21bai_1
XFILLER_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16687_ _16396_/X _19318_/Q _16689_/S vssd1 vssd1 vccd1 vccd1 _16688_/A sky130_fd_sc_hd__mux2_1
X_13899_ _12601_/A _13893_/X _12604_/Y _12607_/Y _13897_/X vssd1 vssd1 vccd1 vccd1
+ _18540_/D sky130_fd_sc_hd__o221a_1
XFILLER_94_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18426_ _19720_/CLK _18426_/D vssd1 vssd1 vccd1 vccd1 _18426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15638_ _18898_/Q _18519_/Q _15644_/S vssd1 vssd1 vccd1 vccd1 _15639_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14783__A1 _18827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18357_ _17640_/X _20010_/Q _18363_/S vssd1 vssd1 vccd1 vccd1 _18358_/A sky130_fd_sc_hd__mux2_1
X_15569_ _15602_/A vssd1 vssd1 vccd1 vccd1 _15578_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__12794__B1 _12154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17308_ _17308_/A vssd1 vssd1 vccd1 vccd1 _19569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18288_ _18288_/A vssd1 vssd1 vccd1 vccd1 _19979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17695__S _17698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17239_ _17138_/X _19539_/Q _17243_/S vssd1 vssd1 vccd1 vccd1 _17240_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09962__A1 _09884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09992_ _10057_/A _09985_/X _09991_/X vssd1 vssd1 vccd1 vccd1 _09992_/X sky130_fd_sc_hd__a21o_1
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14413__A _14413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09507__A _15139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17237__A0 _17135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15799__B1 _15798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12868__A _14865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__A _11772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11285__B1 _11003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11380__S0 _09586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09426_ _09414_/X _09422_/Y _12065_/B _12066_/B _18823_/Q vssd1 vssd1 vccd1 vccd1
+ _09426_/X sky130_fd_sc_hd__a2111o_1
XFILLER_80_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09357_ _09425_/B _09355_/A _09347_/X vssd1 vssd1 vccd1 vccd1 _09358_/B sky130_fd_sc_hd__a21o_1
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09288_ _09501_/B _09290_/B vssd1 vssd1 vccd1 vccd1 _11931_/C sky130_fd_sc_hd__or2_1
XANTENNA__14307__B _14317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_167_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11250_ _11257_/A _11250_/B vssd1 vssd1 vccd1 vccd1 _11250_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10201_ _19218_/Q _19809_/Q _19971_/Q _19186_/Q _10313_/S _09636_/A vssd1 vssd1 vccd1
+ vccd1 _10201_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09953__A1 _09833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11181_ _11181_/A vssd1 vssd1 vccd1 vccd1 _11181_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10851__A _10953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16014__S _16020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14323__A _14407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10132_ _10126_/X _10130_/X _10131_/X _10191_/A _10107_/A vssd1 vssd1 vccd1 vccd1
+ _10137_/B sky130_fd_sc_hd__o221a_1
XFILLER_122_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15138__B _15138_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16949__S _16953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11158__S _11158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10063_ _10270_/A _10063_/B vssd1 vssd1 vccd1 vccd1 _10063_/Y sky130_fd_sc_hd__nor2_1
X_14940_ _14932_/X _14939_/X _15016_/A vssd1 vssd1 vccd1 vccd1 _14941_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10946__S0 _10907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input27_A io_dbus_rdata[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ _14871_/A vssd1 vssd1 vccd1 vccd1 _15234_/B sky130_fd_sc_hd__buf_2
XFILLER_48_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16610_ _16610_/A vssd1 vssd1 vccd1 vccd1 _19283_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11682__A _11682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13822_ _17058_/A vssd1 vssd1 vccd1 vccd1 _13822_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17590_ _17590_/A vssd1 vssd1 vccd1 vccd1 _19698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16541_ _19253_/Q _13851_/X _16541_/S vssd1 vssd1 vccd1 vccd1 _16542_/A sky130_fd_sc_hd__mux2_1
X_13753_ _13753_/A vssd1 vssd1 vccd1 vccd1 _18485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10965_ _10900_/A _10957_/X _10964_/X _09792_/A vssd1 vssd1 vccd1 vccd1 _10965_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14993__A _14993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11371__S0 _11328_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12704_ _09263_/A _12657_/A _12860_/C _11945_/A vssd1 vssd1 vccd1 vccd1 _12705_/B
+ sky130_fd_sc_hd__a22o_1
X_19260_ _19324_/CLK _19260_/D vssd1 vssd1 vccd1 vccd1 _19260_/Q sky130_fd_sc_hd__dfxtp_1
X_16472_ _19223_/Q _13857_/X _16472_/S vssd1 vssd1 vccd1 vccd1 _16473_/A sky130_fd_sc_hd__mux2_1
X_13684_ _13732_/A _19016_/Q vssd1 vssd1 vccd1 vccd1 _13684_/Y sky130_fd_sc_hd__nand2_1
X_10896_ _11032_/A vssd1 vssd1 vccd1 vccd1 _10900_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18211_ _19945_/Q _17634_/A _18219_/S vssd1 vssd1 vccd1 vccd1 _18212_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_184_clock clkbuf_opt_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _18974_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12635_ _09466_/A _12657_/A _12682_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _15474_/A
+ sky130_fd_sc_hd__a211o_4
X_15423_ _15077_/X _15420_/Y _15422_/X _14855_/A vssd1 vssd1 vccd1 vccd1 _15423_/X
+ sky130_fd_sc_hd__a211o_1
X_19191_ _19846_/CLK _19191_/D vssd1 vssd1 vccd1 vccd1 _19191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09867__S1 _09851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13402__A _13439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18142_ _18142_/A vssd1 vssd1 vccd1 vccd1 _19914_/D sky130_fd_sc_hd__clkbuf_1
X_15354_ _15284_/X _15350_/Y _15352_/X _15353_/X vssd1 vssd1 vccd1 vccd1 _15357_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12566_ _12634_/A _12853_/B vssd1 vssd1 vccd1 vccd1 _12566_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11517_ _15958_/C _12850_/B vssd1 vssd1 vccd1 vccd1 _11517_/X sky130_fd_sc_hd__and2_1
X_14305_ _18667_/Q _14312_/C _14304_/Y vssd1 vssd1 vccd1 vccd1 _18667_/D sky130_fd_sc_hd__o21a_1
XFILLER_7_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18073_ _18073_/A vssd1 vssd1 vccd1 vccd1 _19893_/D sky130_fd_sc_hd__clkbuf_1
X_15285_ _15291_/A _15291_/B vssd1 vssd1 vccd1 vccd1 _15285_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12018__A _18757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12497_ _12497_/A _12497_/B vssd1 vssd1 vccd1 vccd1 _12498_/A sky130_fd_sc_hd__xnor2_4
XFILLER_156_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17024_ _19462_/Q _17023_/X _17024_/S vssd1 vssd1 vccd1 vccd1 _17025_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output95_A _12812_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14236_ _14236_/A _14236_/B vssd1 vssd1 vccd1 vccd1 _18647_/D sky130_fd_sc_hd__nor2_1
XFILLER_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11448_ _11401_/A _11445_/X _11447_/X _09788_/A vssd1 vssd1 vccd1 vccd1 _11448_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11426__S1 _11073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12960__B _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11857__A _19006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14167_ _14191_/A _14172_/C vssd1 vssd1 vccd1 vccd1 _14167_/Y sky130_fd_sc_hd__nor2_1
X_11379_ _11206_/A _11378_/X _09557_/A vssd1 vssd1 vccd1 vccd1 _11379_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13145_/A vssd1 vssd1 vccd1 vccd1 _13268_/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_122_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _19876_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11576__B _12866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18975_ _18975_/CLK _18975_/D vssd1 vssd1 vccd1 vccd1 _18975_/Q sky130_fd_sc_hd__dfxtp_1
X_14098_ _14245_/A vssd1 vssd1 vccd1 vccd1 _14146_/A sky130_fd_sc_hd__buf_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16859__S _16859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15493__A2 _15053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17926_ _19834_/Q _17055_/X _17926_/S vssd1 vssd1 vccd1 vccd1 _17927_/A sky130_fd_sc_hd__mux2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _18751_/Q _11778_/Y _11817_/A _18764_/Q _13048_/X vssd1 vssd1 vccd1 vccd1
+ _13053_/A sky130_fd_sc_hd__a221o_1
XFILLER_39_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10937__S0 _10703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17857_ _19803_/Q _17058_/X _17865_/S vssd1 vssd1 vccd1 vccd1 _17858_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16808_ _16361_/X _19371_/Q _16808_/S vssd1 vssd1 vccd1 vccd1 _16809_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_137_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _18741_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17788_ _17788_/A vssd1 vssd1 vccd1 vccd1 _19772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19527_ _20010_/CLK _19527_/D vssd1 vssd1 vccd1 vccd1 _19527_/Q sky130_fd_sc_hd__dfxtp_1
X_16739_ _19340_/Q _13822_/X _16747_/S vssd1 vssd1 vccd1 vccd1 _16740_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16594__S _16602_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09997__A _10200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10001__A _10001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13008__A1 _18459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19458_ _19950_/CLK _19458_/D vssd1 vssd1 vccd1 vccd1 _19458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09211_ _13473_/A vssd1 vssd1 vccd1 vccd1 _13439_/A sky130_fd_sc_hd__clkbuf_4
X_18409_ _18409_/A vssd1 vssd1 vccd1 vccd1 _18418_/S sky130_fd_sc_hd__buf_4
XFILLER_22_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19389_ _19389_/CLK _19389_/D vssd1 vssd1 vccd1 vccd1 _19389_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11114__S0 _09721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09858__S1 _09614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12767__B1 _18547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12870__B _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09935__A1 _09929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13192__B1 _11843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14143__A _14143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11742__B2 _18774_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09975_ _10553_/A vssd1 vssd1 vccd1 vccd1 _10191_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16769__S _16775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10950__C1 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_93_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14444__B1 _15807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10156__S1 _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750_ _19238_/Q _19733_/Q _10750_/S vssd1 vssd1 vccd1 vccd1 _10750_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ _11670_/A _11690_/A _13335_/B vssd1 vssd1 vccd1 vccd1 _09410_/D sky130_fd_sc_hd__nor3_1
XFILLER_13_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ _20024_/Q _19862_/Q _19271_/Q _19041_/Q _09726_/A _10010_/A vssd1 vssd1 vccd1
+ vccd1 _10681_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14747__B2 _12393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16009__S _16009_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12420_ _18469_/Q _12343_/X _12344_/X vssd1 vssd1 vccd1 vccd1 _12420_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10233__A1 _10438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ _12347_/X _12348_/X _12349_/Y _12350_/X vssd1 vssd1 vccd1 vccd1 _12351_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_166_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18224__S _18230_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11302_ _11311_/A _11301_/X _09789_/A vssd1 vssd1 vccd1 vccd1 _11302_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11981__A1 _09882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11981__B2 _12956_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15070_ _15151_/A vssd1 vssd1 vccd1 vccd1 _15365_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12282_ _18767_/Q vssd1 vssd1 vccd1 vccd1 _12283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14021_ _18581_/Q _14017_/B _14020_/Y vssd1 vssd1 vccd1 vccd1 _18581_/D sky130_fd_sc_hd__o21a_1
XANTENNA__09926__A1 _09933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11677__A _14672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ _09755_/A _11228_/X _11232_/X _11095_/A vssd1 vssd1 vccd1 vccd1 _11233_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14053__A _14088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__C1 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12930__B1 _11733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11164_/X sky130_fd_sc_hd__or2_1
XFILLER_45_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16679__S _16685_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10115_ _10191_/A vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18760_ _19063_/CLK _18760_/D vssd1 vssd1 vccd1 vccd1 _18760_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11095_ _11095_/A vssd1 vssd1 vccd1 vccd1 _11095_/X sky130_fd_sc_hd__clkbuf_2
X_15972_ _15978_/A _15978_/B _15972_/C vssd1 vssd1 vccd1 vccd1 _15972_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_54_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19767_/CLK sky130_fd_sc_hd__clkbuf_16
X_17711_ _17710_/X _19742_/Q _17714_/S vssd1 vssd1 vccd1 vccd1 _17712_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10046_ _09884_/X _10033_/X _10044_/X _09913_/X _10045_/Y vssd1 vssd1 vccd1 vccd1
+ _12857_/B sky130_fd_sc_hd__o32a_4
X_14923_ _15100_/A vssd1 vssd1 vccd1 vccd1 _14923_/X sky130_fd_sc_hd__clkbuf_2
X_18691_ _18693_/CLK _18691_/D vssd1 vssd1 vccd1 vccd1 _18691_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16424__A1 _13787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17642_ _17642_/A vssd1 vssd1 vccd1 vccd1 _19720_/D sky130_fd_sc_hd__clkbuf_1
X_14854_ _11971_/B _14852_/X _14854_/S vssd1 vssd1 vccd1 vccd1 _14855_/B sky130_fd_sc_hd__mux2_1
XFILLER_17_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13805_ _13805_/A vssd1 vssd1 vccd1 vccd1 _18500_/D sky130_fd_sc_hd__clkbuf_1
X_17573_ _17112_/X _19691_/Q _17573_/S vssd1 vssd1 vccd1 vccd1 _17574_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_69_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _20040_/CLK sky130_fd_sc_hd__clkbuf_16
X_14785_ _14785_/A vssd1 vssd1 vccd1 vccd1 _18827_/D sky130_fd_sc_hd__clkbuf_1
X_11997_ _12790_/A vssd1 vssd1 vccd1 vccd1 _11997_/X sky130_fd_sc_hd__buf_2
X_19312_ _20035_/CLK _19312_/D vssd1 vssd1 vccd1 vccd1 _19312_/Q sky130_fd_sc_hd__dfxtp_1
X_16524_ _19245_/Q _13826_/X _16530_/S vssd1 vssd1 vccd1 vccd1 _16525_/A sky130_fd_sc_hd__mux2_1
X_10948_ _20018_/Q _19856_/Q _19265_/Q _19035_/Q _10787_/A _10856_/A vssd1 vssd1 vccd1
+ vccd1 _10948_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13736_ _13736_/A vssd1 vssd1 vccd1 vccd1 _18483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19243_ _19771_/CLK _19243_/D vssd1 vssd1 vccd1 vccd1 _19243_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10472__A1 _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09610__A _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14738__A1 _13733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16455_ _19215_/Q _13832_/X _16457_/S vssd1 vssd1 vccd1 vccd1 _16456_/A sky130_fd_sc_hd__mux2_1
X_10879_ _10824_/A _10876_/X _10878_/X vssd1 vssd1 vccd1 vccd1 _10879_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13667_ _13587_/X _13665_/X _13666_/Y _13590_/X _19014_/Q vssd1 vssd1 vccd1 vccd1
+ _13667_/X sky130_fd_sc_hd__a32o_2
X_15406_ _15410_/A _15410_/B vssd1 vssd1 vccd1 vccd1 _15406_/Y sky130_fd_sc_hd__nand2_1
X_19174_ _19959_/CLK _19174_/D vssd1 vssd1 vccd1 vccd1 _19174_/Q sky130_fd_sc_hd__dfxtp_1
X_12618_ _12618_/A vssd1 vssd1 vccd1 vccd1 _15449_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_169_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16386_ _16386_/A vssd1 vssd1 vccd1 vccd1 _19186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13598_ _13598_/A vssd1 vssd1 vccd1 vccd1 _18464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18125_ _18124_/X _19909_/Q _18128_/S vssd1 vssd1 vccd1 vccd1 _18126_/A sky130_fd_sc_hd__mux2_1
X_15337_ _15284_/X _15334_/Y _15336_/X _15268_/X vssd1 vssd1 vccd1 vccd1 _15340_/B
+ sky130_fd_sc_hd__a211o_1
X_12549_ _12497_/A _12497_/B _12546_/Y _12548_/X vssd1 vssd1 vccd1 vccd1 _12550_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_157_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14662__S _14667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11783__A_N _15760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18056_ _18056_/A vssd1 vssd1 vccd1 vccd1 _19888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15268_ _15268_/A vssd1 vssd1 vccd1 vccd1 _15268_/X sky130_fd_sc_hd__clkbuf_2
X_17007_ _17007_/A vssd1 vssd1 vccd1 vccd1 _17007_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14219_ _18645_/Q _14216_/B _14218_/Y vssd1 vssd1 vccd1 vccd1 _18645_/D sky130_fd_sc_hd__o21a_1
XANTENNA__14910__A1 _12664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15199_ _15114_/X _15117_/X _15199_/S vssd1 vssd1 vccd1 vccd1 _15199_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18101__A1 _13677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11724__B2 _19010_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09393__A2 _11777_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16589__S _16591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09760_ _10680_/A vssd1 vssd1 vccd1 vccd1 _10567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18958_ _18958_/CLK _18958_/D vssd1 vssd1 vccd1 vccd1 _18958_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13477__A1 _12897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17909_ _19826_/Q _17030_/X _17915_/S vssd1 vssd1 vccd1 vccd1 _17910_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_115_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09691_ _11543_/A _09677_/X _09679_/X _09690_/X vssd1 vssd1 vccd1 vccd1 _09692_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18889_ _18924_/CLK _18889_/D vssd1 vssd1 vccd1 vccd1 _18889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13307__A _13307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_1_0_clock_A clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18309__S _18313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17213__S _17221_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17915__A1 _17039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10999__C1 _09873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10666__A _10832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13042__A _17656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13977__A _14010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18044__S _18044_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10074__S0 _09597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09958_ _19348_/Q _19619_/Q _19843_/Q _19587_/Q _09939_/X _09940_/X vssd1 vssd1 vccd1
+ vccd1 _09958_/X sky130_fd_sc_hd__mux4_2
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14601__A _14601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13468__A1 _18484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _09891_/A _09888_/X _09837_/X vssd1 vssd1 vccd1 vccd1 _09889_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10377__S1 _10163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _11961_/B _11920_/B _11920_/C _11920_/D vssd1 vssd1 vccd1 vccd1 _11920_/X
+ sky130_fd_sc_hd__or4_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _11851_/A vssd1 vssd1 vccd1 vccd1 _11851_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18219__S _18219_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _09776_/A _10790_/Y _10795_/Y _10801_/Y _09819_/A vssd1 vssd1 vccd1 vccd1
+ _10802_/X sky130_fd_sc_hd__o311a_1
XANTENNA__15432__A _15436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17123__S _17129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _18760_/Q _11801_/A _14601_/A vssd1 vssd1 vccd1 vccd1 _14571_/B sky130_fd_sc_hd__mux2_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11782_ _19062_/Q _12878_/A _12984_/A _18760_/Q vssd1 vssd1 vccd1 vccd1 _11782_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09844__B1 _09843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10733_ _10723_/A _10730_/X _10732_/X vssd1 vssd1 vccd1 vccd1 _10733_/Y sky130_fd_sc_hd__o21ai_1
X_13521_ _13690_/A vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16962__S _16964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ _18483_/Q _11755_/X _11847_/A _18707_/Q _13451_/X vssd1 vssd1 vccd1 vccd1
+ _13452_/X sky130_fd_sc_hd__a221o_1
X_16240_ _16240_/A vssd1 vssd1 vccd1 vccd1 _19133_/D sky130_fd_sc_hd__clkbuf_1
X_10664_ _10664_/A vssd1 vssd1 vccd1 vccd1 _10820_/A sky130_fd_sc_hd__buf_2
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14196__A2 _14197_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12403_ _11997_/X _12401_/Y _12402_/X vssd1 vssd1 vccd1 vccd1 _12403_/X sky130_fd_sc_hd__a21o_2
XFILLER_51_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13383_ _13223_/X _13369_/Y _13382_/X vssd1 vssd1 vccd1 vccd1 _17074_/A sky130_fd_sc_hd__o21ai_4
X_16171_ _13098_/X _19104_/Q _16173_/S vssd1 vssd1 vccd1 vccd1 _16172_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10595_ _10662_/A vssd1 vssd1 vccd1 vccd1 _10596_/A sky130_fd_sc_hd__buf_2
XFILLER_166_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12334_ _12334_/A _12334_/B vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__xnor2_4
X_15122_ _15040_/Y _15120_/Y _15121_/X _15082_/B vssd1 vssd1 vccd1 vccd1 _15122_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19930_ _19995_/CLK _19930_/D vssd1 vssd1 vccd1 vccd1 _19930_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17793__S _17793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15053_ _15978_/A vssd1 vssd1 vccd1 vccd1 _15053_/X sky130_fd_sc_hd__buf_4
X_12265_ _15270_/A _12265_/B vssd1 vssd1 vccd1 vccd1 _12299_/A sky130_fd_sc_hd__xnor2_4
X_14004_ _18576_/Q _14007_/C _13969_/X vssd1 vssd1 vccd1 vccd1 _14004_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10065__S0 _09597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11216_ _11070_/X _11215_/X _09559_/A vssd1 vssd1 vccd1 vccd1 _11216_/Y sky130_fd_sc_hd__o21ai_1
X_19861_ _19861_/CLK _19861_/D vssd1 vssd1 vccd1 vccd1 _19861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12196_ _12196_/A vssd1 vssd1 vccd1 vccd1 _12372_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10914__C1 _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput71 _12871_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_150_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput82 _11971_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[1] sky130_fd_sc_hd__buf_2
X_18812_ _19900_/CLK _18812_/D vssd1 vssd1 vccd1 vccd1 _18812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput93 _11994_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ _11088_/A _11146_/X _09773_/A vssd1 vssd1 vccd1 vccd1 _11147_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16202__S _16206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19792_ _19792_/CLK _19792_/D vssd1 vssd1 vccd1 vccd1 _19792_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13459__A1 _12956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09605__A _10048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18743_ _18744_/CLK _18743_/D vssd1 vssd1 vccd1 vccd1 _18743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15955_ _15955_/A vssd1 vssd1 vccd1 vccd1 _15955_/X sky130_fd_sc_hd__buf_2
X_11078_ _19199_/Q _19790_/Q _19952_/Q _19167_/Q _11121_/S _11077_/X vssd1 vssd1 vccd1
+ vccd1 _11078_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14230__B _14242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ _19938_/Q _19552_/Q _20002_/Q _19121_/Q _10095_/S _10028_/X vssd1 vssd1 vccd1
+ vccd1 _10030_/B sky130_fd_sc_hd__mux4_1
X_14906_ _14906_/A vssd1 vssd1 vccd1 vccd1 _15219_/B sky130_fd_sc_hd__clkbuf_4
X_18674_ _18688_/CLK _18674_/D vssd1 vssd1 vccd1 vccd1 _18674_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11485__A3 _11484_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15886_ _15886_/A vssd1 vssd1 vccd1 vccd1 _18988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17625_ _17625_/A vssd1 vssd1 vccd1 vccd1 _19714_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11890__B1 _11772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14837_ _14869_/A vssd1 vssd1 vccd1 vccd1 _14948_/S sky130_fd_sc_hd__buf_2
XFILLER_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12966__A _19487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17556_ _19684_/Q vssd1 vssd1 vccd1 vccd1 _17557_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_51_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09835__B1 _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14768_ _14780_/A _14768_/B vssd1 vssd1 vccd1 vccd1 _14769_/A sky130_fd_sc_hd__and2_1
XFILLER_60_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16507_ _16507_/A vssd1 vssd1 vccd1 vccd1 _19237_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15908__A0 _18996_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17968__S _17976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09930__S0 _09668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ _11813_/X _13717_/X _13718_/Y _11831_/X _19021_/Q vssd1 vssd1 vccd1 vccd1
+ _13719_/X sky130_fd_sc_hd__a32o_2
X_17487_ _17487_/A vssd1 vssd1 vccd1 vccd1 _19649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14699_ _18801_/Q _11833_/D _14705_/S vssd1 vssd1 vccd1 vccd1 _14700_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19226_ _19485_/CLK _19226_/D vssd1 vssd1 vccd1 vccd1 _19226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16438_ _19207_/Q _13806_/X _16446_/S vssd1 vssd1 vccd1 vccd1 _16439_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13797__A _17033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19157_ _20038_/CLK _19157_/D vssd1 vssd1 vccd1 vccd1 _19157_/Q sky130_fd_sc_hd__dfxtp_1
X_16369_ _16368_/X _19181_/Q _16378_/S vssd1 vssd1 vccd1 vccd1 _16370_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_41_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18108_ _18856_/Q _11879_/X _18118_/S vssd1 vssd1 vccd1 vccd1 _18108_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19088_ _20035_/CLK _19088_/D vssd1 vssd1 vccd1 vccd1 _19088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18039_ _18039_/A vssd1 vssd1 vccd1 vccd1 _19883_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10425__S _10470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20001_ _20032_/CLK _20001_/D vssd1 vssd1 vccd1 vccd1 _20001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09812_ _09891_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _09812_/X sky130_fd_sc_hd__or2_1
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14421__A _14479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__S0 _09733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ _10522_/A vssd1 vssd1 vccd1 vccd1 _10473_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09674_ _10069_/A vssd1 vssd1 vccd1 vccd1 _11547_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09234__B _18989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14567__S _14581_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12876__A _12876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__A _15758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11228__A3 _19165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10436__A1 _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17878__S _17880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16782__S _16786_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11936__A1 _15899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13500__A _17093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10295__S0 _10037_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ _10380_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10380_/X sky130_fd_sc_hd__or2_1
XFILLER_136_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09409__B _11690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18077__A0 _18847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12050_ _12050_/A vssd1 vssd1 vccd1 vccd1 _12791_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11001_ _11001_/A _11001_/B vssd1 vssd1 vccd1 vccd1 _11001_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10598__S1 _10654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15740_ _15740_/A _15740_/B vssd1 vssd1 vccd1 vccd1 _15740_/Y sky130_fd_sc_hd__nand2_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _18616_/Q vssd1 vssd1 vccd1 vccd1 _14133_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11903_ _11903_/A vssd1 vssd1 vccd1 vccd1 _11904_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11872__B1 _14555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15671_ _18913_/Q _12446_/A _15677_/S vssd1 vssd1 vccd1 vccd1 _15672_/A sky130_fd_sc_hd__mux2_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _13164_/B vssd1 vssd1 vccd1 vccd1 _13431_/B sky130_fd_sc_hd__buf_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17410_/A vssd1 vssd1 vccd1 vccd1 _19615_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11690__A _11690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _12508_/A _11764_/X _14632_/S vssd1 vssd1 vccd1 vccd1 _14623_/B sky130_fd_sc_hd__mux2_1
XFILLER_61_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18390_ _17688_/X _20025_/Q _18396_/S vssd1 vssd1 vccd1 vccd1 _18391_/A sky130_fd_sc_hd__mux2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _13926_/A vssd1 vssd1 vccd1 vccd1 _13879_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _17341_/A vssd1 vssd1 vccd1 vccd1 _19584_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _18747_/Q _13910_/A _14670_/S vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__and3_1
XFILLER_13_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14553_ _18994_/Q _12892_/X _14552_/Y _11717_/X vssd1 vssd1 vccd1 vccd1 _14553_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _10934_/A vssd1 vssd1 vccd1 vccd1 _10936_/A sky130_fd_sc_hd__clkbuf_2
X_13504_ _13504_/A _19879_/Q vssd1 vssd1 vccd1 vccd1 _13504_/Y sky130_fd_sc_hd__xnor2_1
X_17272_ _17186_/X _19554_/Q _17276_/S vssd1 vssd1 vccd1 vccd1 _17273_/A sky130_fd_sc_hd__mux2_1
X_11696_ _18694_/Q vssd1 vssd1 vccd1 vccd1 _14398_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14484_ _14485_/A _14485_/C _14483_/Y vssd1 vssd1 vccd1 vccd1 _18727_/D sky130_fd_sc_hd__o21a_1
X_19011_ _19023_/CLK _19011_/D vssd1 vssd1 vccd1 vccd1 _19011_/Q sky130_fd_sc_hd__dfxtp_1
X_16223_ _18352_/A _18352_/B vssd1 vssd1 vccd1 vccd1 _16692_/A sky130_fd_sc_hd__or2_2
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10647_ _10643_/A _10644_/X _10646_/X vssd1 vssd1 vccd1 vccd1 _10647_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ _14105_/B _11851_/X _12887_/X _18642_/Q vssd1 vssd1 vccd1 vccd1 _13435_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11927__A1 _15847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11927__B2 _09468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13366_ _13365_/X _18448_/Q _13366_/S vssd1 vssd1 vccd1 vccd1 _13367_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16154_ _12909_/X _19096_/Q _16162_/S vssd1 vssd1 vccd1 vccd1 _16155_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10578_ _19337_/Q _19608_/Q _19832_/Q _19576_/Q _10574_/S _10522_/A vssd1 vssd1 vccd1
+ vccd1 _10578_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13129__A0 _18843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14225__B _18938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__A2_N _09540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15105_ _15353_/A vssd1 vssd1 vccd1 vccd1 _15105_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12317_ _12317_/A _12588_/A vssd1 vssd1 vccd1 vccd1 _12318_/B sky130_fd_sc_hd__nand2_2
XANTENNA__14940__S _15016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16085_ _12963_/X _19066_/Q _16089_/S vssd1 vssd1 vccd1 vccd1 _16086_/A sky130_fd_sc_hd__mux2_1
X_13297_ _13297_/A vssd1 vssd1 vccd1 vccd1 _13460_/A sky130_fd_sc_hd__buf_2
XANTENNA__18412__S _18418_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__S0 _09657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19913_ _19978_/CLK _19913_/D vssd1 vssd1 vccd1 vccd1 _19913_/Q sky130_fd_sc_hd__dfxtp_1
X_12248_ _12277_/B _12303_/B vssd1 vssd1 vccd1 vccd1 _12258_/A sky130_fd_sc_hd__or2_1
X_15036_ _14910_/X _14913_/X _15039_/S vssd1 vssd1 vccd1 vccd1 _15036_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17028__S _17040_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19844_ _20039_/CLK _19844_/D vssd1 vssd1 vccd1 vccd1 _19844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12179_ _15925_/C _18904_/Q _12179_/S vssd1 vssd1 vccd1 vccd1 _14906_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09335__A _17098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19775_ _19839_/CLK _19775_/D vssd1 vssd1 vccd1 vccd1 _19775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16987_ _16987_/A vssd1 vssd1 vccd1 vccd1 _19450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18726_ _18741_/CLK _18726_/D vssd1 vssd1 vccd1 vccd1 _18726_/Q sky130_fd_sc_hd__dfxtp_1
X_15938_ _15940_/A _15955_/A _15938_/C vssd1 vssd1 vccd1 vccd1 _15938_/X sky130_fd_sc_hd__and3_1
XFILLER_36_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18657_ _18660_/CLK _18657_/D vssd1 vssd1 vccd1 vccd1 _18657_/Q sky130_fd_sc_hd__dfxtp_1
X_15869_ _15869_/A vssd1 vssd1 vccd1 vccd1 _18983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17608_ _17619_/A vssd1 vssd1 vccd1 vccd1 _17617_/S sky130_fd_sc_hd__buf_4
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09390_ _11869_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _11695_/A sky130_fd_sc_hd__or2_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18588_ _18655_/CLK _18588_/D vssd1 vssd1 vccd1 vccd1 _18588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17698__S _17698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17539_ _17539_/A vssd1 vssd1 vccd1 vccd1 _19675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15800__A _15813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11105__A _11158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19209_ _20027_/CLK _19209_/D vssd1 vssd1 vccd1 vccd1 _19209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16107__S _16111_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12040__A0 _11292_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18322__S _18324_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11775__A _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14151__A _14407_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A io_dbus_rdata[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09726_ _09726_/A vssd1 vssd1 vccd1 vccd1 _10574_/S sky130_fd_sc_hd__buf_2
XFILLER_41_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17034__A1 _17033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09657_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09918_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16793__A0 _16339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09588_ _10775_/A vssd1 vssd1 vccd1 vccd1 _10921_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18293__A _18350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17401__S _17409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11015__A _11015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11550_ _09568_/X _11543_/Y _11545_/Y _11547_/Y _11549_/Y vssd1 vssd1 vccd1 vccd1
+ _11550_/X sky130_fd_sc_hd__o32a_1
XFILLER_11_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11082__A1 _09848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11082__B2 _18840_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10501_ _10557_/A _10498_/X _10500_/X _09687_/A vssd1 vssd1 vccd1 vccd1 _10502_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ _11481_/A _11481_/B vssd1 vssd1 vccd1 vccd1 _11481_/X sky130_fd_sc_hd__or2_1
XANTENNA__10854__A _10854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ _13386_/A vssd1 vssd1 vccd1 vccd1 _13284_/S sky130_fd_sc_hd__buf_2
X_10432_ _10159_/X _10427_/X _10429_/Y _10431_/Y _09806_/A vssd1 vssd1 vccd1 vccd1
+ _10432_/X sky130_fd_sc_hd__o221a_1
XFILLER_164_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13151_ _13150_/X _18435_/Q _13203_/S vssd1 vssd1 vccd1 vccd1 _13152_/A sky130_fd_sc_hd__mux2_1
X_10363_ _09566_/A _10358_/X _10360_/X _10362_/X _09555_/A vssd1 vssd1 vccd1 vccd1
+ _10363_/X sky130_fd_sc_hd__a221o_2
XFILLER_12_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17637__A _17736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12102_ _18756_/Q _18789_/Q _12101_/Y _12064_/B vssd1 vssd1 vccd1 vccd1 _12102_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13082_ _13082_/A vssd1 vssd1 vccd1 vccd1 _13082_/X sky130_fd_sc_hd__buf_2
X_10294_ _10294_/A _10294_/B vssd1 vssd1 vccd1 vccd1 _10294_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_input57_A io_ibus_inst[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16910_ _16387_/X _19416_/Q _16914_/S vssd1 vssd1 vccd1 vccd1 _16911_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11685__A _14227_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12033_ _14749_/A _12032_/X _12033_/S vssd1 vssd1 vccd1 vccd1 _12033_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17890_ _17890_/A vssd1 vssd1 vccd1 vccd1 _19817_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16841_ _17201_/A _16841_/B vssd1 vssd1 vccd1 vccd1 _16842_/A sky130_fd_sc_hd__and2_1
XANTENNA__16687__S _16689_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19560_ _19656_/CLK _19560_/D vssd1 vssd1 vccd1 vccd1 _19560_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_9_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16772_ _16772_/A vssd1 vssd1 vccd1 vccd1 _19354_/D sky130_fd_sc_hd__clkbuf_1
X_13984_ _18569_/Q _13984_/B vssd1 vssd1 vccd1 vccd1 _13990_/C sky130_fd_sc_hd__and2_1
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18511_ _19873_/CLK _18511_/D vssd1 vssd1 vccd1 vccd1 _18511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15723_ _11925_/B _15720_/X _15722_/X _15713_/X vssd1 vssd1 vccd1 vccd1 _18935_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19491_ _20010_/CLK _19491_/D vssd1 vssd1 vccd1 vccd1 _19491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12935_ _12875_/X _12933_/X _12934_/Y _12897_/X vssd1 vssd1 vccd1 vccd1 _12935_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_92_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _19865_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13405__A _17078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _15654_/A vssd1 vssd1 vccd1 vccd1 _18905_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _12866_/A _12866_/B _12866_/C vssd1 vssd1 vccd1 vccd1 _12867_/A sky130_fd_sc_hd__and3_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _18770_/Q _13612_/X _14615_/S vssd1 vssd1 vccd1 vccd1 _14606_/B sky130_fd_sc_hd__mux2_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _18373_/A vssd1 vssd1 vccd1 vccd1 _20017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11817_ _11817_/A vssd1 vssd1 vccd1 vccd1 _11817_/X sky130_fd_sc_hd__clkbuf_2
X_15585_ _18875_/Q _18907_/Q _15589_/S vssd1 vssd1 vccd1 vccd1 _15586_/A sky130_fd_sc_hd__mux2_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18407__S _18407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16716__A _16762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12797_ _18787_/Q vssd1 vssd1 vccd1 vccd1 _12799_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17157_/X _19577_/Q _17326_/S vssd1 vssd1 vccd1 vccd1 _17325_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17311__S _17315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14536_ _14548_/A _18751_/Q _14670_/S vssd1 vssd1 vccd1 vccd1 _14537_/A sky130_fd_sc_hd__mux2_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _11731_/X _11746_/X _11747_/Y _11723_/X _19011_/Q vssd1 vssd1 vccd1 vccd1
+ _11748_/X sky130_fd_sc_hd__a32o_4
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17255_ _17255_/A vssd1 vssd1 vccd1 vccd1 _19546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14467_ _14468_/A _14468_/C _14466_/Y vssd1 vssd1 vccd1 vccd1 _18721_/D sky130_fd_sc_hd__o21a_1
X_11679_ _18598_/Q vssd1 vssd1 vccd1 vccd1 _14070_/B sky130_fd_sc_hd__clkbuf_2
X_16206_ _13365_/X _19120_/Q _16206_/S vssd1 vssd1 vccd1 vccd1 _16207_/A sky130_fd_sc_hd__mux2_1
X_13418_ _18577_/Q _13189_/X _13415_/X _13416_/X _13417_/X vssd1 vssd1 vccd1 vccd1
+ _13717_/B sky130_fd_sc_hd__a2111o_1
XFILLER_174_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17186_ _17723_/A vssd1 vssd1 vccd1 vccd1 _17186_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14562__A2 _18995_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14398_ _18695_/Q _14398_/B _14398_/C vssd1 vssd1 vccd1 vccd1 _14399_/C sky130_fd_sc_hd__and3_1
XANTENNA__10033__C1 _09823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16137_ _16137_/A vssd1 vssd1 vccd1 vccd1 _19089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13349_ _18856_/Q _11877_/B _13349_/S vssd1 vssd1 vccd1 vccd1 _13349_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10584__B1 _09913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16068_ _16068_/A vssd1 vssd1 vccd1 vccd1 _19060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17981__S _17987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15019_ _14929_/X _14878_/X _15023_/S vssd1 vssd1 vccd1 vccd1 _15019_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19827_ _19827_/CLK _19827_/D vssd1 vssd1 vccd1 vccd1 _19827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12089__A0 _11223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__A _10279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19758_ _19758_/CLK _19758_/D vssd1 vssd1 vccd1 vccd1 _19758_/Q sky130_fd_sc_hd__dfxtp_1
X_09511_ _11961_/B _09500_/B _14811_/C vssd1 vssd1 vccd1 vccd1 _14804_/D sky130_fd_sc_hd__o21bai_1
X_18709_ _19883_/CLK _18709_/D vssd1 vssd1 vccd1 vccd1 _18709_/Q sky130_fd_sc_hd__dfxtp_1
X_19689_ _20012_/CLK _19689_/D vssd1 vssd1 vccd1 vccd1 _19689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11534__S _11534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09442_ _09442_/A _09442_/B vssd1 vssd1 vccd1 vccd1 _15856_/A sky130_fd_sc_hd__or2_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _09407_/C vssd1 vssd1 vccd1 vccd1 _14227_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_40_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17221__S _17221_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10674__A _10674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14553__A2 _12892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12564__A1 _12554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13985__A _14010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17891__S _17893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10422__S0 _10388_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_163_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09709_ _10211_/A vssd1 vssd1 vccd1 vccd1 _10643_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11827__B1 _11823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10981_ _11270_/S vssd1 vssd1 vccd1 vccd1 _11258_/S sky130_fd_sc_hd__buf_4
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13292__A2 _13071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15870__A1_N input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12720_ _12720_/A _12768_/C vssd1 vssd1 vccd1 vccd1 _12720_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ _12522_/X _12649_/X _12650_/X vssd1 vssd1 vccd1 vccd1 _12651_/X sky130_fd_sc_hd__o21a_1
X_11602_ _11605_/A _11604_/A _11604_/B _10918_/A vssd1 vssd1 vccd1 vccd1 _11602_/X
+ sky130_fd_sc_hd__a31o_1
X_12582_ _18778_/Q _18777_/Q _12582_/C vssd1 vssd1 vccd1 vccd1 _12628_/C sky130_fd_sc_hd__and3_1
X_15370_ _15381_/A _15373_/A vssd1 vssd1 vccd1 vccd1 _15370_/X sky130_fd_sc_hd__or2_1
XFILLER_8_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10802__A1 _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14321_ _14327_/B _14327_/C _14203_/X vssd1 vssd1 vccd1 vccd1 _14321_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11150__S1 _10854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11533_ _11533_/A _11533_/B vssd1 vssd1 vccd1 vccd1 _11533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17040_ _19467_/Q _17039_/X _17040_/S vssd1 vssd1 vccd1 vccd1 _17041_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11464_ _11605_/A _11604_/A _11604_/B _10918_/A _11463_/Y vssd1 vssd1 vccd1 vccd1
+ _11617_/C sky130_fd_sc_hd__a311o_1
X_14252_ _14278_/B _14250_/B _14203_/X vssd1 vssd1 vccd1 vccd1 _14252_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10415_ _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10415_/Y sky130_fd_sc_hd__nor2_1
X_13203_ _13202_/X _18438_/Q _13203_/S vssd1 vssd1 vccd1 vccd1 _13204_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_88_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17367__A _17424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14183_ _14191_/A _14188_/C vssd1 vssd1 vccd1 vccd1 _14183_/Y sky130_fd_sc_hd__nor2_1
X_11395_ _11404_/A _11395_/B vssd1 vssd1 vccd1 vccd1 _11395_/X sky130_fd_sc_hd__or2_1
XFILLER_152_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16271__A _16282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10346_ _10342_/A _10345_/X _09779_/A vssd1 vssd1 vccd1 vccd1 _10346_/Y sky130_fd_sc_hd__o21ai_1
X_13134_ input2/X _13091_/X _13094_/X vssd1 vssd1 vccd1 vccd1 _13134_/X sky130_fd_sc_hd__a21o_1
X_18991_ _18992_/CLK _18991_/D vssd1 vssd1 vccd1 vccd1 _18991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output163_A _12776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17942_ _19841_/Q _17078_/X _17948_/S vssd1 vssd1 vccd1 vccd1 _17943_/A sky130_fd_sc_hd__mux2_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13065_ _17659_/A vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__buf_2
X_10277_ _19375_/Q _19710_/Q _10277_/S vssd1 vssd1 vccd1 vccd1 _10278_/B sky130_fd_sc_hd__mux2_1
XFILLER_112_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12304__A _12340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ _18753_/Q _18748_/Q _12015_/Y _12064_/A vssd1 vssd1 vccd1 vccd1 _12016_/X
+ sky130_fd_sc_hd__a31o_1
X_17873_ _17873_/A vssd1 vssd1 vccd1 vccd1 _19810_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19612_ _19935_/CLK _19612_/D vssd1 vssd1 vccd1 vccd1 _19612_/Q sky130_fd_sc_hd__dfxtp_1
X_16824_ _16384_/X _19378_/Q _16830_/S vssd1 vssd1 vccd1 vccd1 _16825_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19543_ _19960_/CLK _19543_/D vssd1 vssd1 vccd1 vccd1 _19543_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09613__A _09646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16755_ _16755_/A vssd1 vssd1 vccd1 vccd1 _19347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13967_ _13967_/A _13973_/C vssd1 vssd1 vccd1 vccd1 _13967_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10759__A _10760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15706_ _09481_/D _11865_/A _13700_/X _14529_/A vssd1 vssd1 vccd1 vccd1 _15706_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11294__A1 _11186_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19474_ _19868_/CLK _19474_/D vssd1 vssd1 vccd1 vccd1 _19474_/Q sky130_fd_sc_hd__dfxtp_1
X_12918_ _18827_/Q _12918_/B vssd1 vssd1 vccd1 vccd1 _16846_/C sky130_fd_sc_hd__nand2_4
XANTENNA__09332__B _18938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16686_ _16686_/A vssd1 vssd1 vccd1 vccd1 _19317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13898_ _18539_/Q _13893_/X _12580_/X _12584_/Y _13897_/X vssd1 vssd1 vccd1 vccd1
+ _18539_/D sky130_fd_sc_hd__o221a_1
X_18425_ _20010_/CLK _18425_/D vssd1 vssd1 vccd1 vccd1 _18425_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15637_ _15637_/A vssd1 vssd1 vccd1 vccd1 _18897_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13035__A2 _13189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ _12851_/A _12849_/B vssd1 vssd1 vccd1 vccd1 _12849_/Y sky130_fd_sc_hd__nor2_4
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18356_ _18356_/A vssd1 vssd1 vccd1 vccd1 _20009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15568_ _15568_/A vssd1 vssd1 vccd1 vccd1 _18867_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17307_ _17131_/X _19569_/Q _17315_/S vssd1 vssd1 vccd1 vccd1 _17308_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17976__S _17976_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14519_ _14518_/A _14518_/C _18740_/Q vssd1 vssd1 vccd1 vccd1 _14520_/C sky130_fd_sc_hd__a21oi_1
X_18287_ _17643_/X _19979_/Q _18291_/S vssd1 vssd1 vccd1 vccd1 _18288_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15499_ _15384_/X _15494_/Y _15498_/Y vssd1 vssd1 vccd1 vccd1 _15500_/C sky130_fd_sc_hd__a21oi_1
X_17238_ _17238_/A vssd1 vssd1 vccd1 vccd1 _19538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17169_ _17169_/A vssd1 vssd1 vccd1 vccd1 _19511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ _10355_/A _09986_/X _10064_/A vssd1 vssd1 vccd1 vccd1 _09991_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13259__C1 _13307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15799__B2 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13274__A2 _11683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17740__A _17808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12482__B1 _18774_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11380__S1 _11208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09425_ _18822_/Q _09425_/B vssd1 vssd1 vccd1 vccd1 _12066_/B sky130_fd_sc_hd__and2_1
XFILLER_53_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _09354_/B _09352_/Y _13340_/A vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__a21o_2
XANTENNA__16075__B _16075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09287_ _09287_/A _09491_/A _09287_/C _09287_/D vssd1 vssd1 vccd1 vccd1 _09289_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16091__A _16148_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ _10200_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__or2_1
XFILLER_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11180_ _18428_/Q _19457_/Q _19494_/Q _19068_/Q _11293_/A _09737_/A vssd1 vssd1 vccd1
+ vccd1 _11180_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10131_ _19682_/Q _19448_/Q _18513_/Q _19778_/Q _10447_/S _10398_/A vssd1 vssd1 vccd1
+ vccd1 _10131_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11760__A2 _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10062_ _19152_/Q _19413_/Q _19312_/Q _19647_/Q _09918_/S _09646_/A vssd1 vssd1 vccd1
+ vccd1 _10063_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17126__S _17129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10946__S1 _10624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870_ _15254_/B _15449_/B _14908_/S vssd1 vssd1 vccd1 vccd1 _14870_/X sky130_fd_sc_hd__mux2_1
X_13821_ _13821_/A vssd1 vssd1 vccd1 vccd1 _18505_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09433__A _15457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15154__B _15160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_opt_8_0_clock _19379_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_8_0_clock/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16540_ _16540_/A vssd1 vssd1 vccd1 vccd1 _19252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11276__B2 _11278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13752_ _18485_/Q _13751_/X _13752_/S vssd1 vssd1 vccd1 vccd1 _13753_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ _11149_/A _10964_/B vssd1 vssd1 vccd1 vccd1 _10964_/X sky130_fd_sc_hd__or2_1
XFILLER_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11371__S1 _11322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ _18544_/Q _12673_/X _12699_/Y _12702_/Y vssd1 vssd1 vccd1 vccd1 _12703_/X
+ sky130_fd_sc_hd__o22a_4
X_16471_ _16471_/A vssd1 vssd1 vccd1 vccd1 _19222_/D sky130_fd_sc_hd__clkbuf_1
X_13683_ _19016_/Q _13683_/B vssd1 vssd1 vccd1 vccd1 _13683_/X sky130_fd_sc_hd__or2_1
X_10895_ _10905_/A _10895_/B vssd1 vssd1 vccd1 vccd1 _10895_/X sky130_fd_sc_hd__or2_1
XFILLER_31_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18210_ _18278_/S vssd1 vssd1 vccd1 vccd1 _18219_/S sky130_fd_sc_hd__buf_2
X_15422_ _15082_/A _15424_/B _15081_/X _15421_/X vssd1 vssd1 vccd1 vccd1 _15422_/X
+ sky130_fd_sc_hd__o211a_1
X_19190_ _19877_/CLK _19190_/D vssd1 vssd1 vccd1 vccd1 _19190_/Q sky130_fd_sc_hd__dfxtp_1
X_12634_ _12634_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12634_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12776__A1 _18547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17796__S _17804_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18141_ _17640_/X _19914_/Q _18147_/S vssd1 vssd1 vccd1 vccd1 _18142_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15353_ _15353_/A vssd1 vssd1 vccd1 vccd1 _15353_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12565_ _12632_/A _15424_/A _12541_/A vssd1 vssd1 vccd1 vccd1 _12568_/A sky130_fd_sc_hd__a21oi_1
XFILLER_141_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14304_ _14319_/A _14304_/B vssd1 vssd1 vccd1 vccd1 _14304_/Y sky130_fd_sc_hd__nor2_1
X_11516_ _11595_/A _11599_/A _11595_/C _10653_/A _11515_/X vssd1 vssd1 vccd1 vccd1
+ _11592_/C sky130_fd_sc_hd__a311o_1
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18072_ _18071_/X _19893_/Q _18078_/S vssd1 vssd1 vccd1 vccd1 _18073_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15284_ _15366_/A vssd1 vssd1 vccd1 vccd1 _15284_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12496_ _12442_/A _12442_/B _12469_/A _12495_/Y vssd1 vssd1 vccd1 vccd1 _12497_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_144_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17023_ _17023_/A vssd1 vssd1 vccd1 vccd1 _17023_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14235_ _14234_/A _14234_/B _15807_/A vssd1 vssd1 vccd1 vccd1 _14236_/B sky130_fd_sc_hd__a21o_1
X_11447_ _19386_/Q _11447_/B vssd1 vssd1 vccd1 vccd1 _11447_/X sky130_fd_sc_hd__or2_1
XFILLER_153_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output88_A _12671_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10634__S0 _09726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11378_ _18425_/Q _19454_/Q _19491_/Q _19065_/Q _11212_/A _11077_/A vssd1 vssd1 vccd1
+ vccd1 _11378_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11857__B _11857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ _18627_/Q _14166_/B vssd1 vssd1 vccd1 vccd1 _14172_/C sky130_fd_sc_hd__and2_1
XFILLER_113_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11751__A2 _11748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10329_ _10329_/A _10329_/B vssd1 vssd1 vccd1 vccd1 _10329_/X sky130_fd_sc_hd__and2_1
X_13117_ _13117_/A vssd1 vssd1 vccd1 vccd1 _18433_/D sky130_fd_sc_hd__clkbuf_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18420__S _18422_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18974_ _18974_/CLK _18974_/D vssd1 vssd1 vccd1 vccd1 _18974_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _14143_/A _14097_/B _14097_/C vssd1 vssd1 vccd1 vccd1 _18608_/D sky130_fd_sc_hd__nor3_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _17925_/A vssd1 vssd1 vccd1 vccd1 _19833_/D sky130_fd_sc_hd__clkbuf_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _18797_/Q _13048_/B vssd1 vssd1 vccd1 vccd1 _13048_/X sky130_fd_sc_hd__and2_1
XFILLER_59_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12969__A _19488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17856_ _17867_/A vssd1 vssd1 vccd1 vccd1 _17865_/S sky130_fd_sc_hd__buf_6
XFILLER_22_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_1_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16807_ _16807_/A vssd1 vssd1 vccd1 vccd1 _19370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16875__S _16881_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17787_ _17704_/X _19772_/Q _17793_/S vssd1 vssd1 vccd1 vccd1 _17788_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14999_ _14991_/X _15002_/B _14997_/X _14998_/X vssd1 vssd1 vccd1 vccd1 _14999_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11267__A1 _09550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16738_ _16749_/A vssd1 vssd1 vccd1 vccd1 _16747_/S sky130_fd_sc_hd__buf_4
X_19526_ _19526_/CLK _19526_/D vssd1 vssd1 vccd1 vccd1 _19526_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19457_ _19949_/CLK _19457_/D vssd1 vssd1 vccd1 vccd1 _19457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16669_ _16669_/A vssd1 vssd1 vccd1 vccd1 _19309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09210_ _13226_/A vssd1 vssd1 vccd1 vccd1 _13473_/A sky130_fd_sc_hd__clkbuf_1
X_18408_ _18408_/A vssd1 vssd1 vccd1 vccd1 _20033_/D sky130_fd_sc_hd__clkbuf_1
X_19388_ _19526_/CLK _19388_/D vssd1 vssd1 vccd1 vccd1 _19388_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11114__S1 _10854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18339_ _18339_/A vssd1 vssd1 vccd1 vccd1 _20002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10778__B1 _10712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13716__B1 _13700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14424__A _14472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11259__S _11270_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09974_ _10549_/A vssd1 vssd1 vccd1 vccd1 _10553_/A sky130_fd_sc_hd__buf_2
XFILLER_130_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14692__A1 _13572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_36_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09408_ _11785_/A _09408_/B vssd1 vssd1 vccd1 vccd1 _13335_/B sky130_fd_sc_hd__nor2_4
XFILLER_158_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10680_ _10680_/A _10680_/B vssd1 vssd1 vccd1 vccd1 _10680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09339_ _14821_/A _11903_/A _09338_/X vssd1 vssd1 vccd1 vccd1 _09339_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _12350_/A vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10864__S0 _10953_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11301_ _19323_/Q _19594_/Q _19818_/Q _19562_/Q _11230_/X _11021_/A vssd1 vssd1 vccd1
+ vccd1 _11301_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12281_ _18464_/Q _12556_/A _12557_/A vssd1 vssd1 vccd1 vccd1 _12281_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16025__S _16031_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14020_ _18581_/Q _14017_/B _14019_/X vssd1 vssd1 vccd1 vccd1 _14020_/Y sky130_fd_sc_hd__a21oi_1
X_11232_ _11344_/A _11232_/B vssd1 vssd1 vccd1 vccd1 _11232_/X sky130_fd_sc_hd__or2_1
XFILLER_153_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11163_ _19134_/Q _19395_/Q _19294_/Q _19629_/Q _11293_/A _11015_/A vssd1 vssd1 vccd1
+ vccd1 _11164_/B sky130_fd_sc_hd__mux4_1
XFILLER_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10941__B1 _09546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10114_ _10415_/A _10114_/B vssd1 vssd1 vccd1 vccd1 _10114_/Y sky130_fd_sc_hd__nor2_1
X_11094_ _20016_/Q _19854_/Q _19263_/Q _19033_/Q _11158_/S _11022_/A vssd1 vssd1 vccd1
+ vccd1 _11094_/X sky130_fd_sc_hd__mux4_1
X_15971_ _19019_/Q _15951_/X _15970_/X vssd1 vssd1 vccd1 vccd1 _19019_/D sky130_fd_sc_hd__a21o_1
XFILLER_121_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14683__A1 hold7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17710_ _17710_/A vssd1 vssd1 vccd1 vccd1 _17710_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10045_ _18858_/Q vssd1 vssd1 vccd1 vccd1 _10045_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14922_ _14894_/X _14919_/X _14922_/S vssd1 vssd1 vccd1 vccd1 _14922_/X sky130_fd_sc_hd__mux2_1
X_18690_ _19882_/CLK _18690_/D vssd1 vssd1 vccd1 vccd1 _18690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17641_ _17640_/X _19720_/Q _17650_/S vssd1 vssd1 vccd1 vccd1 _17642_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14853_ _14990_/A _15004_/A _14990_/C vssd1 vssd1 vccd1 vccd1 _14854_/S sky130_fd_sc_hd__or3_1
XANTENNA__16695__S _16703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output126_A _12857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13804_ _18500_/Q _13803_/X _13804_/S vssd1 vssd1 vccd1 vccd1 _13805_/A sky130_fd_sc_hd__mux2_1
X_17572_ _17572_/A vssd1 vssd1 vccd1 vccd1 _19690_/D sky130_fd_sc_hd__clkbuf_1
X_14784_ _14800_/A _14784_/B vssd1 vssd1 vccd1 vccd1 _14785_/A sky130_fd_sc_hd__and2_1
XFILLER_16_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11996_ _12583_/A vssd1 vssd1 vccd1 vccd1 _12790_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19311_ _20003_/CLK _19311_/D vssd1 vssd1 vccd1 vccd1 _19311_/Q sky130_fd_sc_hd__dfxtp_1
X_16523_ _16523_/A vssd1 vssd1 vccd1 vccd1 _19244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13735_ _18483_/Q _13734_/X _13752_/S vssd1 vssd1 vccd1 vccd1 _13736_/A sky130_fd_sc_hd__mux2_1
X_10947_ _10947_/A _10947_/B vssd1 vssd1 vccd1 vccd1 _10947_/X sky130_fd_sc_hd__or2_1
XFILLER_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19242_ _19995_/CLK _19242_/D vssd1 vssd1 vccd1 vccd1 _19242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16454_ _16454_/A vssd1 vssd1 vccd1 vccd1 _19214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13666_ _13709_/A _19014_/Q vssd1 vssd1 vccd1 vccd1 _13666_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ _10727_/A _10877_/X _10719_/A vssd1 vssd1 vccd1 vccd1 _10878_/X sky130_fd_sc_hd__o21a_1
X_15405_ _15405_/A vssd1 vssd1 vccd1 vccd1 _15405_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19173_ _19989_/CLK _19173_/D vssd1 vssd1 vccd1 vccd1 _19173_/Q sky130_fd_sc_hd__dfxtp_1
X_12617_ _12617_/A _12617_/B vssd1 vssd1 vccd1 vccd1 _12621_/A sky130_fd_sc_hd__nor2_2
X_16385_ _16384_/X _19186_/Q _16394_/S vssd1 vssd1 vccd1 vccd1 _16386_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _18464_/Q _13596_/X _13617_/S vssd1 vssd1 vccd1 vccd1 _13598_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18124_ _18861_/Q _13727_/X _18130_/S vssd1 vssd1 vccd1 vccd1 _18124_/X sky130_fd_sc_hd__mux2_1
X_15336_ _15286_/X _15338_/B _15287_/X _15335_/X vssd1 vssd1 vccd1 vccd1 _15336_/X
+ sky130_fd_sc_hd__o211a_1
X_12548_ _12518_/A _14886_/A _12547_/X vssd1 vssd1 vccd1 vccd1 _12548_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18055_ _18054_/X _19888_/Q _18061_/S vssd1 vssd1 vccd1 vccd1 _18056_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15267_ _15211_/X _15270_/B _15212_/X _15266_/X vssd1 vssd1 vccd1 vccd1 _15267_/X
+ sky130_fd_sc_hd__o211a_1
X_12479_ _12470_/Y _12478_/Y _12479_/S vssd1 vssd1 vccd1 vccd1 _12479_/X sky130_fd_sc_hd__mux2_1
X_17006_ _17006_/A vssd1 vssd1 vccd1 vccd1 _19456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10607__S0 _10655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ _18645_/Q _14216_/B _14203_/X vssd1 vssd1 vccd1 vccd1 _14218_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15198_ _15113_/X _15110_/X _15198_/S vssd1 vssd1 vccd1 vccd1 _15198_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11724__A2 _11717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14149_ _14153_/B _14153_/C _14148_/Y vssd1 vssd1 vccd1 vccd1 _18622_/D sky130_fd_sc_hd__o21a_1
XANTENNA__18150__S _18158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18957_ _18960_/CLK _18957_/D vssd1 vssd1 vccd1 vccd1 _18957_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17908_ _17908_/A vssd1 vssd1 vccd1 vccd1 _19825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _09690_/A vssd1 vssd1 vccd1 vccd1 _09690_/X sky130_fd_sc_hd__clkbuf_4
X_18888_ _18923_/CLK _18888_/D vssd1 vssd1 vccd1 vccd1 _18888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10160__A1 _10438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17839_ _19795_/Q _17033_/X _17843_/S vssd1 vssd1 vccd1 vccd1 _17840_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11108__A _11108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15803__A _15813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10012__A _10153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19509_ _20028_/CLK _19509_/D vssd1 vssd1 vccd1 vccd1 _19509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11099__S0 _11186_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11412__A1 _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__S0 _10797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11778__A _12060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14154__A _14189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13993__A _14010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10074__S1 _09646_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15311__C1 _15275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09957_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13468__A2 _13511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_183_clock clkbuf_opt_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _18975_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09888_ _18453_/Q _19482_/Q _19519_/Q _19093_/Q _09898_/S _09895_/A vssd1 vssd1 vccd1
+ vccd1 _09888_/X sky130_fd_sc_hd__mux4_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12402__A _12416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10687__C1 _09820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _18802_/Q _11841_/X _11843_/X _12349_/A _11849_/X vssd1 vssd1 vccd1 vccd1
+ _11857_/B sky130_fd_sc_hd__a221o_2
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09711__A _10572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801_ _10843_/A _10798_/X _10800_/X vssd1 vssd1 vccd1 vccd1 _10801_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09844__A1 _09702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ _11817_/A vssd1 vssd1 vccd1 vccd1 _12984_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14329__A _18674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09844__B2 _18863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13520_ _13520_/A vssd1 vssd1 vccd1 vccd1 _13690_/A sky130_fd_sc_hd__clkbuf_2
X_10732_ _11481_/A _10731_/X _09685_/A vssd1 vssd1 vccd1 vccd1 _10732_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09430__B _15719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_121_clock clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 _20038_/CLK sky130_fd_sc_hd__clkbuf_16
X_13451_ _19910_/Q _13451_/B vssd1 vssd1 vccd1 vccd1 _13451_/X sky130_fd_sc_hd__and2_1
X_10663_ _10663_/A vssd1 vssd1 vccd1 vccd1 _10664_/A sky130_fd_sc_hd__buf_2
XANTENNA__18235__S _18241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12402_ _12416_/B _12402_/B vssd1 vssd1 vccd1 vccd1 _12402_/X sky130_fd_sc_hd__and2_1
X_16170_ _16170_/A vssd1 vssd1 vccd1 vccd1 _19103_/D sky130_fd_sc_hd__clkbuf_1
X_10594_ _10824_/A vssd1 vssd1 vccd1 vccd1 _10832_/A sky130_fd_sc_hd__buf_2
XANTENNA__10837__S0 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13382_ _13307_/X _13371_/Y _13372_/Y _13381_/Y _13460_/A vssd1 vssd1 vccd1 vccd1
+ _13382_/X sky130_fd_sc_hd__a221o_2
XFILLER_127_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12791__B _12791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11688__A _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15121_ _15037_/X _15039_/X _15121_/S vssd1 vssd1 vccd1 vccd1 _15121_/X sky130_fd_sc_hd__mux2_1
X_12333_ _12272_/A _12272_/B _12301_/A _12332_/X vssd1 vssd1 vccd1 vccd1 _12334_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__14064__A _14088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_136_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19909_/CLK sky130_fd_sc_hd__clkbuf_16
X_15052_ _15945_/A vssd1 vssd1 vccd1 vccd1 _15978_/A sky130_fd_sc_hd__buf_2
XFILLER_142_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12264_ _12323_/A _12323_/C _12322_/A vssd1 vssd1 vccd1 vccd1 _12265_/B sky130_fd_sc_hd__o21ai_2
XFILLER_141_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14003_ _18575_/Q _14001_/B _14002_/Y vssd1 vssd1 vccd1 vccd1 _18575_/D sky130_fd_sc_hd__o21a_1
X_11215_ _18428_/Q _19457_/Q _19494_/Q _19068_/Q _11125_/S _11065_/X vssd1 vssd1 vccd1
+ vccd1 _11215_/X sky130_fd_sc_hd__mux4_1
X_19860_ _19989_/CLK _19860_/D vssd1 vssd1 vccd1 vccd1 _19860_/Q sky130_fd_sc_hd__dfxtp_1
X_12195_ _12479_/S _12192_/Y _12194_/X _12154_/X vssd1 vssd1 vccd1 vccd1 _12195_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11262__S0 _10977_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput72 _12273_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[10] sky130_fd_sc_hd__buf_2
X_18811_ _19900_/CLK _18811_/D vssd1 vssd1 vccd1 vccd1 _18811_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput83 _12551_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[20] sky130_fd_sc_hd__buf_2
X_11146_ _18430_/Q _19459_/Q _19496_/Q _19070_/Q _11023_/S _11296_/A vssd1 vssd1 vccd1
+ vccd1 _11146_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10390__A1 _10380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19791_ _19824_/CLK _19791_/D vssd1 vssd1 vccd1 vccd1 _19791_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput94 _12791_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[30] sky130_fd_sc_hd__buf_2
XANTENNA__14656__A1 _13727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15954_ _15954_/A vssd1 vssd1 vccd1 vccd1 _15954_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11077_ _11077_/A vssd1 vssd1 vccd1 vccd1 _11077_/X sky130_fd_sc_hd__buf_2
X_18742_ _18744_/CLK _18742_/D vssd1 vssd1 vccd1 vccd1 _18742_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12131__A2 _12124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _10329_/A vssd1 vssd1 vccd1 vccd1 _10028_/X sky130_fd_sc_hd__buf_2
X_14905_ _14900_/X _14903_/X _15113_/S vssd1 vssd1 vccd1 vccd1 _14905_/X sky130_fd_sc_hd__mux2_1
X_18673_ _18677_/CLK _18673_/D vssd1 vssd1 vccd1 vccd1 _18673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15605__A0 _18884_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15885_ _15897_/A _15885_/B vssd1 vssd1 vccd1 vccd1 _15886_/A sky130_fd_sc_hd__and2_1
XANTENNA__12031__B _12031_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17624_ _17186_/X _19714_/Q _17628_/S vssd1 vssd1 vccd1 vccd1 _17625_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12419__B1 _12154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14836_ _14966_/A _12080_/B _15201_/B vssd1 vssd1 vccd1 vccd1 _15346_/A sky130_fd_sc_hd__a21bo_1
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11890__B2 _18711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17555_ _17555_/A vssd1 vssd1 vccd1 vccd1 _19683_/D sky130_fd_sc_hd__clkbuf_1
X_14767_ _14748_/X _14752_/X _14766_/Y _18823_/Q vssd1 vssd1 vccd1 vccd1 _14768_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09835__A1 _09833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14239__A _14239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11979_ _14931_/A _14865_/A _12029_/A vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__o21ai_1
XFILLER_91_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16506_ _19237_/Q _13800_/X _16508_/S vssd1 vssd1 vccd1 vccd1 _16507_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13718_ _13726_/A _19021_/Q vssd1 vssd1 vccd1 vccd1 _13718_/Y sky130_fd_sc_hd__nand2_1
X_17486_ _17183_/X _19649_/Q _17492_/S vssd1 vssd1 vccd1 vccd1 _17487_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09930__S1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14698_ _14698_/A vssd1 vssd1 vccd1 vccd1 _18800_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16437_ _16459_/A vssd1 vssd1 vccd1 vccd1 _16446_/S sky130_fd_sc_hd__buf_4
XFILLER_108_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19225_ _19523_/CLK _19225_/D vssd1 vssd1 vccd1 vccd1 _19225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13649_ _13654_/B _13647_/Y _13648_/X vssd1 vssd1 vccd1 vccd1 _13649_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_31_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18145__S _18147_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19156_ _19747_/CLK _19156_/D vssd1 vssd1 vccd1 vccd1 _19156_/Q sky130_fd_sc_hd__dfxtp_1
X_16368_ _17704_/A vssd1 vssd1 vccd1 vccd1 _16368_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10828__S0 _10764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18107_ _18107_/A vssd1 vssd1 vccd1 vccd1 _19903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15319_ _15286_/X _15321_/B _15287_/X _15318_/X vssd1 vssd1 vccd1 vccd1 _15319_/X
+ sky130_fd_sc_hd__o211a_1
X_19087_ _19583_/CLK _19087_/D vssd1 vssd1 vccd1 vccd1 _19087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16299_ _17426_/A _18208_/B vssd1 vssd1 vccd1 vccd1 _16381_/A sky130_fd_sc_hd__or2_2
XFILLER_173_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13147__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18038_ _18037_/Y _19883_/Q _18044_/S vssd1 vssd1 vccd1 vccd1 _18039_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11253__S0 _11212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20000_ _20032_/CLK _20000_/D vssd1 vssd1 vccd1 vccd1 _20000_/Q sky130_fd_sc_hd__dfxtp_1
X_09811_ _19350_/Q _19621_/Q _19845_/Q _19589_/Q _09898_/S _09895_/A vssd1 vssd1 vccd1
+ vccd1 _09812_/B sky130_fd_sc_hd__mux4_1
XFILLER_28_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19989_ _19989_/CLK _19989_/D vssd1 vssd1 vccd1 vccd1 _19989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09742_ _10638_/A vssd1 vssd1 vccd1 vccd1 _10522_/A sky130_fd_sc_hd__buf_2
XFILLER_140_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11005__S0 _11048_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13318__A _13340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09749__S1 _09895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09673_ _19685_/Q _19451_/Q _18516_/Q _19781_/Q _09855_/A _09642_/A vssd1 vssd1 vccd1
+ vccd1 _09673_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17224__S _17232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11308__S1 _11108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09531__A _19487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13083__B1 _13082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_53_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19960_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15780__C1 _13885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10295__S1 _10329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11492__S0 _10906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14335__B1 _18676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09409__C _13335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19622_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__18077__A1 _13621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11000_ _19921_/Q _19535_/Q _19985_/Q _19104_/Q _11048_/S _10978_/A vssd1 vssd1 vccd1
+ vccd1 _11001_/B sky130_fd_sc_hd__mux4_1
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12649__A0 _12645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13228__A _13360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09425__B _09425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12132__A _18459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ _18792_/Q _11841_/X _12949_/X _12950_/X vssd1 vssd1 vccd1 vccd1 _12951_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16691__C_N _16298_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _12831_/A vssd1 vssd1 vccd1 vccd1 _12827_/A sky130_fd_sc_hd__buf_6
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11872__A1 _18477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15670_ _15670_/A vssd1 vssd1 vccd1 vccd1 _18912_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _18678_/Q vssd1 vssd1 vccd1 vccd1 _14345_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09441__A input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14621_ _14621_/A vssd1 vssd1 vccd1 vccd1 _18774_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _14544_/B _11860_/B _11860_/C _11833_/D vssd1 vssd1 vccd1 vccd1 _11833_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10587__A _10587_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16973__S _16975_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14059__A _14102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17179_/X _19584_/Q _17348_/S vssd1 vssd1 vccd1 vccd1 _17341_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14552_/A _18994_/Q vssd1 vssd1 vccd1 vccd1 _14552_/Y sky130_fd_sc_hd__nand2_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11731_/X _11761_/X _11762_/Y _13660_/A _19012_/Q vssd1 vssd1 vccd1 vccd1
+ _11764_/X sky130_fd_sc_hd__a32o_4
XFILLER_159_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13503_ _13503_/A vssd1 vssd1 vccd1 vccd1 _18455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10836_/A _10715_/B vssd1 vssd1 vccd1 vccd1 _10715_/Y sky130_fd_sc_hd__nor2_1
X_17271_ _17271_/A vssd1 vssd1 vccd1 vccd1 _19553_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14483_ _14485_/A _14485_/C _14465_/X vssd1 vssd1 vccd1 vccd1 _14483_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16563__A1 _13778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11695_ _11695_/A vssd1 vssd1 vccd1 vccd1 _13054_/B sky130_fd_sc_hd__buf_4
XFILLER_9_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19010_ _19010_/CLK _19010_/D vssd1 vssd1 vccd1 vccd1 _19010_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_174_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16222_ _16222_/A vssd1 vssd1 vccd1 vccd1 _19127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13434_ _18610_/Q vssd1 vssd1 vccd1 vccd1 _14105_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ _10630_/A _10645_/X _10579_/A vssd1 vssd1 vccd1 vccd1 _10646_/X sky130_fd_sc_hd__o21a_1
XFILLER_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16153_ _16221_/S vssd1 vssd1 vccd1 vccd1 _16162_/S sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_158_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10286__S1 _10283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13365_ _17713_/A vssd1 vssd1 vccd1 vccd1 _13365_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10577_ _19145_/Q _19406_/Q _19305_/Q _19640_/Q _10521_/X _10522_/X vssd1 vssd1 vccd1
+ vccd1 _10577_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13129__A1 _13588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ _15101_/X _15100_/B _15102_/X _15103_/X vssd1 vssd1 vccd1 vccd1 _15104_/X
+ sky130_fd_sc_hd__o211a_1
X_12316_ _12316_/A _12536_/A _15916_/A vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__and3_2
X_16084_ _16084_/A vssd1 vssd1 vccd1 vccd1 _19065_/D sky130_fd_sc_hd__clkbuf_1
X_13296_ _18853_/Q _13665_/B _13458_/A vssd1 vssd1 vccd1 vccd1 _13296_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17309__S _17315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15035_ _15031_/X _15034_/X _15132_/S vssd1 vssd1 vccd1 vccd1 _15035_/X sky130_fd_sc_hd__mux2_1
X_19912_ _19912_/CLK _19912_/D vssd1 vssd1 vccd1 vccd1 _19912_/Q sky130_fd_sc_hd__dfxtp_1
X_12247_ _18527_/Q vssd1 vssd1 vccd1 vccd1 _12277_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__11235__S0 _11156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16213__S _16217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__S1 _09637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14522__A _14529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09616__A _11538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19843_ _20037_/CLK _19843_/D vssd1 vssd1 vccd1 vccd1 _19843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10363__A1 _09566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ _15219_/A _12178_/B vssd1 vssd1 vccd1 vccd1 _12217_/A sky130_fd_sc_hd__xor2_1
XFILLER_110_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13138__A _13502_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11129_ _19326_/Q _19597_/Q _19821_/Q _19565_/Q _11258_/S _11050_/A vssd1 vssd1 vccd1
+ vccd1 _11129_/X sky130_fd_sc_hd__mux4_1
X_19774_ _20032_/CLK _19774_/D vssd1 vssd1 vccd1 vccd1 _19774_/Q sky130_fd_sc_hd__dfxtp_1
X_16986_ _16393_/X _19450_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16987_/A sky130_fd_sc_hd__mux2_1
X_18725_ _18741_/CLK _18725_/D vssd1 vssd1 vccd1 vccd1 _18725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15937_ _19005_/Q _15927_/X _15928_/X _15936_/Y vssd1 vssd1 vccd1 vccd1 _19005_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12977__A _17004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17044__S _17056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15868_ _15881_/A _16841_/B vssd1 vssd1 vccd1 vccd1 _15869_/A sky130_fd_sc_hd__and2_1
X_18656_ _18660_/CLK _18656_/D vssd1 vssd1 vccd1 vccd1 _18656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17607_ _17607_/A vssd1 vssd1 vccd1 vccd1 _19706_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17979__S _17987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14819_ _14819_/A _14819_/B vssd1 vssd1 vccd1 vccd1 _14819_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15799_ _09481_/B _11860_/A _15798_/X input56/X vssd1 vssd1 vccd1 vccd1 _15800_/B
+ sky130_fd_sc_hd__a22o_1
X_18587_ _18655_/CLK _18587_/D vssd1 vssd1 vccd1 vccd1 _18587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17538_ _19675_/Q vssd1 vssd1 vccd1 vccd1 _17539_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_32_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17469_ _17469_/A vssd1 vssd1 vccd1 vccd1 _19641_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19208_ _19976_/CLK _19208_/D vssd1 vssd1 vccd1 vccd1 _19208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13958__D _13958_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19139_ _19637_/CLK _19139_/D vssd1 vssd1 vccd1 vccd1 _19139_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12040__A1 _18900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10029__S1 _10028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17219__S _17221_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15528__A _15553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__S0 _11293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11551__B1 _09547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15817__B1 _15798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09725_ _09725_/A vssd1 vssd1 vccd1 vccd1 _09726_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13482__S _13502_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11791__A _11791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ _10058_/A vssd1 vssd1 vccd1 vccd1 _09657_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10201__S1 _09636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09261__A _09261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17889__S _17893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16793__S _16797_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09587_ _11273_/A vssd1 vssd1 vccd1 vccd1 _10775_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10200__A _10200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12803__B1 _12866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15710__B _15740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11082__A2 _11060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16545__A1 _13857_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10500_ _10549_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10500_/X sky130_fd_sc_hd__or2_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13511__A _13511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11480_ _19205_/Q _19796_/Q _19958_/Q _19173_/Q _10708_/X _10710_/X vssd1 vssd1 vccd1
+ vccd1 _11481_/B sky130_fd_sc_hd__mux4_1
XFILLER_155_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10431_ _10484_/A _10430_/X _10382_/X vssd1 vssd1 vccd1 vccd1 _10431_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_137_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11465__S0 _10821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09983__A0 _19680_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ _17672_/A vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10362_ _10064_/A _10361_/X _09980_/A vssd1 vssd1 vccd1 vccd1 _10362_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12101_ _18755_/Q _18751_/Q vssd1 vssd1 vccd1 vccd1 _12101_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17129__S _17129_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ _19936_/Q _19550_/Q _20000_/Q _19119_/Q _10037_/S _10329_/A vssd1 vssd1 vccd1
+ vccd1 _10294_/B sky130_fd_sc_hd__mux4_1
XFILLER_124_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11217__S0 _11212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13081_ _13081_/A vssd1 vssd1 vccd1 vccd1 _13081_/X sky130_fd_sc_hd__buf_2
XFILLER_105_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12032_ _18979_/Q vssd1 vssd1 vccd1 vccd1 _12032_/X sky130_fd_sc_hd__buf_4
XANTENNA__11685__B _11790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17653__A _17736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16840_ _16840_/A vssd1 vssd1 vccd1 vccd1 _19385_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14996__B _14996_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16771_ _16307_/X _19354_/Q _16775_/S vssd1 vssd1 vccd1 vccd1 _16772_/A sky130_fd_sc_hd__mux2_1
X_13983_ _13991_/A _13983_/B _13984_/B vssd1 vssd1 vccd1 vccd1 _18568_/D sky130_fd_sc_hd__nor3_1
XFILLER_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13295__B1 _13292_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18510_ _20032_/CLK _18510_/D vssd1 vssd1 vccd1 vccd1 _18510_/Q sky130_fd_sc_hd__dfxtp_1
X_15722_ _18935_/Q _15745_/B vssd1 vssd1 vccd1 vccd1 _15722_/X sky130_fd_sc_hd__or2_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12934_ _12934_/A _12956_/A vssd1 vssd1 vccd1 vccd1 _12934_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _20010_/CLK _19490_/D vssd1 vssd1 vccd1 vccd1 _19490_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_84_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ _19864_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15653_ _18905_/Q _12234_/A _15655_/S vssd1 vssd1 vccd1 vccd1 _15654_/A sky130_fd_sc_hd__mux2_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _12865_/A vssd1 vssd1 vccd1 vccd1 _12865_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14604_/A vssd1 vssd1 vccd1 vccd1 _18769_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11206__A _11206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _17662_/X _20017_/Q _18374_/S vssd1 vssd1 vccd1 vccd1 _18373_/A sky130_fd_sc_hd__mux2_1
X_11816_ _13269_/A vssd1 vssd1 vccd1 vccd1 _11841_/A sky130_fd_sc_hd__clkbuf_2
X_15584_ _15584_/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__clkbuf_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12791_/X _12794_/X _12795_/X vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__o21a_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _17323_/A vssd1 vssd1 vccd1 vccd1 _19576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14535_/A vssd1 vssd1 vccd1 vccd1 _18750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11897_/A _19011_/Q vssd1 vssd1 vccd1 vccd1 _11747_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17254_ _17160_/X _19546_/Q _17254_/S vssd1 vssd1 vccd1 vccd1 _17255_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10281__B1 _10162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14466_ _14468_/A _14468_/C _14465_/X vssd1 vssd1 vccd1 vccd1 _14466_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _11727_/A vssd1 vssd1 vccd1 vccd1 _14670_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_30_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16205_ _16205_/A vssd1 vssd1 vccd1 vccd1 _19119_/D sky130_fd_sc_hd__clkbuf_1
X_13417_ _18609_/Q _11851_/X _13194_/X _18741_/Q vssd1 vssd1 vccd1 vccd1 _13417_/X
+ sky130_fd_sc_hd__a22o_1
X_10629_ _19208_/Q _19799_/Q _19961_/Q _19176_/Q _10691_/S _10626_/X vssd1 vssd1 vccd1
+ vccd1 _10630_/B sky130_fd_sc_hd__mux4_1
X_17185_ _17185_/A vssd1 vssd1 vccd1 vccd1 _19516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14397_ _14398_/B _14398_/C _18695_/Q vssd1 vssd1 vccd1 vccd1 _14399_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14562__A3 _09341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16136_ _13385_/X _19089_/Q _16144_/S vssd1 vssd1 vccd1 vccd1 _16137_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ _13688_/A _13357_/C vssd1 vssd1 vccd1 vccd1 _13348_/X sky130_fd_sc_hd__xor2_1
XFILLER_155_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10584__A1 _09883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16067_ _19060_/Q _16066_/X _16073_/S vssd1 vssd1 vccd1 vccd1 _16068_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13279_ _13068_/X _13278_/X _13005_/X vssd1 vssd1 vccd1 vccd1 _13279_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_170_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15018_ _14925_/X _14928_/X _15023_/S vssd1 vssd1 vccd1 vccd1 _15018_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19826_ _19829_/CLK _19826_/D vssd1 vssd1 vccd1 vccd1 _19826_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17563__A _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12089__A1 _18901_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19757_ _19757_/CLK _19757_/D vssd1 vssd1 vccd1 vccd1 _19757_/Q sky130_fd_sc_hd__dfxtp_1
X_16969_ _16368_/X _19442_/Q _16975_/S vssd1 vssd1 vccd1 vccd1 _16970_/A sky130_fd_sc_hd__mux2_1
X_09510_ _11948_/B _09510_/B vssd1 vssd1 vccd1 vccd1 _09510_/X sky130_fd_sc_hd__or2_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18708_ _19912_/CLK _18708_/D vssd1 vssd1 vccd1 vccd1 _18708_/Q sky130_fd_sc_hd__dfxtp_1
X_19688_ _19720_/CLK _19688_/D vssd1 vssd1 vccd1 vccd1 _19688_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12500__A _12501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__S0 _10354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09441_ input70/X vssd1 vssd1 vccd1 vccd1 _14665_/A sky130_fd_sc_hd__inv_2
XFILLER_25_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18639_ _18688_/CLK _18639_/D vssd1 vssd1 vccd1 vccd1 _18639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09372_ _18952_/Q _18951_/Q _18950_/Q _18949_/Q vssd1 vssd1 vccd1 vccd1 _09407_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09888__S0 _09898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14427__A _14427_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10166__S _10166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18333__S _18335_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10575__A1 _10690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10690__A _10690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10422__S1 _10153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_106_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13277__B1 _13272_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09708_ _11500_/A vssd1 vssd1 vccd1 vccd1 _10211_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10980_ _10980_/A vssd1 vssd1 vccd1 vccd1 _11270_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10186__S0 _09655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16215__A0 _13443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09639_ _09642_/A vssd1 vssd1 vccd1 vccd1 _09639_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17412__S _17420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12650_ _18478_/Q _12010_/X _12530_/A vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__o21a_1
XFILLER_169_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11601_ _11617_/B vssd1 vssd1 vccd1 vccd1 _11601_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _12562_/A _12582_/C _18778_/Q vssd1 vssd1 vccd1 vccd1 _12581_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_169_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14320_ _18671_/Q _14316_/X _14319_/Y vssd1 vssd1 vccd1 vccd1 _18671_/D sky130_fd_sc_hd__o21a_1
X_11532_ _19255_/Q _19750_/Q _11532_/S vssd1 vssd1 vccd1 vccd1 _11533_/B sky130_fd_sc_hd__mux2_1
XFILLER_169_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251_ _18651_/Q _14247_/B _14250_/Y vssd1 vssd1 vccd1 vccd1 _18651_/D sky130_fd_sc_hd__o21a_1
X_11463_ _15936_/B _12839_/B vssd1 vssd1 vccd1 vccd1 _11463_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15741__A2 _15738_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13202_ _17681_/A vssd1 vssd1 vccd1 vccd1 _13202_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10414_ _19212_/Q _19803_/Q _19965_/Q _19180_/Q _10314_/S _10109_/X vssd1 vssd1 vccd1
+ vccd1 _10415_/B sky130_fd_sc_hd__mux4_1
XFILLER_143_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_opt_4_0_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_165_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14182_ _18633_/Q _14182_/B vssd1 vssd1 vccd1 vccd1 _14188_/C sky130_fd_sc_hd__and2_1
XFILLER_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11394_ _19321_/Q _19592_/Q _19816_/Q _19560_/Q _11153_/A _11019_/A vssd1 vssd1 vccd1
+ vccd1 _11395_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10110__S0 _10314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13387__S _13464_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13133_ _13268_/A _13129_/X _13132_/X vssd1 vssd1 vccd1 vccd1 _13133_/X sky130_fd_sc_hd__a21bo_1
XFILLER_174_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10345_ _18446_/Q _19475_/Q _19512_/Q _19086_/Q _10005_/A _10223_/X vssd1 vssd1 vccd1
+ vccd1 _10345_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10661__S1 _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14072__A _14088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18990_ _18992_/CLK _18990_/D vssd1 vssd1 vccd1 vccd1 _18990_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_98_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _17941_/A vssd1 vssd1 vccd1 vccd1 _19840_/D sky130_fd_sc_hd__clkbuf_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _17017_/A vssd1 vssd1 vccd1 vccd1 _17659_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10276_ _09939_/A _10253_/Y _10275_/Y _09747_/A vssd1 vssd1 vccd1 vccd1 _10276_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_105_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output156_A _12608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ _18754_/Q _18749_/Q vssd1 vssd1 vccd1 vccd1 _12015_/Y sky130_fd_sc_hd__nand2_1
X_17872_ _19810_/Q _17081_/X _17876_/S vssd1 vssd1 vccd1 vccd1 _17873_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10105__A _15970_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19611_ _19965_/CLK _19611_/D vssd1 vssd1 vccd1 vccd1 _19611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16823_ _16823_/A vssd1 vssd1 vccd1 vccd1 _19377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19542_ _20024_/CLK _19542_/D vssd1 vssd1 vccd1 vccd1 _19542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16754_ _19347_/Q _13845_/X _16758_/S vssd1 vssd1 vccd1 vccd1 _16755_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13966_ _18563_/Q _13966_/B vssd1 vssd1 vccd1 vccd1 _13973_/C sky130_fd_sc_hd__and2_2
XFILLER_81_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10759__B _12843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12917_ _15735_/A _16474_/B _16150_/B vssd1 vssd1 vccd1 vccd1 _17738_/A sky130_fd_sc_hd__or3_2
X_15705_ _15765_/A vssd1 vssd1 vccd1 vccd1 _15705_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19473_ _19581_/CLK _19473_/D vssd1 vssd1 vccd1 vccd1 _19473_/Q sky130_fd_sc_hd__dfxtp_1
X_16685_ _16393_/X _19317_/Q _16685_/S vssd1 vssd1 vccd1 vccd1 _16686_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18418__S _18418_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897_ _14385_/A vssd1 vssd1 vccd1 vccd1 _13897_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17322__S _17326_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18424_ _20010_/CLK _18424_/D vssd1 vssd1 vccd1 vccd1 _18424_/Q sky130_fd_sc_hd__dfxtp_1
X_12848_ _12851_/A _12848_/B vssd1 vssd1 vccd1 vccd1 _12848_/Y sky130_fd_sc_hd__nor2_4
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15636_ _18897_/Q _18518_/Q _15644_/S vssd1 vssd1 vccd1 vccd1 _15637_/A sky130_fd_sc_hd__mux2_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18355_ _17634_/X _20009_/Q _18363_/S vssd1 vssd1 vccd1 vccd1 _18356_/A sky130_fd_sc_hd__mux2_1
X_15567_ _13504_/A _18899_/Q _15567_/S vssd1 vssd1 vccd1 vccd1 _15568_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _14993_/A _12755_/A _12758_/B vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14247__A _14265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17306_ _17352_/S vssd1 vssd1 vccd1 vccd1 _17315_/S sky130_fd_sc_hd__clkbuf_4
X_14518_ _14518_/A _18740_/Q _14518_/C vssd1 vssd1 vccd1 vccd1 _14520_/B sky130_fd_sc_hd__and3_1
XFILLER_147_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18286_ _18286_/A vssd1 vssd1 vccd1 vccd1 _19978_/D sky130_fd_sc_hd__clkbuf_1
X_15498_ _15498_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _15498_/Y sky130_fd_sc_hd__nor2_1
X_17237_ _17135_/X _19538_/Q _17243_/S vssd1 vssd1 vccd1 vccd1 _17238_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14449_ _14450_/A _14450_/B _14448_/Y vssd1 vssd1 vccd1 vccd1 _18715_/D sky130_fd_sc_hd__o21a_1
XFILLER_128_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13743__A1 _13742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17168_ _17167_/X _19511_/Q _17177_/S vssd1 vssd1 vccd1 vccd1 _17169_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16119_ _16119_/A vssd1 vssd1 vccd1 vccd1 _19081_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17992__S _17998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09990_ _10305_/A vssd1 vssd1 vccd1 vccd1 _10064_/A sky130_fd_sc_hd__buf_2
X_17099_ _17180_/A vssd1 vssd1 vccd1 vccd1 _17199_/S sky130_fd_sc_hd__buf_4
XFILLER_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11506__B1 _09820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09804__A _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19809_ _19971_/CLK _19809_/D vssd1 vssd1 vccd1 vccd1 _19809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15799__A2 _11860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12482__A1 _12452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17232__S _17232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13760__S _13772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _15777_/A _11770_/B vssd1 vssd1 vccd1 vccd1 _12065_/B sky130_fd_sc_hd__nor2_2
XFILLER_13_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12884__B _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09355_ _09355_/A vssd1 vssd1 vccd1 vccd1 _13340_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15971__A2 _15951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09286_ _14761_/B _09245_/A _11961_/C _09313_/A vssd1 vssd1 vccd1 vccd1 _09287_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_32_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13734__A1 _13733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11745__B1 _11744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10130_ _10185_/A _10129_/X _09988_/A vssd1 vssd1 vccd1 vccd1 _10130_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17407__S _17409_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10061_ _10270_/A _10055_/X _10057_/Y _10060_/Y vssd1 vssd1 vccd1 vccd1 _10061_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16311__S _16314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13820_ _18505_/Q _13819_/X _13820_/S vssd1 vssd1 vccd1 vccd1 _13821_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13751_ _12347_/A _13746_/Y _16075_/B vssd1 vssd1 vccd1 vccd1 _13751_/X sky130_fd_sc_hd__a21o_1
X_10963_ _19137_/Q _19398_/Q _19297_/Q _19632_/Q _10962_/X _10893_/A vssd1 vssd1 vccd1
+ vccd1 _10964_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13670__A0 _18474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17142__S _17145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ _12750_/C _12701_/Y _12425_/X vssd1 vssd1 vccd1 vccd1 _12702_/Y sky130_fd_sc_hd__o21ai_1
X_16470_ _19222_/Q _13854_/X _16472_/S vssd1 vssd1 vccd1 vccd1 _16471_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13682_ _13693_/C _13681_/Y _13648_/X vssd1 vssd1 vccd1 vccd1 _13682_/Y sky130_fd_sc_hd__a21oi_2
X_10894_ _19923_/Q _19537_/Q _19987_/Q _19106_/Q _10892_/X _10893_/X vssd1 vssd1 vccd1
+ vccd1 _10895_/B sky130_fd_sc_hd__mux4_1
X_15421_ _15553_/A _15424_/A vssd1 vssd1 vccd1 vccd1 _15421_/X sky130_fd_sc_hd__or2_1
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12633_ _12756_/A _15463_/A _12613_/A vssd1 vssd1 vccd1 vccd1 _12636_/A sky130_fd_sc_hd__a21oi_1
XFILLER_70_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18140_ _18140_/A vssd1 vssd1 vccd1 vccd1 _19913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15352_ _15286_/X _15355_/B _15287_/X _15351_/X vssd1 vssd1 vccd1 vccd1 _15352_/X
+ sky130_fd_sc_hd__o211a_1
X_12564_ _12554_/A _12553_/X _12559_/Y _12563_/X vssd1 vssd1 vccd1 vccd1 _12564_/X
+ sky130_fd_sc_hd__o22a_4
XANTENNA__11984__A0 _18970_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15175__A0 _18838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14303_ _18667_/Q _18666_/Q _14306_/D vssd1 vssd1 vccd1 vccd1 _14304_/B sky130_fd_sc_hd__and3_1
XFILLER_156_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11515_ _15952_/C _12848_/B vssd1 vssd1 vccd1 vccd1 _11515_/X sky130_fd_sc_hd__and2_1
XFILLER_12_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18071_ _18845_/Q _11860_/D _18084_/S vssd1 vssd1 vccd1 vccd1 _18071_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17378__A _17424_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15283_ _15247_/X _15134_/X _14986_/X vssd1 vssd1 vccd1 vccd1 _15283_/X sky130_fd_sc_hd__o21a_1
XFILLER_145_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16282__A _16282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12495_ _12495_/A _12495_/B vssd1 vssd1 vccd1 vccd1 _12495_/Y sky130_fd_sc_hd__nor2_1
X_17022_ _17022_/A vssd1 vssd1 vccd1 vccd1 _19461_/D sky130_fd_sc_hd__clkbuf_1
X_14234_ _14234_/A _14234_/B vssd1 vssd1 vccd1 vccd1 _14236_/A sky130_fd_sc_hd__nor2_1
XFILLER_144_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11446_ _19128_/Q _19389_/Q _19288_/Q _19623_/Q _11153_/A _19385_/Q vssd1 vssd1 vccd1
+ vccd1 _11447_/B sky130_fd_sc_hd__mux4_1
XFILLER_172_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11736__B1 _11855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14165_ _14189_/A _14165_/B _14166_/B vssd1 vssd1 vccd1 vccd1 _18626_/D sky130_fd_sc_hd__nor3_1
XANTENNA__10634__S1 _10626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11377_ _11421_/A _11377_/B vssd1 vssd1 vccd1 vccd1 _11377_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ _13115_/X _18433_/Q _13116_/S vssd1 vssd1 vccd1 vccd1 _13117_/A sky130_fd_sc_hd__mux2_1
X_10328_ _19374_/Q _19709_/Q _10328_/S vssd1 vssd1 vccd1 vccd1 _10329_/B sky130_fd_sc_hd__mux2_1
XFILLER_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18973_ _18975_/CLK _18973_/D vssd1 vssd1 vccd1 vccd1 _18973_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _14095_/A _14095_/C _18608_/Q vssd1 vssd1 vccd1 vccd1 _14097_/C sky130_fd_sc_hd__a21oi_1
XFILLER_106_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _19833_/Q _17052_/X _17926_/S vssd1 vssd1 vccd1 vccd1 _17925_/A sky130_fd_sc_hd__mux2_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13047_/A _13088_/B vssd1 vssd1 vccd1 vccd1 _13047_/Y sky130_fd_sc_hd__nor2_1
X_10259_ _10266_/A _10259_/B vssd1 vssd1 vccd1 vccd1 _10259_/X sky130_fd_sc_hd__or2_1
XANTENNA__16221__S _16221_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17855_ _17855_/A vssd1 vssd1 vccd1 vccd1 _19802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16806_ _16358_/X _19370_/Q _16808_/S vssd1 vssd1 vccd1 vccd1 _16807_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17786_ _17786_/A vssd1 vssd1 vccd1 vccd1 _19771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14998_ _15353_/A vssd1 vssd1 vccd1 vccd1 _14998_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19525_ _19526_/CLK _19525_/D vssd1 vssd1 vccd1 vccd1 _19525_/Q sky130_fd_sc_hd__dfxtp_1
X_16737_ _16737_/A vssd1 vssd1 vccd1 vccd1 _19339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13949_ _13967_/A _13956_/C vssd1 vssd1 vccd1 vccd1 _13949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_5_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19456_ _19948_/CLK _19456_/D vssd1 vssd1 vccd1 vccd1 _19456_/Q sky130_fd_sc_hd__dfxtp_1
X_16668_ _16368_/X _19309_/Q _16674_/S vssd1 vssd1 vccd1 vccd1 _16669_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17987__S _17987_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18407_ _17713_/X _20033_/Q _18407_/S vssd1 vssd1 vccd1 vccd1 _18408_/A sky130_fd_sc_hd__mux2_1
X_15619_ _15619_/A vssd1 vssd1 vccd1 vccd1 _18890_/D sky130_fd_sc_hd__clkbuf_1
X_19387_ _19526_/CLK _19387_/D vssd1 vssd1 vccd1 vccd1 _19387_/Q sky130_fd_sc_hd__dfxtp_1
X_16599_ _16599_/A vssd1 vssd1 vccd1 vccd1 _19278_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15953__A2 _15951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18338_ _17716_/X _20002_/Q _18346_/S vssd1 vssd1 vccd1 vccd1 _18339_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18269_ _18269_/A vssd1 vssd1 vccd1 vccd1 _19971_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12924__S _13003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14913__A0 _15160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12225__A _12234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15469__A1 _18856_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09973_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _09973_/X sky130_fd_sc_hd__or2_1
XFILLER_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16131__S _16133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17751__A _17808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12455__A1 _11982_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12895__A _12895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10466__B1 _09539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09407_ _14227_/A _11697_/C _09407_/C vssd1 vssd1 vccd1 vccd1 _11690_/A sky130_fd_sc_hd__nor3_4
XFILLER_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09338_ _09909_/B _09909_/C vssd1 vssd1 vccd1 vccd1 _09338_/X sky130_fd_sc_hd__and2_1
XFILLER_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ _11919_/B _11951_/B vssd1 vssd1 vccd1 vccd1 _09520_/B sky130_fd_sc_hd__or2_2
XFILLER_5_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ _19131_/Q _19392_/Q _19291_/Q _19626_/Q _11171_/X _11172_/X vssd1 vssd1 vccd1
+ vccd1 _11300_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09709__A _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12280_ _12814_/S _12273_/A _12279_/X _12722_/B vssd1 vssd1 vccd1 vccd1 _12280_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11231_ _20014_/Q _19852_/Q _19261_/Q _19031_/Q _11230_/X _11108_/A vssd1 vssd1 vccd1
+ vccd1 _11232_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10354__S _10354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15837__A1_N input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11194__A1 _11095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12930__A2 _11732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _19326_/Q _19597_/Q _19821_/Q _19565_/Q _11017_/A _11015_/X vssd1 vssd1 vccd1
+ vccd1 _11162_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10113_ _19219_/Q _19810_/Q _19972_/Q _19187_/Q _09595_/A _10109_/X vssd1 vssd1 vccd1
+ vccd1 _10114_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11093_ _11441_/S vssd1 vssd1 vccd1 vccd1 _11158_/S sky130_fd_sc_hd__buf_4
X_15970_ _15978_/A _15978_/B _15970_/C vssd1 vssd1 vccd1 vccd1 _15970_/X sky130_fd_sc_hd__and3_1
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15880__A1 _09261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A io_dbus_rdata[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10044_ _09799_/A _10039_/X _10041_/Y _10043_/Y _09807_/X vssd1 vssd1 vccd1 vccd1
+ _10044_/X sky130_fd_sc_hd__o221a_1
XANTENNA__15880__B2 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14921_ _15100_/A vssd1 vssd1 vccd1 vccd1 _14922_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17640_ _17640_/A vssd1 vssd1 vccd1 vccd1 _17640_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14852_ _09289_/B _12870_/B _14957_/S vssd1 vssd1 vccd1 vccd1 _14852_/X sky130_fd_sc_hd__a21o_1
XFILLER_76_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13803_ _17039_/A vssd1 vssd1 vccd1 vccd1 _13803_/X sky130_fd_sc_hd__clkbuf_2
X_14783_ _18827_/Q _14778_/A _14782_/X _14748_/X vssd1 vssd1 vccd1 vccd1 _14784_/B
+ sky130_fd_sc_hd__a22o_1
X_17571_ _17109_/X _19690_/Q _17573_/S vssd1 vssd1 vccd1 vccd1 _17572_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13643__A0 _11748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11995_ _12285_/A vssd1 vssd1 vccd1 vccd1 _12583_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output119_A _12850_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19310_ _19581_/CLK _19310_/D vssd1 vssd1 vccd1 vccd1 _19310_/Q sky130_fd_sc_hd__dfxtp_1
X_16522_ _19244_/Q _13822_/X _16530_/S vssd1 vssd1 vccd1 vccd1 _16523_/A sky130_fd_sc_hd__mux2_1
X_13734_ _13730_/Y _13733_/X _16066_/S vssd1 vssd1 vccd1 vccd1 _13734_/X sky130_fd_sc_hd__mux2_1
X_10946_ _19201_/Q _19792_/Q _19954_/Q _19169_/Q _10907_/S _10624_/A vssd1 vssd1 vccd1
+ vccd1 _10947_/B sky130_fd_sc_hd__mux4_1
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17385__A1 _17036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19241_ _19641_/CLK _19241_/D vssd1 vssd1 vccd1 vccd1 _19241_/Q sky130_fd_sc_hd__dfxtp_1
X_16453_ _19214_/Q _13829_/X _16457_/S vssd1 vssd1 vccd1 vccd1 _16454_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13413__B _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13665_ _19014_/Q _13665_/B vssd1 vssd1 vccd1 vccd1 _13665_/X sky130_fd_sc_hd__or2_1
XANTENNA__10529__S _10529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ _19330_/Q _19601_/Q _19825_/Q _19569_/Q _10703_/A _10663_/A vssd1 vssd1 vccd1
+ vccd1 _10877_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17600__S _17606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ _12641_/A _12642_/A vssd1 vssd1 vccd1 vccd1 _12617_/B sky130_fd_sc_hd__and2b_1
X_15404_ _18851_/Q _15363_/X _15403_/X vssd1 vssd1 vccd1 vccd1 _18851_/D sky130_fd_sc_hd__o21a_1
X_16384_ _17720_/A vssd1 vssd1 vccd1 vccd1 _16384_/X sky130_fd_sc_hd__clkbuf_2
X_19172_ _19827_/CLK _19172_/D vssd1 vssd1 vccd1 vccd1 _19172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13596_ _13591_/X _13594_/Y _13623_/S vssd1 vssd1 vccd1 vccd1 _13596_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10304__S0 _09655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18123_ _18123_/A vssd1 vssd1 vccd1 vccd1 _19908_/D sky130_fd_sc_hd__clkbuf_1
X_15335_ _15381_/A _15338_/A vssd1 vssd1 vccd1 vccd1 _15335_/X sky130_fd_sc_hd__or2_1
X_12547_ _12493_/A _12519_/A _12518_/A _14886_/A vssd1 vssd1 vccd1 vccd1 _12547_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15699__A1 _18547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18054_ _18840_/Q _13563_/A _18067_/S vssd1 vssd1 vccd1 vccd1 _18054_/X sky130_fd_sc_hd__mux2_1
X_15266_ _15302_/A _15270_/A vssd1 vssd1 vccd1 vccd1 _15266_/X sky130_fd_sc_hd__or2_1
XANTENNA__09619__A _11206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ _12478_/A _12524_/C vssd1 vssd1 vccd1 vccd1 _12478_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11709__B1 _13164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17005_ _19456_/Q _17004_/X _17008_/S vssd1 vssd1 vccd1 vccd1 _17006_/A sky130_fd_sc_hd__mux2_1
X_14217_ _18644_/Q _14215_/B _14216_/Y vssd1 vssd1 vccd1 vccd1 _18644_/D sky130_fd_sc_hd__o21a_1
XFILLER_172_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11429_ _11291_/A _11419_/X _11428_/X _10078_/A _12895_/A vssd1 vssd1 vccd1 vccd1
+ _11967_/A sky130_fd_sc_hd__o32a_2
XANTENNA__10607__S1 _09607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15197_ _15197_/A vssd1 vssd1 vccd1 vccd1 _18839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16648__A0 _16339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14148_ _14153_/B _14153_/C _14102_/X vssd1 vssd1 vccd1 vccd1 _14148_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17047__S _17056_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__A _14102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14079_ _14078_/A _14078_/C _18602_/Q vssd1 vssd1 vccd1 vccd1 _14080_/C sky130_fd_sc_hd__a21oi_1
X_18956_ _18956_/CLK _18956_/D vssd1 vssd1 vccd1 vccd1 _18956_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13331__C1 _11869_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17907_ _19825_/Q _17026_/X _17915_/S vssd1 vssd1 vccd1 vccd1 _17908_/A sky130_fd_sc_hd__mux2_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16886__S _16892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18887_ _19055_/CLK _18887_/D vssd1 vssd1 vccd1 vccd1 _18887_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13882__B1 _14447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17838_ _17838_/A vssd1 vssd1 vccd1 vccd1 _19794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13634__A0 _18469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17769_ _17678_/X _19764_/Q _17771_/S vssd1 vssd1 vccd1 vccd1 _17770_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19508_ _19864_/CLK _19508_/D vssd1 vssd1 vccd1 vccd1 _19508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19439_ _19995_/CLK _19439_/D vssd1 vssd1 vccd1 vccd1 _19439_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15926__A2 _15921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11124__A _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11099__S1 _11022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9_0_clock_A clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11176__A1 _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10384__C1 _09807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09956_ _19156_/Q _19417_/Q _19316_/Q _19651_/Q _09950_/S _09824_/A vssd1 vssd1 vccd1
+ vccd1 _09957_/B sky130_fd_sc_hd__mux4_1
XFILLER_89_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10136__C1 _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09887_ _11572_/A _09887_/B vssd1 vssd1 vccd1 vccd1 _09887_/Y sky130_fd_sc_hd__nor2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _11500_/A _10799_/X _09775_/A vssd1 vssd1 vccd1 vccd1 _10800_/X sky130_fd_sc_hd__o21a_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _15758_/A _11780_/B vssd1 vssd1 vccd1 vccd1 _11817_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11100__A1 _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10731_ _19334_/Q _19605_/Q _19829_/Q _19573_/Q _11468_/S _10597_/A vssd1 vssd1 vccd1
+ vccd1 _10731_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13233__B _13368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17420__S _17420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13450_ _13448_/Y _13476_/B _12960_/A vssd1 vssd1 vccd1 vccd1 _13450_/Y sky130_fd_sc_hd__o21ai_1
X_10662_ _10662_/A vssd1 vssd1 vccd1 vccd1 _10663_/A sky130_fd_sc_hd__buf_2
XFILLER_90_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _12394_/X _12397_/Y _12400_/X vssd1 vssd1 vccd1 vccd1 _12401_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11969__A _14865_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ _13439_/A _13702_/B vssd1 vssd1 vccd1 vccd1 _13381_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16036__S _16042_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10837__S1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ _10934_/A vssd1 vssd1 vccd1 vccd1 _10824_/A sky130_fd_sc_hd__buf_2
XFILLER_167_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15120_ _15055_/S _14983_/B _15132_/S vssd1 vssd1 vccd1 vccd1 _15120_/Y sky130_fd_sc_hd__a21oi_1
X_12332_ _12297_/A _14859_/A _12331_/X vssd1 vssd1 vccd1 vccd1 _12332_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09439__A _15393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14353__A1 _14355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15051_ _15051_/A vssd1 vssd1 vccd1 vccd1 _18834_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15550__A0 _18863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12263_ _12263_/A _15254_/A vssd1 vssd1 vccd1 vccd1 _12323_/C sky130_fd_sc_hd__or2_1
XANTENNA__17656__A _17656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16560__A _16617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14002_ _14010_/A _14007_/C vssd1 vssd1 vccd1 vccd1 _14002_/Y sky130_fd_sc_hd__nor2_1
X_11214_ _11257_/A _11214_/B vssd1 vssd1 vccd1 vccd1 _11214_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12194_ _12279_/A _12393_/B _12393_/C _12186_/Y vssd1 vssd1 vccd1 vccd1 _12194_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__10914__A1 _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__S1 _11045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18810_ _18819_/CLK _18810_/D vssd1 vssd1 vccd1 vccd1 _18810_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput73 _12301_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[11] sky130_fd_sc_hd__buf_2
X_11145_ _11145_/A _11145_/B vssd1 vssd1 vccd1 vccd1 _11145_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14080__A _14088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 _12574_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[21] sky130_fd_sc_hd__buf_2
X_19790_ _19821_/CLK _19790_/D vssd1 vssd1 vccd1 vccd1 _19790_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput95 _12812_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[31] sky130_fd_sc_hd__buf_2
XANTENNA__15853__A1 _12032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15853__B2 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18741_ _18741_/CLK _18741_/D vssd1 vssd1 vccd1 vccd1 _18741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15953_ _19011_/Q _15951_/X _15952_/X vssd1 vssd1 vccd1 vccd1 _19011_/D sky130_fd_sc_hd__a21o_1
X_11076_ _19523_/Q vssd1 vssd1 vccd1 vccd1 _11077_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10027_ _10027_/A vssd1 vssd1 vccd1 vccd1 _10329_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10678__B1 _09539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14904_ _15020_/A vssd1 vssd1 vccd1 vccd1 _15113_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_1_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18672_ _18677_/CLK _18672_/D vssd1 vssd1 vccd1 vccd1 _18672_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11875__C1 _11874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15884_ _09263_/A _15875_/X _15879_/X input53/X vssd1 vssd1 vccd1 vccd1 _15885_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_154_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10773__S0 _10704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17623_ _17623_/A vssd1 vssd1 vccd1 vccd1 _19713_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09902__A _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13616__A0 _13612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14835_ _15097_/A vssd1 vssd1 vccd1 vccd1 _14835_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11890__A2 _12943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17554_ _19683_/Q vssd1 vssd1 vccd1 vccd1 _17555_/A sky130_fd_sc_hd__clkbuf_1
X_14766_ _14766_/A _14766_/B vssd1 vssd1 vccd1 vccd1 _14766_/Y sky130_fd_sc_hd__nor2_1
X_11978_ _12366_/B _11971_/Y _11977_/X _13861_/C _18519_/Q vssd1 vssd1 vccd1 vccd1
+ _13864_/B sky130_fd_sc_hd__a32o_4
XFILLER_72_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16505_ _16505_/A vssd1 vssd1 vccd1 vccd1 _19236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10929_ _10929_/A _10929_/B vssd1 vssd1 vccd1 vccd1 _10929_/Y sky130_fd_sc_hd__nor2_1
X_13717_ _19021_/Q _13717_/B vssd1 vssd1 vccd1 vccd1 _13717_/X sky130_fd_sc_hd__or2_1
X_17485_ _17485_/A vssd1 vssd1 vccd1 vccd1 _19648_/D sky130_fd_sc_hd__clkbuf_1
X_14697_ _18800_/Q _13591_/X _14705_/S vssd1 vssd1 vccd1 vccd1 _14698_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19224_ _19485_/CLK _19224_/D vssd1 vssd1 vccd1 vccd1 _19224_/Q sky130_fd_sc_hd__dfxtp_1
X_16436_ _16436_/A vssd1 vssd1 vccd1 vccd1 _19206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13648_ _13648_/A vssd1 vssd1 vccd1 vccd1 _13648_/X sky130_fd_sc_hd__buf_2
XFILLER_158_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19842_/CLK _19155_/D vssd1 vssd1 vccd1 vccd1 _19155_/Q sky130_fd_sc_hd__dfxtp_1
X_16367_ _16367_/A vssd1 vssd1 vccd1 vccd1 _19180_/D sky130_fd_sc_hd__clkbuf_1
X_13579_ _13528_/X _13577_/X _13578_/Y _13532_/X _19003_/Q vssd1 vssd1 vccd1 vccd1
+ _13579_/X sky130_fd_sc_hd__a32o_4
XANTENNA__14255__A _18653_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18106_ _18105_/X _19903_/Q _18112_/S vssd1 vssd1 vccd1 vccd1 _18107_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15318_ _15381_/A _15321_/A vssd1 vssd1 vccd1 vccd1 _15318_/X sky130_fd_sc_hd__or2_1
XFILLER_173_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19086_ _19999_/CLK _19086_/D vssd1 vssd1 vccd1 vccd1 _19086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16298_ _16691_/A _16474_/B _16298_/C vssd1 vssd1 vccd1 vccd1 _18208_/B sky130_fd_sc_hd__nand3_4
XFILLER_173_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_79_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18037_ _12956_/B _13648_/A _16069_/B vssd1 vssd1 vccd1 vccd1 _18037_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_173_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18161__S _18169_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15249_ _15544_/A vssd1 vssd1 vccd1 vccd1 _15323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11253__S1 _11045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09810_ _09950_/S vssd1 vssd1 vccd1 vccd1 _09898_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_113_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19988_ _20020_/CLK _19988_/D vssd1 vssd1 vccd1 vccd1 _19988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15844__A1 _09458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ _11487_/A vssd1 vssd1 vccd1 vccd1 _10638_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15844__B2 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18939_ _18975_/CLK _18939_/D vssd1 vssd1 vccd1 vccd1 _18939_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__11119__A _18840_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _09920_/S vssd1 vssd1 vccd1 vccd1 _09855_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10023__A _10470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12649__S _12770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14864__S _14948_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10841__B1 _10078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14165__A _14189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11397__A1 _11181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11492__S1 _10625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14335__A1 _14336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15296__C1 _15275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09939_ _09939_/A vssd1 vssd1 vccd1 vccd1 _09939_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13228__B _18849_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15724__A _16846_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ _19061_/Q _12878_/X _12879_/A _12020_/X vssd1 vssd1 vccd1 vccd1 _12950_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11321__A1 _11199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _18711_/Q _11884_/X _11865_/X _15732_/B _11900_/X vssd1 vssd1 vccd1 vccd1
+ _18711_/D sky130_fd_sc_hd__o32a_1
XFILLER_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _12881_/A vssd1 vssd1 vccd1 vccd1 _12881_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _14629_/A _14620_/B vssd1 vssd1 vccd1 vccd1 _14621_/A sky130_fd_sc_hd__and2_1
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11832_ _11813_/X _11828_/X _11830_/Y _11831_/X _19005_/Q vssd1 vssd1 vccd1 vccd1
+ _11833_/D sky130_fd_sc_hd__a32o_4
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10507__S0 _10125_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _18756_/Q _14547_/X _14550_/Y vssd1 vssd1 vccd1 vccd1 _18756_/D sky130_fd_sc_hd__o21a_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11763_ _11831_/A vssd1 vssd1 vccd1 vccd1 _13660_/A sky130_fd_sc_hd__buf_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18246__S _18252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11180__S0 _11293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _19206_/Q _19797_/Q _19959_/Q _19174_/Q _09650_/A _10049_/A vssd1 vssd1 vccd1
+ vccd1 _10715_/B sky130_fd_sc_hd__mux4_1
XFILLER_159_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13502_ _13501_/X _18455_/Q _13502_/S vssd1 vssd1 vccd1 vccd1 _13503_/A sky130_fd_sc_hd__mux2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _17183_/X _19553_/Q _17276_/S vssd1 vssd1 vccd1 vccd1 _17271_/A sky130_fd_sc_hd__mux2_1
X_14482_ _18726_/Q _14478_/B _14481_/Y vssd1 vssd1 vccd1 vccd1 _18726_/D sky130_fd_sc_hd__o21a_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11694_ _14070_/B _11683_/X _11687_/X _18630_/Q _11693_/X vssd1 vssd1 vccd1 vccd1
+ _13227_/A sky130_fd_sc_hd__a221o_2
X_16221_ _13501_/X _19127_/Q _16221_/S vssd1 vssd1 vccd1 vccd1 _16222_/A sky130_fd_sc_hd__mux2_1
X_13433_ _18818_/Q _13269_/X _12879_/X _18785_/Q _13432_/X vssd1 vssd1 vccd1 vccd1
+ _13433_/X sky130_fd_sc_hd__a221o_1
X_10645_ _19336_/Q _19607_/Q _19831_/Q _19575_/Q _10749_/S _10638_/A vssd1 vssd1 vccd1
+ vccd1 _10645_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16152_ _16208_/A vssd1 vssd1 vccd1 vccd1 _16221_/S sky130_fd_sc_hd__buf_4
XFILLER_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13364_ _17071_/A vssd1 vssd1 vccd1 vccd1 _17713_/A sky130_fd_sc_hd__clkbuf_2
X_10576_ _10223_/A _10573_/X _10575_/X vssd1 vssd1 vccd1 vccd1 _10576_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_80_clock_A _19379_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10060__A1 _11533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12315_ _12315_/A vssd1 vssd1 vccd1 vccd1 _15916_/A sky130_fd_sc_hd__clkbuf_2
X_15103_ _15517_/A _15103_/B vssd1 vssd1 vccd1 vccd1 _15103_/X sky130_fd_sc_hd__or2_1
XANTENNA__14225__D _14225_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16083_ _12939_/X _19065_/Q _16089_/S vssd1 vssd1 vccd1 vccd1 _16084_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13295_ _18570_/Q _13070_/X _13292_/X _13293_/X _13294_/X vssd1 vssd1 vccd1 vccd1
+ _13665_/B sky130_fd_sc_hd__a2111o_1
XFILLER_155_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14803__A _15954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15034_ _15032_/X _15033_/X _15041_/S vssd1 vssd1 vccd1 vccd1 _15034_/X sky130_fd_sc_hd__mux2_1
X_19911_ _19912_/CLK _19911_/D vssd1 vssd1 vccd1 vccd1 _19911_/Q sky130_fd_sc_hd__dfxtp_1
X_12246_ _12246_/A _12246_/B vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__xor2_4
XFILLER_135_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11235__S1 _11172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19842_ _19842_/CLK _19842_/D vssd1 vssd1 vccd1 vccd1 _19842_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13419__A _13439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12177_ _12080_/B _15178_/B _12209_/C _12208_/A vssd1 vssd1 vccd1 vccd1 _12178_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_150_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _11122_/X _11126_/X _11127_/X _11252_/A _11003_/X vssd1 vssd1 vccd1 vccd1
+ _11133_/B sky130_fd_sc_hd__o221a_1
X_19773_ _19935_/CLK _19773_/D vssd1 vssd1 vccd1 vccd1 _19773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16985_ _16985_/A vssd1 vssd1 vccd1 vccd1 _19449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15634__A _15690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18724_ _18724_/CLK _18724_/D vssd1 vssd1 vccd1 vccd1 _18724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11059_ _11137_/A _11052_/X _11056_/X _11058_/X vssd1 vssd1 vccd1 vccd1 _11059_/X
+ sky130_fd_sc_hd__o211a_1
X_15936_ _15936_/A _15936_/B vssd1 vssd1 vccd1 vccd1 _15936_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11312__A1 _11181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09632__A _09933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18655_ _18655_/CLK _18655_/D vssd1 vssd1 vccd1 vccd1 _18655_/Q sky130_fd_sc_hd__dfxtp_1
X_15867_ _09454_/B _15856_/X _15788_/X input48/X vssd1 vssd1 vccd1 vccd1 _16841_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17606_ _17160_/X _19706_/Q _17606_/S vssd1 vssd1 vccd1 vccd1 _17607_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14818_ _14818_/A vssd1 vssd1 vccd1 vccd1 _15368_/A sky130_fd_sc_hd__buf_2
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18586_ _18719_/CLK _18586_/D vssd1 vssd1 vccd1 vccd1 _18586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15798_ _15834_/A vssd1 vssd1 vccd1 vccd1 _15798_/X sky130_fd_sc_hd__buf_2
X_17537_ _17537_/A vssd1 vssd1 vccd1 vccd1 _19674_/D sky130_fd_sc_hd__clkbuf_1
X_14749_ _14749_/A _14749_/B _09467_/X _09454_/B vssd1 vssd1 vccd1 vccd1 _14750_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18156__S _18158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17060__S _17072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17468_ _17157_/X _19641_/Q _17470_/S vssd1 vssd1 vccd1 vccd1 _17469_/A sky130_fd_sc_hd__mux2_1
X_19207_ _20024_/CLK _19207_/D vssd1 vssd1 vccd1 vccd1 _19207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_182_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _18997_/CLK sky130_fd_sc_hd__clkbuf_16
X_16419_ _16419_/A vssd1 vssd1 vccd1 vccd1 _19198_/D sky130_fd_sc_hd__clkbuf_1
X_17399_ _17399_/A vssd1 vssd1 vccd1 vccd1 _19610_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11379__A1 _11206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19138_ _19633_/CLK _19138_/D vssd1 vssd1 vccd1 vccd1 _19138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09992__A1 _10057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19069_ _19693_/CLK _19069_/D vssd1 vssd1 vccd1 vccd1 _19069_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15514__B1 _15513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_197_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19389_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09807__A _09807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__S1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11551__A1 _09862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15817__B2 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_120_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19873_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13763__S _13772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _10859_/S vssd1 vssd1 vccd1 vccd1 _09725_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__17235__S _17243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09655_ _09655_/A vssd1 vssd1 vccd1 vccd1 _10058_/A sky130_fd_sc_hd__buf_2
XANTENNA__10511__C1 _10668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13064__A _17017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_135_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19910_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09261__B _09261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _09586_/A vssd1 vssd1 vccd1 vccd1 _11273_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12803__A1 _12316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12803__B2 _11904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__S0 _11017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_102_clock_A clkbuf_4_15_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13003__S _13003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ _19340_/Q _19611_/Q _19835_/Q _19579_/Q _10209_/S _10163_/X vssd1 vssd1 vccd1
+ vccd1 _10430_/X sky130_fd_sc_hd__mux4_1
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10361_ _19341_/Q _19612_/Q _19836_/Q _19580_/Q _10058_/A _10261_/A vssd1 vssd1 vccd1
+ vccd1 _10361_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15719__A _15719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16314__S _16314_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12100_ _18760_/Q _12069_/B _12071_/X vssd1 vssd1 vccd1 vccd1 _12108_/A sky130_fd_sc_hd__a21o_1
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13080_ _18654_/Q vssd1 vssd1 vccd1 vccd1 _14279_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10292_ _10292_/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10292_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11217__S1 _11208_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _12208_/A _12031_/B vssd1 vssd1 vccd1 vccd1 _12038_/A sky130_fd_sc_hd__nand2_1
XFILLER_105_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_1_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17145__S _17145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16770_ _16770_/A vssd1 vssd1 vccd1 vccd1 _19353_/D sky130_fd_sc_hd__clkbuf_1
X_13982_ _18568_/Q _18567_/Q _13982_/C vssd1 vssd1 vccd1 vccd1 _13984_/B sky130_fd_sc_hd__and3_1
XFILLER_101_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ _15747_/A vssd1 vssd1 vccd1 vccd1 _15745_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _18551_/Q _12877_/X _12928_/X _12930_/X _12932_/X vssd1 vssd1 vccd1 vccd1
+ _12933_/X sky130_fd_sc_hd__a2111o_2
XANTENNA_clkbuf_leaf_27_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16984__S _16986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _20026_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _15652_/A vssd1 vssd1 vccd1 vccd1 _18904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12866_/A _12866_/B _12864_/C vssd1 vssd1 vccd1 vccd1 _12865_/A sky130_fd_sc_hd__and3_2
XANTENNA__17981__A1 _17030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14603_ _14612_/A _14603_/B vssd1 vssd1 vccd1 vccd1 _14604_/A sky130_fd_sc_hd__and2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _11815_/A vssd1 vssd1 vccd1 vccd1 _11815_/X sky130_fd_sc_hd__clkbuf_4
X_18371_ _18371_/A vssd1 vssd1 vccd1 vccd1 _20016_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output101_A _12221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12795_ _18484_/Q _12010_/X _12530_/A vssd1 vssd1 vccd1 vccd1 _12795_/X sky130_fd_sc_hd__o21a_1
X_15583_ _13110_/A _18906_/Q _15589_/S vssd1 vssd1 vccd1 vccd1 _15584_/A sky130_fd_sc_hd__mux2_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17154_/X _19576_/Q _17326_/S vssd1 vssd1 vccd1 vccd1 _17323_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ _18750_/Q _14533_/X _14534_/S vssd1 vssd1 vccd1 vccd1 _14535_/A sky130_fd_sc_hd__mux2_1
X_11746_ _19011_/Q _13245_/B _11745_/Y vssd1 vssd1 vccd1 vccd1 _11746_/X sky130_fd_sc_hd__or3b_1
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17253_ _17253_/A vssd1 vssd1 vccd1 vccd1 _19545_/D sky130_fd_sc_hd__clkbuf_1
X_11677_ _14672_/B _11677_/B vssd1 vssd1 vccd1 vccd1 _11727_/A sky130_fd_sc_hd__nand2_1
X_14465_ _14507_/A vssd1 vssd1 vccd1 vccd1 _14465_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16204_ _13354_/X _19119_/Q _16206_/S vssd1 vssd1 vccd1 vccd1 _16205_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11222__A _11291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10628_ _10643_/A _10628_/B vssd1 vssd1 vccd1 vccd1 _10628_/Y sky130_fd_sc_hd__nor2_1
X_13416_ _18673_/Q _11815_/X _12887_/X _18641_/Q vssd1 vssd1 vccd1 vccd1 _13416_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17184_ _17183_/X _19516_/Q _17193_/S vssd1 vssd1 vccd1 vccd1 _17185_/A sky130_fd_sc_hd__mux2_1
X_14396_ _14398_/B _14398_/C _14395_/Y vssd1 vssd1 vccd1 vccd1 _18694_/D sky130_fd_sc_hd__o21a_1
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16135_ _16135_/A vssd1 vssd1 vccd1 vccd1 _16144_/S sky130_fd_sc_hd__buf_4
X_13347_ _18888_/Q vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__clkbuf_2
X_10559_ _10508_/A _10558_/X _09687_/A vssd1 vssd1 vccd1 vccd1 _10559_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09627__A _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16066_ _12069_/B _14562_/X _16066_/S vssd1 vssd1 vccd1 vccd1 _16066_/X sky130_fd_sc_hd__mux2_1
X_13278_ _18852_/Q _13657_/B _13458_/A vssd1 vssd1 vccd1 vccd1 _13278_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13149__A _17030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15017_ _15012_/X _15015_/X _15198_/S vssd1 vssd1 vccd1 vccd1 _15017_/X sky130_fd_sc_hd__mux2_1
X_12229_ _18462_/Q _12012_/X _13700_/A vssd1 vssd1 vccd1 vccd1 _12229_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19825_ _19957_/CLK _19825_/D vssd1 vssd1 vccd1 vccd1 _19825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16472__A1 _13857_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15364__A _15458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19756_ _20016_/CLK _19756_/D vssd1 vssd1 vccd1 vccd1 _19756_/Q sky130_fd_sc_hd__dfxtp_1
X_16968_ _16968_/A vssd1 vssd1 vccd1 vccd1 _19441_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_52_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19828_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09362__A _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18707_ _18744_/CLK _18707_/D vssd1 vssd1 vccd1 vccd1 _18707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15919_ _15053_/X _15928_/A _12118_/Y _15918_/X vssd1 vssd1 vccd1 vccd1 _18999_/D
+ sky130_fd_sc_hd__a31o_1
X_19687_ _19720_/CLK _19687_/D vssd1 vssd1 vccd1 vccd1 _19687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16899_ _16371_/X _19411_/Q _16903_/S vssd1 vssd1 vccd1 vccd1 _16900_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10195__S1 _10182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ _15517_/A vssd1 vssd1 vccd1 vccd1 _15139_/A sky130_fd_sc_hd__buf_2
XFILLER_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18638_ _18719_/CLK _18638_/D vssd1 vssd1 vccd1 vccd1 _18638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14235__B1 _15807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14786__A1 _09188_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09371_ _09394_/A vssd1 vssd1 vccd1 vccd1 _11705_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18569_ _20005_/CLK _18569_/D vssd1 vssd1 vccd1 vccd1 _18569_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15983__B1 _15928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_67_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19846_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11144__S0 _11017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__S1 _09895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12261__A2 _12837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13210__A1 _18469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10971__A _11131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09537__A _09537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14710__A1 _11724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12721__A0 _12717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09707_ _10952_/A vssd1 vssd1 vccd1 vccd1 _11500_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11827__A2 _11815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13506__B _18996_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10186__S1 _10185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10211__A _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _10057_/A vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__buf_2
XFILLER_83_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09569_ _19524_/Q vssd1 vssd1 vccd1 vccd1 _11325_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11600_ _11600_/A _11600_/B vssd1 vssd1 vccd1 vccd1 _11600_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_24_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12580_ _12522_/X _12578_/X _12579_/X vssd1 vssd1 vccd1 vccd1 _12580_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11531_ _19686_/Q _19452_/Q _18517_/Q _19782_/Q _11532_/S _09614_/X vssd1 vssd1 vccd1
+ vccd1 _11531_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14250_ _14265_/A _14250_/B vssd1 vssd1 vccd1 vccd1 _14250_/Y sky130_fd_sc_hd__nor2_1
X_11462_ _11462_/A _11462_/B _11462_/C vssd1 vssd1 vccd1 vccd1 _11604_/B sky130_fd_sc_hd__nand3_1
XFILLER_165_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _17039_/A vssd1 vssd1 vccd1 vccd1 _17681_/A sky130_fd_sc_hd__buf_2
XFILLER_99_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10413_ _10462_/A _10412_/X _09565_/A vssd1 vssd1 vccd1 vccd1 _10413_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14181_ _14189_/A _14181_/B _14182_/B vssd1 vssd1 vccd1 vccd1 _18632_/D sky130_fd_sc_hd__nor3_1
XANTENNA__15449__A _15449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11393_ _19129_/Q _19390_/Q _19289_/Q _19624_/Q _11154_/A _11107_/A vssd1 vssd1 vccd1
+ vccd1 _11393_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13132_ _13175_/A _13132_/B _13143_/B vssd1 vssd1 vccd1 vccd1 _13132_/X sky130_fd_sc_hd__or3_1
X_10344_ _10344_/A _10344_/B vssd1 vssd1 vccd1 vccd1 _10344_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09447__A _14665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input62_A io_ibus_inst[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17940_ _19840_/Q _17074_/X _17948_/S vssd1 vssd1 vccd1 vccd1 _17941_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14701__A1 _11860_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13063_ input30/X _12906_/X _13062_/X _12874_/X vssd1 vssd1 vccd1 vccd1 _17017_/A
+ sky130_fd_sc_hd__a22o_4
X_10275_ _10275_/A _19247_/Q vssd1 vssd1 vccd1 vccd1 _10275_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12014_ _18456_/Q _12012_/X _13700_/A vssd1 vssd1 vccd1 vccd1 _12014_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17871_ _17871_/A vssd1 vssd1 vccd1 vccd1 _19809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10105__B _12857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output149_A _12454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19610_ _19972_/CLK _19610_/D vssd1 vssd1 vccd1 vccd1 _19610_/Q sky130_fd_sc_hd__dfxtp_1
X_16822_ _16380_/X _19377_/Q _16830_/S vssd1 vssd1 vccd1 vccd1 _16823_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12601__A _12601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19541_ _19990_/CLK _19541_/D vssd1 vssd1 vccd1 vccd1 _19541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16753_ _16753_/A vssd1 vssd1 vccd1 vccd1 _19346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13965_ _13991_/A _13965_/B _13966_/B vssd1 vssd1 vccd1 vccd1 _18562_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15704_ _15704_/A vssd1 vssd1 vccd1 vccd1 _18928_/D sky130_fd_sc_hd__clkbuf_1
X_19472_ _20028_/CLK _19472_/D vssd1 vssd1 vccd1 vccd1 _19472_/Q sky130_fd_sc_hd__dfxtp_1
X_12916_ _18939_/Q vssd1 vssd1 vccd1 vccd1 _16474_/B sky130_fd_sc_hd__buf_4
XFILLER_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16684_ _16684_/A vssd1 vssd1 vccd1 vccd1 _19316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13896_ _12554_/A _13893_/X _12559_/Y _12563_/X _13890_/X vssd1 vssd1 vccd1 vccd1
+ _18538_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18423_ _18423_/A vssd1 vssd1 vccd1 vccd1 _20040_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15635_ _15703_/S vssd1 vssd1 vccd1 vccd1 _15644_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__12228__C1 _12556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15965__B1 _15955_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _12851_/A _12847_/B vssd1 vssd1 vccd1 vccd1 _12847_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__16219__S _16221_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14528__A _14528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _18422_/S vssd1 vssd1 vccd1 vccd1 _18363_/S sky130_fd_sc_hd__clkbuf_4
X_15566_ _15566_/A vssd1 vssd1 vccd1 vccd1 _18866_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09644__B1 _09568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12778_ _12778_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _15542_/A sky130_fd_sc_hd__or2_2
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17305_ _17305_/A vssd1 vssd1 vccd1 vccd1 _19568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14517_ _14518_/A _14518_/C _14516_/Y vssd1 vssd1 vccd1 vccd1 _18739_/D sky130_fd_sc_hd__o21a_1
X_11729_ _14670_/S _11724_/X _11728_/X vssd1 vssd1 vccd1 vccd1 _18749_/D sky130_fd_sc_hd__o21a_1
X_18285_ _17640_/X _19978_/Q _18291_/S vssd1 vssd1 vccd1 vccd1 _18286_/A sky130_fd_sc_hd__mux2_1
X_15497_ _14991_/X _15494_/Y _15496_/X _14998_/X vssd1 vssd1 vccd1 vccd1 _15500_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_159_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17236_ _17236_/A vssd1 vssd1 vccd1 vccd1 _19537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14448_ _14450_/A _14450_/B _14427_/X vssd1 vssd1 vccd1 vccd1 _14448_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ _17704_/A vssd1 vssd1 vccd1 vccd1 _17167_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12400__C1 _12188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14379_ _14399_/A _14379_/B _14384_/C vssd1 vssd1 vccd1 vccd1 _18689_/D sky130_fd_sc_hd__nor3_1
XFILLER_116_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16118_ _13250_/X _19081_/Q _16122_/S vssd1 vssd1 vccd1 vccd1 _16119_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16142__A0 _13443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15078__B _15078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17098_ _17098_/A _17098_/B _17098_/C vssd1 vssd1 vccd1 vccd1 _17180_/A sky130_fd_sc_hd__or3_4
XFILLER_115_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16049_ _13423_/X _19053_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16050_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15094__A _15094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19808_ _20002_/CLK _19808_/D vssd1 vssd1 vccd1 vccd1 _19808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13259__A1 _12956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19739_ _19997_/CLK _19739_/D vssd1 vssd1 vccd1 vccd1 _19739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11365__S0 _11124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09423_ _11716_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _11770_/B sky130_fd_sc_hd__or2_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09820__A _09820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16129__S _16133_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09354_ _09354_/A _09354_/B vssd1 vssd1 vccd1 vccd1 _09355_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15708__B1 _14529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _18973_/Q _09434_/A _09285_/C _09435_/A vssd1 vssd1 vccd1 vccd1 _11961_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_138_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18344__S _18346_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09406__A_N _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14173__A _14189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10060_ _11533_/A _10059_/X _09973_/A vssd1 vssd1 vccd1 vccd1 _10060_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15732__A _16691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13750_ _18053_/A _13750_/B vssd1 vssd1 vccd1 vccd1 _16075_/B sky130_fd_sc_hd__and2_2
X_10962_ _11023_/S vssd1 vssd1 vccd1 vccd1 _10962_/X sky130_fd_sc_hd__buf_2
XFILLER_90_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09730__A _10166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ _18783_/Q _12700_/B _12170_/X vssd1 vssd1 vccd1 vccd1 _12701_/Y sky130_fd_sc_hd__o21ai_1
X_10893_ _10893_/A vssd1 vssd1 vccd1 vccd1 _10893_/X sky130_fd_sc_hd__buf_2
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13681_ _18887_/Q _13681_/B vssd1 vssd1 vccd1 vccd1 _13681_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15420_ _15424_/A _15424_/B vssd1 vssd1 vccd1 vccd1 _15420_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12632_ _12632_/A vssd1 vssd1 vccd1 vccd1 _12756_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12563_ _12347_/X _12561_/X _12562_/Y _12350_/X vssd1 vssd1 vccd1 vccd1 _12563_/X
+ sky130_fd_sc_hd__a31o_1
X_15351_ _15381_/A _15355_/A vssd1 vssd1 vccd1 vccd1 _15351_/X sky130_fd_sc_hd__or2_1
XFILLER_156_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11514_ _11616_/A _11616_/B _11598_/A _10759_/X vssd1 vssd1 vccd1 vccd1 _11595_/C
+ sky130_fd_sc_hd__a211o_1
X_14302_ _14312_/C _14302_/B vssd1 vssd1 vccd1 vccd1 _18666_/D sky130_fd_sc_hd__nor2_1
X_18070_ _18104_/A vssd1 vssd1 vccd1 vccd1 _18084_/S sky130_fd_sc_hd__clkbuf_2
X_12494_ _12437_/A _12467_/A _12465_/A vssd1 vssd1 vccd1 vccd1 _12495_/B sky130_fd_sc_hd__a21oi_1
X_15282_ _15365_/A vssd1 vssd1 vccd1 vccd1 _15282_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17021_ _19461_/Q _17020_/X _17024_/S vssd1 vssd1 vccd1 vccd1 _17022_/A sky130_fd_sc_hd__mux2_1
X_11445_ _19320_/Q _19591_/Q _19815_/Q _19559_/Q _11154_/A _11107_/A vssd1 vssd1 vccd1
+ vccd1 _11445_/X sky130_fd_sc_hd__mux4_1
X_14233_ _18647_/Q vssd1 vssd1 vccd1 vccd1 _14234_/A sky130_fd_sc_hd__inv_2
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12933__B1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14164_ _18626_/Q _18625_/Q _14164_/C vssd1 vssd1 vccd1 vccd1 _14166_/B sky130_fd_sc_hd__and3_1
X_11376_ _19914_/Q _19528_/Q _19978_/Q _19097_/Q _11328_/X _11322_/X vssd1 vssd1 vccd1
+ vccd1 _11377_/B sky130_fd_sc_hd__mux4_2
XFILLER_125_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13115_ _17665_/A vssd1 vssd1 vccd1 vccd1 _13115_/X sky130_fd_sc_hd__clkbuf_2
X_10327_ _15964_/B vssd1 vssd1 vccd1 vccd1 _10351_/A sky130_fd_sc_hd__inv_2
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18972_ _18972_/CLK _18972_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_2
X_14095_ _14095_/A _18608_/Q _14095_/C vssd1 vssd1 vccd1 vccd1 _14097_/B sky130_fd_sc_hd__and3_1
XANTENNA__16502__S _16508_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14811__A _14811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13489__B2 _18788_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _17923_/A vssd1 vssd1 vccd1 vccd1 _19832_/D sky130_fd_sc_hd__clkbuf_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13046_/A _18872_/Q _13046_/C vssd1 vssd1 vccd1 vccd1 _13088_/B sky130_fd_sc_hd__and3_1
X_10258_ _19151_/Q _19412_/Q _19311_/Q _19646_/Q _09657_/A _09637_/A vssd1 vssd1 vccd1
+ vccd1 _10259_/B sky130_fd_sc_hd__mux4_1
XFILLER_61_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17854_ _19802_/Q _17055_/X _17854_/S vssd1 vssd1 vccd1 vccd1 _17855_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10189_ _19346_/Q _19617_/Q _19841_/Q _19585_/Q _10354_/S _10185_/X vssd1 vssd1 vccd1
+ vccd1 _10189_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16805_ _16805_/A vssd1 vssd1 vccd1 vccd1 _19369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17785_ _17700_/X _19771_/Q _17793_/S vssd1 vssd1 vccd1 vccd1 _17786_/A sky130_fd_sc_hd__mux2_1
X_14997_ _15139_/A _15055_/S _14994_/X _14996_/X vssd1 vssd1 vccd1 vccd1 _14997_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17333__S _17337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19524_ _19524_/CLK _19524_/D vssd1 vssd1 vccd1 vccd1 _19524_/Q sky130_fd_sc_hd__dfxtp_1
X_16736_ _19339_/Q _13819_/X _16736_/S vssd1 vssd1 vccd1 vccd1 _16737_/A sky130_fd_sc_hd__mux2_1
X_13948_ _13958_/D vssd1 vssd1 vccd1 vccd1 _13956_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19455_ _19947_/CLK _19455_/D vssd1 vssd1 vccd1 vccd1 _19455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16667_ _16667_/A vssd1 vssd1 vccd1 vccd1 _19308_/D sky130_fd_sc_hd__clkbuf_1
X_13879_ _13879_/A vssd1 vssd1 vccd1 vccd1 _15833_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18406_ _18406_/A vssd1 vssd1 vccd1 vccd1 _20032_/D sky130_fd_sc_hd__clkbuf_1
X_15618_ _13699_/A _18922_/Q _15622_/S vssd1 vssd1 vccd1 vccd1 _15619_/A sky130_fd_sc_hd__mux2_1
X_19386_ _19526_/CLK _19386_/D vssd1 vssd1 vccd1 vccd1 _19386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16598_ _19278_/Q _13829_/X _16602_/S vssd1 vssd1 vccd1 vccd1 _16599_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18337_ _18337_/A vssd1 vssd1 vccd1 vccd1 _18346_/S sky130_fd_sc_hd__buf_4
XFILLER_148_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15549_ _15602_/A vssd1 vssd1 vccd1 vccd1 _15567_/S sky130_fd_sc_hd__buf_2
X_18268_ _19971_/Q _17720_/A _18274_/S vssd1 vssd1 vccd1 vccd1 _18269_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_149_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17219_ _17109_/X _19530_/Q _17221_/S vssd1 vssd1 vccd1 vccd1 _17220_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14913__A1 _12715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18199_ _18199_/A vssd1 vssd1 vccd1 vccd1 _19940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10026__A _10153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09972_ _19217_/Q _19808_/Q _19970_/Q _19185_/Q _09967_/X _09612_/A vssd1 vssd1 vccd1
+ vccd1 _09973_/B sky130_fd_sc_hd__mux4_1
XANTENNA__12940__S _13003_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16418__A1 _13778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17243__S _17243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13652__A1 _18472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12895__B _12956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__A _09550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__A1 _09849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10466__B2 _18852_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09406_ _09394_/A _11777_/B _09406_/C _11699_/A vssd1 vssd1 vccd1 vccd1 _11670_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13404__A1 _13223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09337_ _09699_/A _09337_/B _09337_/C vssd1 vssd1 vccd1 vccd1 _09909_/C sky130_fd_sc_hd__and3_1
XFILLER_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13800__A _17036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _09284_/A vssd1 vssd1 vccd1 vccd1 _11663_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09199_ _09274_/A _11919_/B _09282_/D _12003_/B vssd1 vssd1 vccd1 vccd1 _11939_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ _11442_/S vssd1 vssd1 vccd1 vccd1 _11230_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11320__A _11320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17418__S _17420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _11157_/X _11159_/X _11160_/X _11145_/A _09773_/A vssd1 vssd1 vccd1 vccd1
+ _11166_/B sky130_fd_sc_hd__o221a_1
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14631__A _14648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10112_ _10112_/A vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09725__A _09725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11092_ _11153_/A vssd1 vssd1 vccd1 vccd1 _11441_/S sky130_fd_sc_hd__buf_2
XANTENNA__15446__B _15449_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14350__B _14350_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10043_ _10007_/A _10042_/X _09799_/A vssd1 vssd1 vccd1 vccd1 _10043_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_121_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14920_ _15103_/B vssd1 vssd1 vccd1 vccd1 _15100_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13891__A1 _12446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13891__B2 _12453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input25_A io_dbus_rdata[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851_ _15268_/A vssd1 vssd1 vccd1 vccd1 _14855_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11329__S0 _11328_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13802_ _13802_/A vssd1 vssd1 vccd1 vccd1 _18499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17570_ _17570_/A vssd1 vssd1 vccd1 vccd1 _19689_/D sky130_fd_sc_hd__clkbuf_1
X_14782_ _14782_/A _14782_/B _14782_/C _14782_/D vssd1 vssd1 vccd1 vccd1 _14782_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13643__A1 _13642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17909__A1 _17030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11994_ _11994_/A vssd1 vssd1 vccd1 vccd1 _11994_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_44_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16521_ _16532_/A vssd1 vssd1 vccd1 vccd1 _16530_/S sky130_fd_sc_hd__buf_4
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13733_ _13656_/X _13731_/X _13732_/Y _13660_/X _19023_/Q vssd1 vssd1 vccd1 vccd1
+ _13733_/X sky130_fd_sc_hd__a32o_2
X_10945_ _10900_/A _10944_/X _09774_/A vssd1 vssd1 vccd1 vccd1 _10945_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19240_ _19767_/CLK _19240_/D vssd1 vssd1 vccd1 vccd1 _19240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16452_ _16452_/A vssd1 vssd1 vccd1 vccd1 _19213_/D sky130_fd_sc_hd__clkbuf_1
X_13664_ _13664_/A _13672_/C vssd1 vssd1 vccd1 vccd1 _13664_/Y sky130_fd_sc_hd__xnor2_1
X_10876_ _19138_/Q _19399_/Q _19298_/Q _19633_/Q _10776_/X _10710_/A vssd1 vssd1 vccd1
+ vccd1 _10876_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15403_ _12498_/Y _15364_/X _15402_/X _15360_/X vssd1 vssd1 vccd1 vccd1 _15403_/X
+ sky130_fd_sc_hd__a211o_1
X_19171_ _20020_/CLK _19171_/D vssd1 vssd1 vccd1 vccd1 _19171_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17389__A _17411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12615_ _12642_/A _12641_/A vssd1 vssd1 vccd1 vccd1 _12617_/A sky130_fd_sc_hd__and2b_1
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16383_ _16383_/A vssd1 vssd1 vccd1 vccd1 _19185_/D sky130_fd_sc_hd__clkbuf_1
X_13595_ _13595_/A vssd1 vssd1 vccd1 vccd1 _13623_/S sky130_fd_sc_hd__buf_2
XANTENNA__10304__S1 _10185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11501__S0 _10787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18122_ _18121_/X _19908_/Q _18128_/S vssd1 vssd1 vccd1 vccd1 _18123_/A sky130_fd_sc_hd__mux2_1
X_15334_ _15338_/A _15338_/B vssd1 vssd1 vccd1 vccd1 _15334_/Y sky130_fd_sc_hd__nand2_1
X_12546_ _12546_/A vssd1 vssd1 vccd1 vccd1 _12546_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_150_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18053_ _18053_/A vssd1 vssd1 vccd1 vccd1 _18067_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_8_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15265_ _15270_/A _15270_/B vssd1 vssd1 vccd1 vccd1 _15265_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12477_ _18534_/Q _18535_/Q _12477_/C _12477_/D vssd1 vssd1 vccd1 vccd1 _12524_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__11709__A1 _18754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14244__C _14279_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ _17004_/A vssd1 vssd1 vccd1 vccd1 _17004_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_output93_A _11994_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10068__S0 _09918_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _14239_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _14216_/Y sky130_fd_sc_hd__nor2_1
X_11428_ _11421_/Y _11423_/Y _11425_/Y _11427_/Y _19526_/Q vssd1 vssd1 vccd1 vccd1
+ _11428_/X sky130_fd_sc_hd__o221a_1
XFILLER_153_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15196_ _18839_/Q _15195_/X _15480_/S vssd1 vssd1 vccd1 vccd1 _15197_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11359_ _11401_/A _11359_/B vssd1 vssd1 vccd1 vccd1 _11359_/X sky130_fd_sc_hd__or2_1
X_14147_ _18621_/Q _14143_/C _14146_/Y vssd1 vssd1 vccd1 vccd1 _18621_/D sky130_fd_sc_hd__o21a_1
XFILLER_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16232__S _16236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09635__A _09668_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14078_ _14078_/A _18602_/Q _14078_/C vssd1 vssd1 vccd1 vccd1 _14080_/B sky130_fd_sc_hd__and3_1
X_18955_ _18956_/CLK _18955_/D vssd1 vssd1 vccd1 vccd1 _18955_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11568__S0 _11553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13331__B1 _09405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17906_ _17952_/S vssd1 vssd1 vccd1 vccd1 _17915_/S sky130_fd_sc_hd__buf_2
XFILLER_112_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13029_ _19887_/Q _13209_/B vssd1 vssd1 vccd1 vccd1 _13029_/X sky130_fd_sc_hd__and2_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18886_ _18923_/CLK _18886_/D vssd1 vssd1 vccd1 vccd1 _18886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12685__A2 _15487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17837_ _19794_/Q _17030_/X _17843_/S vssd1 vssd1 vccd1 vccd1 _17838_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11893__B1 _11852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17063__S _17072_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17768_ _17768_/A vssd1 vssd1 vccd1 vccd1 _19763_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_75_clock_A clkbuf_4_12_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14831__A0 _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10299__A1_N _18856_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16719_ _19331_/Q _13794_/X _16725_/S vssd1 vssd1 vccd1 vccd1 _16720_/A sky130_fd_sc_hd__mux2_1
X_19507_ _19864_/CLK _19507_/D vssd1 vssd1 vccd1 vccd1 _19507_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17998__S _17998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17699_ _17699_/A vssd1 vssd1 vccd1 vccd1 _19738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19438_ _19641_/CLK _19438_/D vssd1 vssd1 vccd1 vccd1 _19438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19369_ _19641_/CLK _19369_/D vssd1 vssd1 vccd1 vccd1 _19369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16407__S _16413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18089__A0 _18088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15790__A2_N _15788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13766__S _13772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16142__S _16144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09545__A _11291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15311__A1 _12335_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09955_ _09946_/A _09954_/X _09837_/A vssd1 vssd1 vccd1 vccd1 _09955_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11559__S0 _11553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17762__A _17808_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ _19942_/Q _19556_/Q _20006_/Q _19125_/Q _11553_/A _09826_/A vssd1 vssd1 vccd1
+ vccd1 _09887_/B sky130_fd_sc_hd__mux4_1
XFILLER_97_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10730_ _19142_/Q _19403_/Q _19302_/Q _19637_/Q _09650_/A _10049_/A vssd1 vssd1 vccd1
+ vccd1 _10730_/X sky130_fd_sc_hd__mux4_2
XANTENNA__15378__A1 _12443_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13389__B1 _13368_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ _19335_/Q _19606_/Q _19830_/Q _19574_/Q _10586_/S _10050_/A vssd1 vssd1 vccd1
+ vccd1 _10661_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _12399_/A _12424_/C _12399_/Y _12188_/X vssd1 vssd1 vccd1 vccd1 _12400_/X
+ sky130_fd_sc_hd__a211o_1
X_13380_ _18575_/Q _13189_/X _13375_/X _13376_/X _13379_/X vssd1 vssd1 vccd1 vccd1
+ _13702_/B sky130_fd_sc_hd__a2111o_1
X_10592_ _10587_/Y _10589_/Y _10591_/Y vssd1 vssd1 vccd1 vccd1 _10592_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11969__B _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12331_ _12299_/A _12298_/A _12297_/A _14859_/A vssd1 vssd1 vccd1 vccd1 _12331_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11050__A _11050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15050_ _09425_/B _15049_/X _15127_/S vssd1 vssd1 vccd1 vccd1 _15051_/A sky130_fd_sc_hd__mux2_1
X_12262_ _12323_/B vssd1 vssd1 vccd1 vccd1 _15270_/A sky130_fd_sc_hd__buf_2
XFILLER_119_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15550__A1 _15547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11213_ _19917_/Q _19531_/Q _19981_/Q _19100_/Q _11212_/X _11208_/X vssd1 vssd1 vccd1
+ vccd1 _11214_/B sky130_fd_sc_hd__mux4_2
X_14001_ _18575_/Q _14001_/B vssd1 vssd1 vccd1 vccd1 _14007_/C sky130_fd_sc_hd__and2_1
XFILLER_141_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15457__A _15457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12193_ _12193_/A vssd1 vssd1 vccd1 vccd1 _12279_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11144_ _19919_/Q _19533_/Q _19983_/Q _19102_/Q _11017_/A _11015_/X vssd1 vssd1 vccd1
+ vccd1 _11145_/B sky130_fd_sc_hd__mux4_1
Xoutput74 _12335_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[12] sky130_fd_sc_hd__buf_2
Xoutput85 _12599_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[22] sky130_fd_sc_hd__buf_2
XFILLER_96_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput96 _12046_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[3] sky130_fd_sc_hd__buf_2
XANTENNA__13313__B1 _11687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18740_ _18741_/CLK _18740_/D vssd1 vssd1 vccd1 vccd1 _18740_/Q sky130_fd_sc_hd__dfxtp_1
X_15952_ _15966_/A _15966_/B _15952_/C vssd1 vssd1 vccd1 vccd1 _15952_/X sky130_fd_sc_hd__and3_1
X_11075_ _11283_/A _11075_/B vssd1 vssd1 vccd1 vccd1 _11075_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10026_ _10153_/A vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__buf_2
XANTENNA__10678__A1 _09849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14903_ _14902_/X _15201_/B _15032_/S vssd1 vssd1 vccd1 vccd1 _14903_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10678__B2 _18848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18671_ _18677_/CLK _18671_/D vssd1 vssd1 vccd1 vccd1 _18671_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11875__B1 _09402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ _15883_/A vssd1 vssd1 vccd1 vccd1 _15897_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output131_A _12825_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10773__S1 _10048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ _17183_/X _19713_/Q _17628_/S vssd1 vssd1 vccd1 vccd1 _17623_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14834_ _15183_/A _14983_/B vssd1 vssd1 vccd1 vccd1 _15097_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13616__A1 _13615_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12419__A2 _12413_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17553_ _17553_/A vssd1 vssd1 vccd1 vccd1 _19682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14765_ _14765_/A _14765_/B _14815_/C _14765_/D vssd1 vssd1 vccd1 vccd1 _14766_/B
+ sky130_fd_sc_hd__or4_1
X_11977_ _14744_/B _12196_/A _12050_/A vssd1 vssd1 vccd1 vccd1 _11977_/X sky130_fd_sc_hd__and3_1
XFILLER_72_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17611__S _17617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16504_ _19236_/Q _13797_/X _16508_/S vssd1 vssd1 vccd1 vccd1 _16505_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13716_ _13723_/B _13715_/Y _13700_/X vssd1 vssd1 vccd1 vccd1 _13716_/Y sky130_fd_sc_hd__a21oi_1
X_17484_ _17179_/X _19648_/Q _17492_/S vssd1 vssd1 vccd1 vccd1 _17485_/A sky130_fd_sc_hd__mux2_1
X_10928_ _19329_/Q _19600_/Q _19824_/Q _19568_/Q _10776_/A _10709_/A vssd1 vssd1 vccd1
+ vccd1 _10929_/B sky130_fd_sc_hd__mux4_1
X_14696_ _14742_/S vssd1 vssd1 vccd1 vccd1 _14705_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19223_ _19846_/CLK _19223_/D vssd1 vssd1 vccd1 vccd1 _19223_/Q sky130_fd_sc_hd__dfxtp_1
X_16435_ _19206_/Q _13803_/X _16435_/S vssd1 vssd1 vccd1 vccd1 _16436_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13647_ _13642_/A _13646_/C _13256_/B vssd1 vssd1 vccd1 vccd1 _13647_/Y sky130_fd_sc_hd__o21ai_2
X_10859_ _19363_/Q _19698_/Q _10859_/S vssd1 vssd1 vccd1 vccd1 _10859_/X sky130_fd_sc_hd__mux2_1
X_19154_ _19942_/CLK _19154_/D vssd1 vssd1 vccd1 vccd1 _19154_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16364_/X _19180_/Q _16378_/S vssd1 vssd1 vccd1 vccd1 _16367_/A sky130_fd_sc_hd__mux2_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13578_ _13589_/A _19003_/Q vssd1 vssd1 vccd1 vccd1 _13578_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18105_ _18855_/Q _13685_/X _18118_/S vssd1 vssd1 vccd1 vccd1 _18105_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15317_ _15393_/A vssd1 vssd1 vccd1 vccd1 _15381_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19085_ _19966_/CLK _19085_/D vssd1 vssd1 vccd1 vccd1 _19085_/Q sky130_fd_sc_hd__dfxtp_1
X_12529_ _18053_/A vssd1 vssd1 vccd1 vccd1 _12530_/A sky130_fd_sc_hd__clkbuf_2
X_16297_ _17634_/A vssd1 vssd1 vccd1 vccd1 _16297_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18036_ _18036_/A vssd1 vssd1 vccd1 vccd1 _19882_/D sky130_fd_sc_hd__clkbuf_1
X_15248_ _15247_/X _15192_/X _15074_/X vssd1 vssd1 vccd1 vccd1 _15248_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15179_ _15101_/X _15177_/B _14994_/X _15178_/X vssd1 vssd1 vccd1 vccd1 _15179_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11563__C1 _09807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10461__S0 _10180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16897__S _16903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19987_ _20021_/CLK _19987_/D vssd1 vssd1 vccd1 vccd1 _19987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09740_ _10793_/A vssd1 vssd1 vccd1 vccd1 _11487_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18938_ _18975_/CLK _18938_/D vssd1 vssd1 vccd1 vccd1 _18938_/Q sky130_fd_sc_hd__dfxtp_2
.ends

