VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Core
  CLASS BLOCK ;
  FOREIGN Core ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 496.000 96.970 500.000 ;
    END
  END clock
  PIN io_dbus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END io_dbus_addr[0]
  PIN io_dbus_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_dbus_addr[10]
  PIN io_dbus_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END io_dbus_addr[11]
  PIN io_dbus_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 214.240 500.000 214.840 ;
    END
  END io_dbus_addr[12]
  PIN io_dbus_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 496.000 322.370 500.000 ;
    END
  END io_dbus_addr[13]
  PIN io_dbus_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 496.000 29.350 500.000 ;
    END
  END io_dbus_addr[14]
  PIN io_dbus_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END io_dbus_addr[15]
  PIN io_dbus_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 37.440 500.000 38.040 ;
    END
  END io_dbus_addr[16]
  PIN io_dbus_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 496.000 480.150 500.000 ;
    END
  END io_dbus_addr[17]
  PIN io_dbus_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_dbus_addr[18]
  PIN io_dbus_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END io_dbus_addr[19]
  PIN io_dbus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END io_dbus_addr[1]
  PIN io_dbus_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END io_dbus_addr[20]
  PIN io_dbus_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 85.040 500.000 85.640 ;
    END
  END io_dbus_addr[21]
  PIN io_dbus_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 496.000 232.210 500.000 ;
    END
  END io_dbus_addr[22]
  PIN io_dbus_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 380.840 500.000 381.440 ;
    END
  END io_dbus_addr[23]
  PIN io_dbus_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END io_dbus_addr[24]
  PIN io_dbus_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 496.000 219.330 500.000 ;
    END
  END io_dbus_addr[25]
  PIN io_dbus_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 496.000 286.950 500.000 ;
    END
  END io_dbus_addr[26]
  PIN io_dbus_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END io_dbus_addr[27]
  PIN io_dbus_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 391.040 500.000 391.640 ;
    END
  END io_dbus_addr[28]
  PIN io_dbus_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END io_dbus_addr[29]
  PIN io_dbus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 496.000 119.510 500.000 ;
    END
  END io_dbus_addr[2]
  PIN io_dbus_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END io_dbus_addr[30]
  PIN io_dbus_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END io_dbus_addr[31]
  PIN io_dbus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 47.640 500.000 48.240 ;
    END
  END io_dbus_addr[3]
  PIN io_dbus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 476.040 500.000 476.640 ;
    END
  END io_dbus_addr[4]
  PIN io_dbus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 496.000 64.770 500.000 ;
    END
  END io_dbus_addr[5]
  PIN io_dbus_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END io_dbus_addr[6]
  PIN io_dbus_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END io_dbus_addr[7]
  PIN io_dbus_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END io_dbus_addr[8]
  PIN io_dbus_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END io_dbus_addr[9]
  PIN io_dbus_ld_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END io_dbus_ld_type[0]
  PIN io_dbus_ld_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 71.440 500.000 72.040 ;
    END
  END io_dbus_ld_type[1]
  PIN io_dbus_ld_type[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END io_dbus_ld_type[2]
  PIN io_dbus_rd_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END io_dbus_rd_en
  PIN io_dbus_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 496.000 42.230 500.000 ;
    END
  END io_dbus_rdata[0]
  PIN io_dbus_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 496.000 19.690 500.000 ;
    END
  END io_dbus_rdata[10]
  PIN io_dbus_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END io_dbus_rdata[11]
  PIN io_dbus_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 496.000 444.730 500.000 ;
    END
  END io_dbus_rdata[12]
  PIN io_dbus_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 319.640 500.000 320.240 ;
    END
  END io_dbus_rdata[13]
  PIN io_dbus_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 496.000 309.490 500.000 ;
    END
  END io_dbus_rdata[14]
  PIN io_dbus_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 496.000 399.650 500.000 ;
    END
  END io_dbus_rdata[15]
  PIN io_dbus_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END io_dbus_rdata[16]
  PIN io_dbus_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END io_dbus_rdata[17]
  PIN io_dbus_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 496.000 457.610 500.000 ;
    END
  END io_dbus_rdata[18]
  PIN io_dbus_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END io_dbus_rdata[19]
  PIN io_dbus_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END io_dbus_rdata[1]
  PIN io_dbus_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 404.640 500.000 405.240 ;
    END
  END io_dbus_rdata[20]
  PIN io_dbus_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 272.040 500.000 272.640 ;
    END
  END io_dbus_rdata[21]
  PIN io_dbus_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 496.000 467.270 500.000 ;
    END
  END io_dbus_rdata[22]
  PIN io_dbus_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 496.000 209.670 500.000 ;
    END
  END io_dbus_rdata[23]
  PIN io_dbus_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 248.240 500.000 248.840 ;
    END
  END io_dbus_rdata[24]
  PIN io_dbus_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 496.000 132.390 500.000 ;
    END
  END io_dbus_rdata[25]
  PIN io_dbus_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_dbus_rdata[26]
  PIN io_dbus_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 496.000 174.250 500.000 ;
    END
  END io_dbus_rdata[27]
  PIN io_dbus_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 343.440 500.000 344.040 ;
    END
  END io_dbus_rdata[28]
  PIN io_dbus_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END io_dbus_rdata[29]
  PIN io_dbus_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 496.000 435.070 500.000 ;
    END
  END io_dbus_rdata[2]
  PIN io_dbus_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 496.000 499.470 500.000 ;
    END
  END io_dbus_rdata[30]
  PIN io_dbus_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 496.000 187.130 500.000 ;
    END
  END io_dbus_rdata[31]
  PIN io_dbus_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END io_dbus_rdata[3]
  PIN io_dbus_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 156.440 500.000 157.040 ;
    END
  END io_dbus_rdata[4]
  PIN io_dbus_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 23.840 500.000 24.440 ;
    END
  END io_dbus_rdata[5]
  PIN io_dbus_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 496.000 299.830 500.000 ;
    END
  END io_dbus_rdata[6]
  PIN io_dbus_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 438.640 500.000 439.240 ;
    END
  END io_dbus_rdata[7]
  PIN io_dbus_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 176.840 500.000 177.440 ;
    END
  END io_dbus_rdata[8]
  PIN io_dbus_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END io_dbus_rdata[9]
  PIN io_dbus_st_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END io_dbus_st_type[0]
  PIN io_dbus_st_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 496.000 344.910 500.000 ;
    END
  END io_dbus_st_type[1]
  PIN io_dbus_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 452.240 500.000 452.840 ;
    END
  END io_dbus_valid
  PIN io_dbus_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 496.000 142.050 500.000 ;
    END
  END io_dbus_wdata[0]
  PIN io_dbus_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 309.440 500.000 310.040 ;
    END
  END io_dbus_wdata[10]
  PIN io_dbus_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END io_dbus_wdata[11]
  PIN io_dbus_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END io_dbus_wdata[12]
  PIN io_dbus_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END io_dbus_wdata[13]
  PIN io_dbus_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 496.000 412.530 500.000 ;
    END
  END io_dbus_wdata[14]
  PIN io_dbus_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_dbus_wdata[15]
  PIN io_dbus_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END io_dbus_wdata[16]
  PIN io_dbus_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END io_dbus_wdata[17]
  PIN io_dbus_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_dbus_wdata[18]
  PIN io_dbus_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 200.640 500.000 201.240 ;
    END
  END io_dbus_wdata[19]
  PIN io_dbus_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 119.040 500.000 119.640 ;
    END
  END io_dbus_wdata[1]
  PIN io_dbus_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END io_dbus_wdata[20]
  PIN io_dbus_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 496.000 196.790 500.000 ;
    END
  END io_dbus_wdata[21]
  PIN io_dbus_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END io_dbus_wdata[22]
  PIN io_dbus_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 414.840 500.000 415.440 ;
    END
  END io_dbus_wdata[23]
  PIN io_dbus_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_dbus_wdata[24]
  PIN io_dbus_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END io_dbus_wdata[25]
  PIN io_dbus_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 357.040 500.000 357.640 ;
    END
  END io_dbus_wdata[26]
  PIN io_dbus_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 0.040 500.000 0.640 ;
    END
  END io_dbus_wdata[27]
  PIN io_dbus_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 132.640 500.000 133.240 ;
    END
  END io_dbus_wdata[28]
  PIN io_dbus_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END io_dbus_wdata[29]
  PIN io_dbus_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 224.440 500.000 225.040 ;
    END
  END io_dbus_wdata[2]
  PIN io_dbus_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END io_dbus_wdata[30]
  PIN io_dbus_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END io_dbus_wdata[31]
  PIN io_dbus_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 261.840 500.000 262.440 ;
    END
  END io_dbus_wdata[3]
  PIN io_dbus_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END io_dbus_wdata[4]
  PIN io_dbus_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END io_dbus_wdata[5]
  PIN io_dbus_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 496.000 264.410 500.000 ;
    END
  END io_dbus_wdata[6]
  PIN io_dbus_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END io_dbus_wdata[7]
  PIN io_dbus_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END io_dbus_wdata[8]
  PIN io_dbus_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 462.440 500.000 463.040 ;
    END
  END io_dbus_wdata[9]
  PIN io_dbus_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END io_dbus_wr_en
  PIN io_ibus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 496.000 277.290 500.000 ;
    END
  END io_ibus_addr[0]
  PIN io_ibus_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END io_ibus_addr[10]
  PIN io_ibus_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 496.000 332.030 500.000 ;
    END
  END io_ibus_addr[11]
  PIN io_ibus_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END io_ibus_addr[12]
  PIN io_ibus_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END io_ibus_addr[13]
  PIN io_ibus_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 61.240 500.000 61.840 ;
    END
  END io_ibus_addr[14]
  PIN io_ibus_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END io_ibus_addr[15]
  PIN io_ibus_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 496.000 109.850 500.000 ;
    END
  END io_ibus_addr[16]
  PIN io_ibus_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 496.000 154.930 500.000 ;
    END
  END io_ibus_addr[17]
  PIN io_ibus_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 496.000 377.110 500.000 ;
    END
  END io_ibus_addr[18]
  PIN io_ibus_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END io_ibus_addr[19]
  PIN io_ibus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 108.840 500.000 109.440 ;
    END
  END io_ibus_addr[1]
  PIN io_ibus_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 285.640 500.000 286.240 ;
    END
  END io_ibus_addr[20]
  PIN io_ibus_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 496.000 164.590 500.000 ;
    END
  END io_ibus_addr[21]
  PIN io_ibus_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 190.440 500.000 191.040 ;
    END
  END io_ibus_addr[22]
  PIN io_ibus_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 496.000 51.890 500.000 ;
    END
  END io_ibus_addr[23]
  PIN io_ibus_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END io_ibus_addr[24]
  PIN io_ibus_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 367.240 500.000 367.840 ;
    END
  END io_ibus_addr[25]
  PIN io_ibus_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 496.000 389.990 500.000 ;
    END
  END io_ibus_addr[26]
  PIN io_ibus_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END io_ibus_addr[27]
  PIN io_ibus_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 142.840 500.000 143.440 ;
    END
  END io_ibus_addr[28]
  PIN io_ibus_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END io_ibus_addr[29]
  PIN io_ibus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 13.640 500.000 14.240 ;
    END
  END io_ibus_addr[2]
  PIN io_ibus_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 496.000 74.430 500.000 ;
    END
  END io_ibus_addr[30]
  PIN io_ibus_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END io_ibus_addr[31]
  PIN io_ibus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END io_ibus_addr[3]
  PIN io_ibus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END io_ibus_addr[4]
  PIN io_ibus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END io_ibus_addr[5]
  PIN io_ibus_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 428.440 500.000 429.040 ;
    END
  END io_ibus_addr[6]
  PIN io_ibus_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 295.840 500.000 296.440 ;
    END
  END io_ibus_addr[7]
  PIN io_ibus_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END io_ibus_addr[8]
  PIN io_ibus_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END io_ibus_addr[9]
  PIN io_ibus_inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 166.640 500.000 167.240 ;
    END
  END io_ibus_inst[0]
  PIN io_ibus_inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END io_ibus_inst[10]
  PIN io_ibus_inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END io_ibus_inst[11]
  PIN io_ibus_inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 486.240 500.000 486.840 ;
    END
  END io_ibus_inst[12]
  PIN io_ibus_inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END io_ibus_inst[13]
  PIN io_ibus_inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 496.000 489.810 500.000 ;
    END
  END io_ibus_inst[14]
  PIN io_ibus_inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END io_ibus_inst[15]
  PIN io_ibus_inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END io_ibus_inst[16]
  PIN io_ibus_inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END io_ibus_inst[17]
  PIN io_ibus_inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_ibus_inst[18]
  PIN io_ibus_inst[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END io_ibus_inst[19]
  PIN io_ibus_inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END io_ibus_inst[1]
  PIN io_ibus_inst[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_ibus_inst[20]
  PIN io_ibus_inst[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 496.000 254.750 500.000 ;
    END
  END io_ibus_inst[21]
  PIN io_ibus_inst[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END io_ibus_inst[22]
  PIN io_ibus_inst[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END io_ibus_inst[23]
  PIN io_ibus_inst[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_ibus_inst[24]
  PIN io_ibus_inst[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END io_ibus_inst[25]
  PIN io_ibus_inst[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 496.000 241.870 500.000 ;
    END
  END io_ibus_inst[26]
  PIN io_ibus_inst[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END io_ibus_inst[27]
  PIN io_ibus_inst[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 496.000 422.190 500.000 ;
    END
  END io_ibus_inst[28]
  PIN io_ibus_inst[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.240 500.000 95.840 ;
    END
  END io_ibus_inst[29]
  PIN io_ibus_inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END io_ibus_inst[2]
  PIN io_ibus_inst[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END io_ibus_inst[30]
  PIN io_ibus_inst[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END io_ibus_inst[31]
  PIN io_ibus_inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END io_ibus_inst[3]
  PIN io_ibus_inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END io_ibus_inst[4]
  PIN io_ibus_inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 333.240 500.000 333.840 ;
    END
  END io_ibus_inst[5]
  PIN io_ibus_inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END io_ibus_inst[6]
  PIN io_ibus_inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 496.000 367.450 500.000 ;
    END
  END io_ibus_inst[7]
  PIN io_ibus_inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 496.000 354.570 500.000 ;
    END
  END io_ibus_inst[8]
  PIN io_ibus_inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 496.000 6.810 500.000 ;
    END
  END io_ibus_inst[9]
  PIN io_ibus_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 496.000 87.310 500.000 ;
    END
  END io_ibus_valid
  PIN io_irq_motor_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END io_irq_motor_irq
  PIN io_irq_spi_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_irq_spi_irq
  PIN io_irq_uart_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END io_irq_uart_irq
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 238.040 500.000 238.640 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 0.070 8.540 499.490 488.200 ;
      LAYER met2 ;
        RECT 0.100 495.720 6.250 496.925 ;
        RECT 7.090 495.720 19.130 496.925 ;
        RECT 19.970 495.720 28.790 496.925 ;
        RECT 29.630 495.720 41.670 496.925 ;
        RECT 42.510 495.720 51.330 496.925 ;
        RECT 52.170 495.720 64.210 496.925 ;
        RECT 65.050 495.720 73.870 496.925 ;
        RECT 74.710 495.720 86.750 496.925 ;
        RECT 87.590 495.720 96.410 496.925 ;
        RECT 97.250 495.720 109.290 496.925 ;
        RECT 110.130 495.720 118.950 496.925 ;
        RECT 119.790 495.720 131.830 496.925 ;
        RECT 132.670 495.720 141.490 496.925 ;
        RECT 142.330 495.720 154.370 496.925 ;
        RECT 155.210 495.720 164.030 496.925 ;
        RECT 164.870 495.720 173.690 496.925 ;
        RECT 174.530 495.720 186.570 496.925 ;
        RECT 187.410 495.720 196.230 496.925 ;
        RECT 197.070 495.720 209.110 496.925 ;
        RECT 209.950 495.720 218.770 496.925 ;
        RECT 219.610 495.720 231.650 496.925 ;
        RECT 232.490 495.720 241.310 496.925 ;
        RECT 242.150 495.720 254.190 496.925 ;
        RECT 255.030 495.720 263.850 496.925 ;
        RECT 264.690 495.720 276.730 496.925 ;
        RECT 277.570 495.720 286.390 496.925 ;
        RECT 287.230 495.720 299.270 496.925 ;
        RECT 300.110 495.720 308.930 496.925 ;
        RECT 309.770 495.720 321.810 496.925 ;
        RECT 322.650 495.720 331.470 496.925 ;
        RECT 332.310 495.720 344.350 496.925 ;
        RECT 345.190 495.720 354.010 496.925 ;
        RECT 354.850 495.720 366.890 496.925 ;
        RECT 367.730 495.720 376.550 496.925 ;
        RECT 377.390 495.720 389.430 496.925 ;
        RECT 390.270 495.720 399.090 496.925 ;
        RECT 399.930 495.720 411.970 496.925 ;
        RECT 412.810 495.720 421.630 496.925 ;
        RECT 422.470 495.720 434.510 496.925 ;
        RECT 435.350 495.720 444.170 496.925 ;
        RECT 445.010 495.720 457.050 496.925 ;
        RECT 457.890 495.720 466.710 496.925 ;
        RECT 467.550 495.720 479.590 496.925 ;
        RECT 480.430 495.720 489.250 496.925 ;
        RECT 490.090 495.720 498.910 496.925 ;
        RECT 0.100 4.280 499.460 495.720 ;
        RECT 0.650 0.155 9.470 4.280 ;
        RECT 10.310 0.155 19.130 4.280 ;
        RECT 19.970 0.155 32.010 4.280 ;
        RECT 32.850 0.155 41.670 4.280 ;
        RECT 42.510 0.155 54.550 4.280 ;
        RECT 55.390 0.155 64.210 4.280 ;
        RECT 65.050 0.155 77.090 4.280 ;
        RECT 77.930 0.155 86.750 4.280 ;
        RECT 87.590 0.155 99.630 4.280 ;
        RECT 100.470 0.155 109.290 4.280 ;
        RECT 110.130 0.155 122.170 4.280 ;
        RECT 123.010 0.155 131.830 4.280 ;
        RECT 132.670 0.155 144.710 4.280 ;
        RECT 145.550 0.155 154.370 4.280 ;
        RECT 155.210 0.155 167.250 4.280 ;
        RECT 168.090 0.155 176.910 4.280 ;
        RECT 177.750 0.155 189.790 4.280 ;
        RECT 190.630 0.155 199.450 4.280 ;
        RECT 200.290 0.155 212.330 4.280 ;
        RECT 213.170 0.155 221.990 4.280 ;
        RECT 222.830 0.155 234.870 4.280 ;
        RECT 235.710 0.155 244.530 4.280 ;
        RECT 245.370 0.155 257.410 4.280 ;
        RECT 258.250 0.155 267.070 4.280 ;
        RECT 267.910 0.155 279.950 4.280 ;
        RECT 280.790 0.155 289.610 4.280 ;
        RECT 290.450 0.155 302.490 4.280 ;
        RECT 303.330 0.155 312.150 4.280 ;
        RECT 312.990 0.155 325.030 4.280 ;
        RECT 325.870 0.155 334.690 4.280 ;
        RECT 335.530 0.155 344.350 4.280 ;
        RECT 345.190 0.155 357.230 4.280 ;
        RECT 358.070 0.155 366.890 4.280 ;
        RECT 367.730 0.155 379.770 4.280 ;
        RECT 380.610 0.155 389.430 4.280 ;
        RECT 390.270 0.155 402.310 4.280 ;
        RECT 403.150 0.155 411.970 4.280 ;
        RECT 412.810 0.155 424.850 4.280 ;
        RECT 425.690 0.155 434.510 4.280 ;
        RECT 435.350 0.155 447.390 4.280 ;
        RECT 448.230 0.155 457.050 4.280 ;
        RECT 457.890 0.155 469.930 4.280 ;
        RECT 470.770 0.155 479.590 4.280 ;
        RECT 480.430 0.155 492.470 4.280 ;
        RECT 493.310 0.155 499.460 4.280 ;
      LAYER met3 ;
        RECT 4.400 496.040 496.000 496.905 ;
        RECT 4.000 487.240 496.000 496.040 ;
        RECT 4.000 485.840 495.600 487.240 ;
        RECT 4.000 483.840 496.000 485.840 ;
        RECT 4.400 482.440 496.000 483.840 ;
        RECT 4.000 477.040 496.000 482.440 ;
        RECT 4.000 475.640 495.600 477.040 ;
        RECT 4.000 473.640 496.000 475.640 ;
        RECT 4.400 472.240 496.000 473.640 ;
        RECT 4.000 463.440 496.000 472.240 ;
        RECT 4.000 462.040 495.600 463.440 ;
        RECT 4.000 460.040 496.000 462.040 ;
        RECT 4.400 458.640 496.000 460.040 ;
        RECT 4.000 453.240 496.000 458.640 ;
        RECT 4.000 451.840 495.600 453.240 ;
        RECT 4.000 449.840 496.000 451.840 ;
        RECT 4.400 448.440 496.000 449.840 ;
        RECT 4.000 439.640 496.000 448.440 ;
        RECT 4.000 438.240 495.600 439.640 ;
        RECT 4.000 436.240 496.000 438.240 ;
        RECT 4.400 434.840 496.000 436.240 ;
        RECT 4.000 429.440 496.000 434.840 ;
        RECT 4.000 428.040 495.600 429.440 ;
        RECT 4.000 426.040 496.000 428.040 ;
        RECT 4.400 424.640 496.000 426.040 ;
        RECT 4.000 415.840 496.000 424.640 ;
        RECT 4.000 414.440 495.600 415.840 ;
        RECT 4.000 412.440 496.000 414.440 ;
        RECT 4.400 411.040 496.000 412.440 ;
        RECT 4.000 405.640 496.000 411.040 ;
        RECT 4.000 404.240 495.600 405.640 ;
        RECT 4.000 402.240 496.000 404.240 ;
        RECT 4.400 400.840 496.000 402.240 ;
        RECT 4.000 392.040 496.000 400.840 ;
        RECT 4.000 390.640 495.600 392.040 ;
        RECT 4.000 388.640 496.000 390.640 ;
        RECT 4.400 387.240 496.000 388.640 ;
        RECT 4.000 381.840 496.000 387.240 ;
        RECT 4.000 380.440 495.600 381.840 ;
        RECT 4.000 378.440 496.000 380.440 ;
        RECT 4.400 377.040 496.000 378.440 ;
        RECT 4.000 368.240 496.000 377.040 ;
        RECT 4.000 366.840 495.600 368.240 ;
        RECT 4.000 364.840 496.000 366.840 ;
        RECT 4.400 363.440 496.000 364.840 ;
        RECT 4.000 358.040 496.000 363.440 ;
        RECT 4.000 356.640 495.600 358.040 ;
        RECT 4.000 354.640 496.000 356.640 ;
        RECT 4.400 353.240 496.000 354.640 ;
        RECT 4.000 344.440 496.000 353.240 ;
        RECT 4.000 343.040 495.600 344.440 ;
        RECT 4.000 341.040 496.000 343.040 ;
        RECT 4.400 339.640 496.000 341.040 ;
        RECT 4.000 334.240 496.000 339.640 ;
        RECT 4.000 332.840 495.600 334.240 ;
        RECT 4.000 330.840 496.000 332.840 ;
        RECT 4.400 329.440 496.000 330.840 ;
        RECT 4.000 320.640 496.000 329.440 ;
        RECT 4.400 319.240 495.600 320.640 ;
        RECT 4.000 310.440 496.000 319.240 ;
        RECT 4.000 309.040 495.600 310.440 ;
        RECT 4.000 307.040 496.000 309.040 ;
        RECT 4.400 305.640 496.000 307.040 ;
        RECT 4.000 296.840 496.000 305.640 ;
        RECT 4.400 295.440 495.600 296.840 ;
        RECT 4.000 286.640 496.000 295.440 ;
        RECT 4.000 285.240 495.600 286.640 ;
        RECT 4.000 283.240 496.000 285.240 ;
        RECT 4.400 281.840 496.000 283.240 ;
        RECT 4.000 273.040 496.000 281.840 ;
        RECT 4.400 271.640 495.600 273.040 ;
        RECT 4.000 262.840 496.000 271.640 ;
        RECT 4.000 261.440 495.600 262.840 ;
        RECT 4.000 259.440 496.000 261.440 ;
        RECT 4.400 258.040 496.000 259.440 ;
        RECT 4.000 249.240 496.000 258.040 ;
        RECT 4.400 247.840 495.600 249.240 ;
        RECT 4.000 239.040 496.000 247.840 ;
        RECT 4.000 237.640 495.600 239.040 ;
        RECT 4.000 235.640 496.000 237.640 ;
        RECT 4.400 234.240 496.000 235.640 ;
        RECT 4.000 225.440 496.000 234.240 ;
        RECT 4.400 224.040 495.600 225.440 ;
        RECT 4.000 215.240 496.000 224.040 ;
        RECT 4.000 213.840 495.600 215.240 ;
        RECT 4.000 211.840 496.000 213.840 ;
        RECT 4.400 210.440 496.000 211.840 ;
        RECT 4.000 201.640 496.000 210.440 ;
        RECT 4.400 200.240 495.600 201.640 ;
        RECT 4.000 191.440 496.000 200.240 ;
        RECT 4.000 190.040 495.600 191.440 ;
        RECT 4.000 188.040 496.000 190.040 ;
        RECT 4.400 186.640 496.000 188.040 ;
        RECT 4.000 177.840 496.000 186.640 ;
        RECT 4.400 176.440 495.600 177.840 ;
        RECT 4.000 167.640 496.000 176.440 ;
        RECT 4.000 166.240 495.600 167.640 ;
        RECT 4.000 164.240 496.000 166.240 ;
        RECT 4.400 162.840 496.000 164.240 ;
        RECT 4.000 157.440 496.000 162.840 ;
        RECT 4.000 156.040 495.600 157.440 ;
        RECT 4.000 154.040 496.000 156.040 ;
        RECT 4.400 152.640 496.000 154.040 ;
        RECT 4.000 143.840 496.000 152.640 ;
        RECT 4.000 142.440 495.600 143.840 ;
        RECT 4.000 140.440 496.000 142.440 ;
        RECT 4.400 139.040 496.000 140.440 ;
        RECT 4.000 133.640 496.000 139.040 ;
        RECT 4.000 132.240 495.600 133.640 ;
        RECT 4.000 130.240 496.000 132.240 ;
        RECT 4.400 128.840 496.000 130.240 ;
        RECT 4.000 120.040 496.000 128.840 ;
        RECT 4.000 118.640 495.600 120.040 ;
        RECT 4.000 116.640 496.000 118.640 ;
        RECT 4.400 115.240 496.000 116.640 ;
        RECT 4.000 109.840 496.000 115.240 ;
        RECT 4.000 108.440 495.600 109.840 ;
        RECT 4.000 106.440 496.000 108.440 ;
        RECT 4.400 105.040 496.000 106.440 ;
        RECT 4.000 96.240 496.000 105.040 ;
        RECT 4.000 94.840 495.600 96.240 ;
        RECT 4.000 92.840 496.000 94.840 ;
        RECT 4.400 91.440 496.000 92.840 ;
        RECT 4.000 86.040 496.000 91.440 ;
        RECT 4.000 84.640 495.600 86.040 ;
        RECT 4.000 82.640 496.000 84.640 ;
        RECT 4.400 81.240 496.000 82.640 ;
        RECT 4.000 72.440 496.000 81.240 ;
        RECT 4.000 71.040 495.600 72.440 ;
        RECT 4.000 69.040 496.000 71.040 ;
        RECT 4.400 67.640 496.000 69.040 ;
        RECT 4.000 62.240 496.000 67.640 ;
        RECT 4.000 60.840 495.600 62.240 ;
        RECT 4.000 58.840 496.000 60.840 ;
        RECT 4.400 57.440 496.000 58.840 ;
        RECT 4.000 48.640 496.000 57.440 ;
        RECT 4.000 47.240 495.600 48.640 ;
        RECT 4.000 45.240 496.000 47.240 ;
        RECT 4.400 43.840 496.000 45.240 ;
        RECT 4.000 38.440 496.000 43.840 ;
        RECT 4.000 37.040 495.600 38.440 ;
        RECT 4.000 35.040 496.000 37.040 ;
        RECT 4.400 33.640 496.000 35.040 ;
        RECT 4.000 24.840 496.000 33.640 ;
        RECT 4.000 23.440 495.600 24.840 ;
        RECT 4.000 21.440 496.000 23.440 ;
        RECT 4.400 20.040 496.000 21.440 ;
        RECT 4.000 14.640 496.000 20.040 ;
        RECT 4.000 13.240 495.600 14.640 ;
        RECT 4.000 11.240 496.000 13.240 ;
        RECT 4.400 9.840 496.000 11.240 ;
        RECT 4.000 1.040 496.000 9.840 ;
        RECT 4.000 0.175 495.600 1.040 ;
      LAYER met4 ;
        RECT 10.415 487.520 489.145 489.425 ;
        RECT 10.415 10.240 20.640 487.520 ;
        RECT 23.040 10.240 97.440 487.520 ;
        RECT 99.840 10.240 174.240 487.520 ;
        RECT 176.640 10.240 251.040 487.520 ;
        RECT 253.440 10.240 327.840 487.520 ;
        RECT 330.240 10.240 404.640 487.520 ;
        RECT 407.040 10.240 481.440 487.520 ;
        RECT 483.840 10.240 489.145 487.520 ;
        RECT 10.415 9.695 489.145 10.240 ;
  END
END Core
END LIBRARY

