magic
tech sky130A
magscale 1 2
timestamp 1647770261
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2128 98808 97424
<< metal2 >>
rect 3514 99200 3570 100000
rect 10598 99200 10654 100000
rect 17774 99200 17830 100000
rect 24858 99200 24914 100000
rect 32034 99200 32090 100000
rect 39210 99200 39266 100000
rect 46294 99200 46350 100000
rect 53470 99200 53526 100000
rect 60646 99200 60702 100000
rect 67730 99200 67786 100000
rect 74906 99200 74962 100000
rect 82082 99200 82138 100000
rect 89166 99200 89222 100000
rect 96342 99200 96398 100000
rect 4986 0 5042 800
rect 14922 0 14978 800
rect 24950 0 25006 800
rect 34978 0 35034 800
rect 44914 0 44970 800
rect 54942 0 54998 800
rect 64970 0 65026 800
rect 74906 0 74962 800
rect 84934 0 84990 800
rect 94962 0 95018 800
<< obsm2 >>
rect 1398 99144 3458 99362
rect 3626 99144 10542 99362
rect 10710 99144 17718 99362
rect 17886 99144 24802 99362
rect 24970 99144 31978 99362
rect 32146 99144 39154 99362
rect 39322 99144 46238 99362
rect 46406 99144 53414 99362
rect 53582 99144 60590 99362
rect 60758 99144 67674 99362
rect 67842 99144 74850 99362
rect 75018 99144 82026 99362
rect 82194 99144 89110 99362
rect 89278 99144 96286 99362
rect 96454 99144 98238 99362
rect 1398 856 98238 99144
rect 1398 800 4930 856
rect 5098 800 14866 856
rect 15034 800 24894 856
rect 25062 800 34922 856
rect 35090 800 44858 856
rect 45026 800 54886 856
rect 55054 800 64914 856
rect 65082 800 74850 856
rect 75018 800 84878 856
rect 85046 800 94906 856
rect 95074 800 98238 856
<< metal3 >>
rect 0 99016 800 99136
rect 0 97384 800 97504
rect 0 95752 800 95872
rect 99200 95344 100000 95464
rect 0 94120 800 94240
rect 0 92352 800 92472
rect 0 90720 800 90840
rect 0 89088 800 89208
rect 0 87456 800 87576
rect 99200 86232 100000 86352
rect 0 85688 800 85808
rect 0 84056 800 84176
rect 0 82424 800 82544
rect 0 80792 800 80912
rect 0 79024 800 79144
rect 0 77392 800 77512
rect 99200 77120 100000 77240
rect 0 75760 800 75880
rect 0 74128 800 74248
rect 0 72360 800 72480
rect 0 70728 800 70848
rect 0 69096 800 69216
rect 99200 68008 100000 68128
rect 0 67464 800 67584
rect 0 65696 800 65816
rect 0 64064 800 64184
rect 0 62432 800 62552
rect 0 60800 800 60920
rect 0 59032 800 59152
rect 99200 58896 100000 59016
rect 0 57400 800 57520
rect 0 55768 800 55888
rect 0 54136 800 54256
rect 0 52368 800 52488
rect 0 50736 800 50856
rect 99200 49920 100000 50040
rect 0 49104 800 49224
rect 0 47472 800 47592
rect 0 45704 800 45824
rect 0 44072 800 44192
rect 0 42440 800 42560
rect 0 40808 800 40928
rect 99200 40808 100000 40928
rect 0 39040 800 39160
rect 0 37408 800 37528
rect 0 35776 800 35896
rect 0 34144 800 34264
rect 0 32376 800 32496
rect 99200 31696 100000 31816
rect 0 30744 800 30864
rect 0 29112 800 29232
rect 0 27480 800 27600
rect 0 25712 800 25832
rect 0 24080 800 24200
rect 0 22448 800 22568
rect 99200 22584 100000 22704
rect 0 20816 800 20936
rect 0 19048 800 19168
rect 0 17416 800 17536
rect 0 15784 800 15904
rect 0 14152 800 14272
rect 99200 13472 100000 13592
rect 0 12384 800 12504
rect 0 10752 800 10872
rect 0 9120 800 9240
rect 0 7488 800 7608
rect 0 5720 800 5840
rect 99200 4496 100000 4616
rect 0 4088 800 4208
rect 0 2456 800 2576
rect 0 824 800 944
<< obsm3 >>
rect 880 98936 99200 99109
rect 800 97584 99200 98936
rect 880 97304 99200 97584
rect 800 95952 99200 97304
rect 880 95672 99200 95952
rect 800 95544 99200 95672
rect 800 95264 99120 95544
rect 800 94320 99200 95264
rect 880 94040 99200 94320
rect 800 92552 99200 94040
rect 880 92272 99200 92552
rect 800 90920 99200 92272
rect 880 90640 99200 90920
rect 800 89288 99200 90640
rect 880 89008 99200 89288
rect 800 87656 99200 89008
rect 880 87376 99200 87656
rect 800 86432 99200 87376
rect 800 86152 99120 86432
rect 800 85888 99200 86152
rect 880 85608 99200 85888
rect 800 84256 99200 85608
rect 880 83976 99200 84256
rect 800 82624 99200 83976
rect 880 82344 99200 82624
rect 800 80992 99200 82344
rect 880 80712 99200 80992
rect 800 79224 99200 80712
rect 880 78944 99200 79224
rect 800 77592 99200 78944
rect 880 77320 99200 77592
rect 880 77312 99120 77320
rect 800 77040 99120 77312
rect 800 75960 99200 77040
rect 880 75680 99200 75960
rect 800 74328 99200 75680
rect 880 74048 99200 74328
rect 800 72560 99200 74048
rect 880 72280 99200 72560
rect 800 70928 99200 72280
rect 880 70648 99200 70928
rect 800 69296 99200 70648
rect 880 69016 99200 69296
rect 800 68208 99200 69016
rect 800 67928 99120 68208
rect 800 67664 99200 67928
rect 880 67384 99200 67664
rect 800 65896 99200 67384
rect 880 65616 99200 65896
rect 800 64264 99200 65616
rect 880 63984 99200 64264
rect 800 62632 99200 63984
rect 880 62352 99200 62632
rect 800 61000 99200 62352
rect 880 60720 99200 61000
rect 800 59232 99200 60720
rect 880 59096 99200 59232
rect 880 58952 99120 59096
rect 800 58816 99120 58952
rect 800 57600 99200 58816
rect 880 57320 99200 57600
rect 800 55968 99200 57320
rect 880 55688 99200 55968
rect 800 54336 99200 55688
rect 880 54056 99200 54336
rect 800 52568 99200 54056
rect 880 52288 99200 52568
rect 800 50936 99200 52288
rect 880 50656 99200 50936
rect 800 50120 99200 50656
rect 800 49840 99120 50120
rect 800 49304 99200 49840
rect 880 49024 99200 49304
rect 800 47672 99200 49024
rect 880 47392 99200 47672
rect 800 45904 99200 47392
rect 880 45624 99200 45904
rect 800 44272 99200 45624
rect 880 43992 99200 44272
rect 800 42640 99200 43992
rect 880 42360 99200 42640
rect 800 41008 99200 42360
rect 880 40728 99120 41008
rect 800 39240 99200 40728
rect 880 38960 99200 39240
rect 800 37608 99200 38960
rect 880 37328 99200 37608
rect 800 35976 99200 37328
rect 880 35696 99200 35976
rect 800 34344 99200 35696
rect 880 34064 99200 34344
rect 800 32576 99200 34064
rect 880 32296 99200 32576
rect 800 31896 99200 32296
rect 800 31616 99120 31896
rect 800 30944 99200 31616
rect 880 30664 99200 30944
rect 800 29312 99200 30664
rect 880 29032 99200 29312
rect 800 27680 99200 29032
rect 880 27400 99200 27680
rect 800 25912 99200 27400
rect 880 25632 99200 25912
rect 800 24280 99200 25632
rect 880 24000 99200 24280
rect 800 22784 99200 24000
rect 800 22648 99120 22784
rect 880 22504 99120 22648
rect 880 22368 99200 22504
rect 800 21016 99200 22368
rect 880 20736 99200 21016
rect 800 19248 99200 20736
rect 880 18968 99200 19248
rect 800 17616 99200 18968
rect 880 17336 99200 17616
rect 800 15984 99200 17336
rect 880 15704 99200 15984
rect 800 14352 99200 15704
rect 880 14072 99200 14352
rect 800 13672 99200 14072
rect 800 13392 99120 13672
rect 800 12584 99200 13392
rect 880 12304 99200 12584
rect 800 10952 99200 12304
rect 880 10672 99200 10952
rect 800 9320 99200 10672
rect 880 9040 99200 9320
rect 800 7688 99200 9040
rect 880 7408 99200 7688
rect 800 5920 99200 7408
rect 880 5640 99200 5920
rect 800 4696 99200 5640
rect 800 4416 99120 4696
rect 800 4288 99200 4416
rect 880 4008 99200 4288
rect 800 2656 99200 4008
rect 880 2376 99200 2656
rect 800 1024 99200 2376
rect 880 851 99200 1024
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 6867 2619 19488 96661
rect 19968 2619 34848 96661
rect 35328 2619 50208 96661
rect 50688 2619 65261 96661
<< labels >>
rlabel metal2 s 3514 99200 3570 100000 6 clock
port 1 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 io_ba_match
port 2 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 io_motor_irq
port 3 nsew signal output
rlabel metal3 s 99200 4496 100000 4616 6 io_pwm_high
port 4 nsew signal output
rlabel metal3 s 99200 13472 100000 13592 6 io_pwm_low
port 5 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 io_qei_ch_a
port 6 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 io_qei_ch_b
port 7 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 io_wbs_ack_o
port 8 nsew signal output
rlabel metal2 s 17774 99200 17830 100000 6 io_wbs_data_o[0]
port 9 nsew signal output
rlabel metal3 s 99200 40808 100000 40928 6 io_wbs_data_o[10]
port 10 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 io_wbs_data_o[11]
port 11 nsew signal output
rlabel metal2 s 53470 99200 53526 100000 6 io_wbs_data_o[12]
port 12 nsew signal output
rlabel metal2 s 60646 99200 60702 100000 6 io_wbs_data_o[13]
port 13 nsew signal output
rlabel metal3 s 99200 49920 100000 50040 6 io_wbs_data_o[14]
port 14 nsew signal output
rlabel metal2 s 67730 99200 67786 100000 6 io_wbs_data_o[15]
port 15 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 io_wbs_data_o[16]
port 16 nsew signal output
rlabel metal2 s 74906 99200 74962 100000 6 io_wbs_data_o[17]
port 17 nsew signal output
rlabel metal3 s 99200 58896 100000 59016 6 io_wbs_data_o[18]
port 18 nsew signal output
rlabel metal3 s 99200 68008 100000 68128 6 io_wbs_data_o[19]
port 19 nsew signal output
rlabel metal2 s 24858 99200 24914 100000 6 io_wbs_data_o[1]
port 20 nsew signal output
rlabel metal2 s 82082 99200 82138 100000 6 io_wbs_data_o[20]
port 21 nsew signal output
rlabel metal2 s 89166 99200 89222 100000 6 io_wbs_data_o[21]
port 22 nsew signal output
rlabel metal2 s 96342 99200 96398 100000 6 io_wbs_data_o[22]
port 23 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 io_wbs_data_o[23]
port 24 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 io_wbs_data_o[24]
port 25 nsew signal output
rlabel metal3 s 99200 77120 100000 77240 6 io_wbs_data_o[25]
port 26 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 io_wbs_data_o[26]
port 27 nsew signal output
rlabel metal3 s 99200 86232 100000 86352 6 io_wbs_data_o[27]
port 28 nsew signal output
rlabel metal3 s 99200 95344 100000 95464 6 io_wbs_data_o[28]
port 29 nsew signal output
rlabel metal3 s 0 97384 800 97504 6 io_wbs_data_o[29]
port 30 nsew signal output
rlabel metal3 s 0 92352 800 92472 6 io_wbs_data_o[2]
port 31 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 io_wbs_data_o[30]
port 32 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 io_wbs_data_o[31]
port 33 nsew signal output
rlabel metal2 s 32034 99200 32090 100000 6 io_wbs_data_o[3]
port 34 nsew signal output
rlabel metal2 s 39210 99200 39266 100000 6 io_wbs_data_o[4]
port 35 nsew signal output
rlabel metal3 s 99200 22584 100000 22704 6 io_wbs_data_o[5]
port 36 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 io_wbs_data_o[6]
port 37 nsew signal output
rlabel metal3 s 0 94120 800 94240 6 io_wbs_data_o[7]
port 38 nsew signal output
rlabel metal2 s 46294 99200 46350 100000 6 io_wbs_data_o[8]
port 39 nsew signal output
rlabel metal3 s 99200 31696 100000 31816 6 io_wbs_data_o[9]
port 40 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 io_wbs_m2s_addr[0]
port 41 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 io_wbs_m2s_addr[10]
port 42 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 io_wbs_m2s_addr[11]
port 43 nsew signal input
rlabel metal3 s 0 50736 800 50856 6 io_wbs_m2s_addr[12]
port 44 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 io_wbs_m2s_addr[13]
port 45 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 io_wbs_m2s_addr[14]
port 46 nsew signal input
rlabel metal3 s 0 60800 800 60920 6 io_wbs_m2s_addr[15]
port 47 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 io_wbs_m2s_addr[1]
port 48 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 io_wbs_m2s_addr[2]
port 49 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_wbs_m2s_addr[3]
port 50 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 io_wbs_m2s_addr[4]
port 51 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 io_wbs_m2s_addr[5]
port 52 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 io_wbs_m2s_addr[6]
port 53 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 io_wbs_m2s_addr[7]
port 54 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 io_wbs_m2s_addr[8]
port 55 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 io_wbs_m2s_addr[9]
port 56 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 io_wbs_m2s_data[0]
port 57 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 io_wbs_m2s_data[10]
port 58 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 io_wbs_m2s_data[11]
port 59 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 io_wbs_m2s_data[12]
port 60 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 io_wbs_m2s_data[13]
port 61 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 io_wbs_m2s_data[14]
port 62 nsew signal input
rlabel metal3 s 0 62432 800 62552 6 io_wbs_m2s_data[15]
port 63 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 io_wbs_m2s_data[16]
port 64 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 io_wbs_m2s_data[17]
port 65 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 io_wbs_m2s_data[18]
port 66 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 io_wbs_m2s_data[19]
port 67 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 io_wbs_m2s_data[1]
port 68 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 io_wbs_m2s_data[20]
port 69 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 io_wbs_m2s_data[21]
port 70 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 io_wbs_m2s_data[22]
port 71 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 io_wbs_m2s_data[23]
port 72 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 io_wbs_m2s_data[24]
port 73 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 io_wbs_m2s_data[25]
port 74 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 io_wbs_m2s_data[26]
port 75 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 io_wbs_m2s_data[27]
port 76 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 io_wbs_m2s_data[28]
port 77 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 io_wbs_m2s_data[29]
port 78 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 io_wbs_m2s_data[2]
port 79 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 io_wbs_m2s_data[30]
port 80 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 io_wbs_m2s_data[31]
port 81 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 io_wbs_m2s_data[3]
port 82 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 io_wbs_m2s_data[4]
port 83 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 io_wbs_m2s_data[5]
port 84 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 io_wbs_m2s_data[6]
port 85 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 io_wbs_m2s_data[7]
port 86 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 io_wbs_m2s_data[8]
port 87 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 io_wbs_m2s_data[9]
port 88 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 io_wbs_m2s_sel[0]
port 89 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 io_wbs_m2s_sel[1]
port 90 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 io_wbs_m2s_sel[2]
port 91 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 io_wbs_m2s_sel[3]
port 92 nsew signal input
rlabel metal3 s 0 824 800 944 6 io_wbs_m2s_stb
port 93 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 io_wbs_m2s_we
port 94 nsew signal input
rlabel metal2 s 10598 99200 10654 100000 6 reset
port 95 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 96 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 97 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 97 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 97 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17572260
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/Motor_Top/runs/Motor_Top/results/finishing/Motor_Top.magic.gds
string GDS_START 1042594
<< end >>

