VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Core
  CLASS BLOCK ;
  FOREIGN Core ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END clock
  PIN io_dbus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 9.560 500.000 10.160 ;
    END
  END io_dbus_addr[0]
  PIN io_dbus_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 112.240 500.000 112.840 ;
    END
  END io_dbus_addr[10]
  PIN io_dbus_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 121.080 500.000 121.680 ;
    END
  END io_dbus_addr[11]
  PIN io_dbus_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 129.920 500.000 130.520 ;
    END
  END io_dbus_addr[12]
  PIN io_dbus_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 138.760 500.000 139.360 ;
    END
  END io_dbus_addr[13]
  PIN io_dbus_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 146.920 500.000 147.520 ;
    END
  END io_dbus_addr[14]
  PIN io_dbus_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 155.760 500.000 156.360 ;
    END
  END io_dbus_addr[15]
  PIN io_dbus_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 164.600 500.000 165.200 ;
    END
  END io_dbus_addr[16]
  PIN io_dbus_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 173.440 500.000 174.040 ;
    END
  END io_dbus_addr[17]
  PIN io_dbus_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 182.280 500.000 182.880 ;
    END
  END io_dbus_addr[18]
  PIN io_dbus_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 191.120 500.000 191.720 ;
    END
  END io_dbus_addr[19]
  PIN io_dbus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 24.520 500.000 25.120 ;
    END
  END io_dbus_addr[1]
  PIN io_dbus_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 199.960 500.000 200.560 ;
    END
  END io_dbus_addr[20]
  PIN io_dbus_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 208.800 500.000 209.400 ;
    END
  END io_dbus_addr[21]
  PIN io_dbus_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 217.640 500.000 218.240 ;
    END
  END io_dbus_addr[22]
  PIN io_dbus_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 225.800 500.000 226.400 ;
    END
  END io_dbus_addr[23]
  PIN io_dbus_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 234.640 500.000 235.240 ;
    END
  END io_dbus_addr[24]
  PIN io_dbus_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 243.480 500.000 244.080 ;
    END
  END io_dbus_addr[25]
  PIN io_dbus_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 252.320 500.000 252.920 ;
    END
  END io_dbus_addr[26]
  PIN io_dbus_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 261.160 500.000 261.760 ;
    END
  END io_dbus_addr[27]
  PIN io_dbus_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 270.000 500.000 270.600 ;
    END
  END io_dbus_addr[28]
  PIN io_dbus_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 278.840 500.000 279.440 ;
    END
  END io_dbus_addr[29]
  PIN io_dbus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 38.800 500.000 39.400 ;
    END
  END io_dbus_addr[2]
  PIN io_dbus_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 287.680 500.000 288.280 ;
    END
  END io_dbus_addr[30]
  PIN io_dbus_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 296.520 500.000 297.120 ;
    END
  END io_dbus_addr[31]
  PIN io_dbus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 51.040 500.000 51.640 ;
    END
  END io_dbus_addr[3]
  PIN io_dbus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 59.200 500.000 59.800 ;
    END
  END io_dbus_addr[4]
  PIN io_dbus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 68.040 500.000 68.640 ;
    END
  END io_dbus_addr[5]
  PIN io_dbus_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 76.880 500.000 77.480 ;
    END
  END io_dbus_addr[6]
  PIN io_dbus_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 85.720 500.000 86.320 ;
    END
  END io_dbus_addr[7]
  PIN io_dbus_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 94.560 500.000 95.160 ;
    END
  END io_dbus_addr[8]
  PIN io_dbus_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 103.400 500.000 104.000 ;
    END
  END io_dbus_addr[9]
  PIN io_dbus_ld_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 12.960 500.000 13.560 ;
    END
  END io_dbus_ld_type[0]
  PIN io_dbus_ld_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 27.240 500.000 27.840 ;
    END
  END io_dbus_ld_type[1]
  PIN io_dbus_ld_type[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 42.200 500.000 42.800 ;
    END
  END io_dbus_ld_type[2]
  PIN io_dbus_rd_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 1.400 500.000 2.000 ;
    END
  END io_dbus_rd_en
  PIN io_dbus_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 15.680 500.000 16.280 ;
    END
  END io_dbus_rdata[0]
  PIN io_dbus_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 114.960 500.000 115.560 ;
    END
  END io_dbus_rdata[10]
  PIN io_dbus_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 123.800 500.000 124.400 ;
    END
  END io_dbus_rdata[11]
  PIN io_dbus_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 132.640 500.000 133.240 ;
    END
  END io_dbus_rdata[12]
  PIN io_dbus_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 141.480 500.000 142.080 ;
    END
  END io_dbus_rdata[13]
  PIN io_dbus_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 150.320 500.000 150.920 ;
    END
  END io_dbus_rdata[14]
  PIN io_dbus_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 159.160 500.000 159.760 ;
    END
  END io_dbus_rdata[15]
  PIN io_dbus_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 168.000 500.000 168.600 ;
    END
  END io_dbus_rdata[16]
  PIN io_dbus_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 176.160 500.000 176.760 ;
    END
  END io_dbus_rdata[17]
  PIN io_dbus_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 185.000 500.000 185.600 ;
    END
  END io_dbus_rdata[18]
  PIN io_dbus_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 193.840 500.000 194.440 ;
    END
  END io_dbus_rdata[19]
  PIN io_dbus_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 29.960 500.000 30.560 ;
    END
  END io_dbus_rdata[1]
  PIN io_dbus_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 202.680 500.000 203.280 ;
    END
  END io_dbus_rdata[20]
  PIN io_dbus_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 211.520 500.000 212.120 ;
    END
  END io_dbus_rdata[21]
  PIN io_dbus_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 220.360 500.000 220.960 ;
    END
  END io_dbus_rdata[22]
  PIN io_dbus_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 229.200 500.000 229.800 ;
    END
  END io_dbus_rdata[23]
  PIN io_dbus_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 238.040 500.000 238.640 ;
    END
  END io_dbus_rdata[24]
  PIN io_dbus_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 246.880 500.000 247.480 ;
    END
  END io_dbus_rdata[25]
  PIN io_dbus_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 255.040 500.000 255.640 ;
    END
  END io_dbus_rdata[26]
  PIN io_dbus_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 263.880 500.000 264.480 ;
    END
  END io_dbus_rdata[27]
  PIN io_dbus_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 272.720 500.000 273.320 ;
    END
  END io_dbus_rdata[28]
  PIN io_dbus_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 281.560 500.000 282.160 ;
    END
  END io_dbus_rdata[29]
  PIN io_dbus_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.920 500.000 45.520 ;
    END
  END io_dbus_rdata[2]
  PIN io_dbus_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 290.400 500.000 291.000 ;
    END
  END io_dbus_rdata[30]
  PIN io_dbus_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 299.240 500.000 299.840 ;
    END
  END io_dbus_rdata[31]
  PIN io_dbus_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 53.760 500.000 54.360 ;
    END
  END io_dbus_rdata[3]
  PIN io_dbus_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 62.600 500.000 63.200 ;
    END
  END io_dbus_rdata[4]
  PIN io_dbus_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 71.440 500.000 72.040 ;
    END
  END io_dbus_rdata[5]
  PIN io_dbus_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 80.280 500.000 80.880 ;
    END
  END io_dbus_rdata[6]
  PIN io_dbus_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 88.440 500.000 89.040 ;
    END
  END io_dbus_rdata[7]
  PIN io_dbus_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 97.280 500.000 97.880 ;
    END
  END io_dbus_rdata[8]
  PIN io_dbus_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 106.120 500.000 106.720 ;
    END
  END io_dbus_rdata[9]
  PIN io_dbus_st_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 18.400 500.000 19.000 ;
    END
  END io_dbus_st_type[0]
  PIN io_dbus_st_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 33.360 500.000 33.960 ;
    END
  END io_dbus_st_type[1]
  PIN io_dbus_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 4.120 500.000 4.720 ;
    END
  END io_dbus_valid
  PIN io_dbus_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 21.800 500.000 22.400 ;
    END
  END io_dbus_wdata[0]
  PIN io_dbus_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 117.680 500.000 118.280 ;
    END
  END io_dbus_wdata[10]
  PIN io_dbus_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 126.520 500.000 127.120 ;
    END
  END io_dbus_wdata[11]
  PIN io_dbus_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 135.360 500.000 135.960 ;
    END
  END io_dbus_wdata[12]
  PIN io_dbus_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 144.200 500.000 144.800 ;
    END
  END io_dbus_wdata[13]
  PIN io_dbus_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 153.040 500.000 153.640 ;
    END
  END io_dbus_wdata[14]
  PIN io_dbus_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 161.880 500.000 162.480 ;
    END
  END io_dbus_wdata[15]
  PIN io_dbus_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 170.720 500.000 171.320 ;
    END
  END io_dbus_wdata[16]
  PIN io_dbus_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 179.560 500.000 180.160 ;
    END
  END io_dbus_wdata[17]
  PIN io_dbus_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 188.400 500.000 189.000 ;
    END
  END io_dbus_wdata[18]
  PIN io_dbus_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 196.560 500.000 197.160 ;
    END
  END io_dbus_wdata[19]
  PIN io_dbus_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 36.080 500.000 36.680 ;
    END
  END io_dbus_wdata[1]
  PIN io_dbus_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 205.400 500.000 206.000 ;
    END
  END io_dbus_wdata[20]
  PIN io_dbus_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 214.240 500.000 214.840 ;
    END
  END io_dbus_wdata[21]
  PIN io_dbus_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 223.080 500.000 223.680 ;
    END
  END io_dbus_wdata[22]
  PIN io_dbus_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 231.920 500.000 232.520 ;
    END
  END io_dbus_wdata[23]
  PIN io_dbus_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 240.760 500.000 241.360 ;
    END
  END io_dbus_wdata[24]
  PIN io_dbus_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 249.600 500.000 250.200 ;
    END
  END io_dbus_wdata[25]
  PIN io_dbus_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 258.440 500.000 259.040 ;
    END
  END io_dbus_wdata[26]
  PIN io_dbus_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 267.280 500.000 267.880 ;
    END
  END io_dbus_wdata[27]
  PIN io_dbus_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 276.120 500.000 276.720 ;
    END
  END io_dbus_wdata[28]
  PIN io_dbus_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 284.280 500.000 284.880 ;
    END
  END io_dbus_wdata[29]
  PIN io_dbus_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 47.640 500.000 48.240 ;
    END
  END io_dbus_wdata[2]
  PIN io_dbus_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 293.120 500.000 293.720 ;
    END
  END io_dbus_wdata[30]
  PIN io_dbus_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 301.960 500.000 302.560 ;
    END
  END io_dbus_wdata[31]
  PIN io_dbus_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 56.480 500.000 57.080 ;
    END
  END io_dbus_wdata[3]
  PIN io_dbus_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 65.320 500.000 65.920 ;
    END
  END io_dbus_wdata[4]
  PIN io_dbus_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 74.160 500.000 74.760 ;
    END
  END io_dbus_wdata[5]
  PIN io_dbus_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 83.000 500.000 83.600 ;
    END
  END io_dbus_wdata[6]
  PIN io_dbus_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 91.840 500.000 92.440 ;
    END
  END io_dbus_wdata[7]
  PIN io_dbus_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 100.680 500.000 101.280 ;
    END
  END io_dbus_wdata[8]
  PIN io_dbus_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 109.520 500.000 110.120 ;
    END
  END io_dbus_wdata[9]
  PIN io_dbus_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 6.840 500.000 7.440 ;
    END
  END io_dbus_wr_en
  PIN io_ibus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 308.080 500.000 308.680 ;
    END
  END io_ibus_addr[0]
  PIN io_ibus_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 366.560 500.000 367.160 ;
    END
  END io_ibus_addr[10]
  PIN io_ibus_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 372.000 500.000 372.600 ;
    END
  END io_ibus_addr[11]
  PIN io_ibus_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 378.120 500.000 378.720 ;
    END
  END io_ibus_addr[12]
  PIN io_ibus_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 384.240 500.000 384.840 ;
    END
  END io_ibus_addr[13]
  PIN io_ibus_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 389.680 500.000 390.280 ;
    END
  END io_ibus_addr[14]
  PIN io_ibus_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 395.800 500.000 396.400 ;
    END
  END io_ibus_addr[15]
  PIN io_ibus_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 401.240 500.000 401.840 ;
    END
  END io_ibus_addr[16]
  PIN io_ibus_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 407.360 500.000 407.960 ;
    END
  END io_ibus_addr[17]
  PIN io_ibus_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 413.480 500.000 414.080 ;
    END
  END io_ibus_addr[18]
  PIN io_ibus_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 418.920 500.000 419.520 ;
    END
  END io_ibus_addr[19]
  PIN io_ibus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 313.520 500.000 314.120 ;
    END
  END io_ibus_addr[1]
  PIN io_ibus_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 425.040 500.000 425.640 ;
    END
  END io_ibus_addr[20]
  PIN io_ibus_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 430.480 500.000 431.080 ;
    END
  END io_ibus_addr[21]
  PIN io_ibus_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 436.600 500.000 437.200 ;
    END
  END io_ibus_addr[22]
  PIN io_ibus_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 442.720 500.000 443.320 ;
    END
  END io_ibus_addr[23]
  PIN io_ibus_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 448.160 500.000 448.760 ;
    END
  END io_ibus_addr[24]
  PIN io_ibus_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 454.280 500.000 454.880 ;
    END
  END io_ibus_addr[25]
  PIN io_ibus_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 459.720 500.000 460.320 ;
    END
  END io_ibus_addr[26]
  PIN io_ibus_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 465.840 500.000 466.440 ;
    END
  END io_ibus_addr[27]
  PIN io_ibus_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 471.960 500.000 472.560 ;
    END
  END io_ibus_addr[28]
  PIN io_ibus_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 477.400 500.000 478.000 ;
    END
  END io_ibus_addr[29]
  PIN io_ibus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 319.640 500.000 320.240 ;
    END
  END io_ibus_addr[2]
  PIN io_ibus_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 483.520 500.000 484.120 ;
    END
  END io_ibus_addr[30]
  PIN io_ibus_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 488.960 500.000 489.560 ;
    END
  END io_ibus_addr[31]
  PIN io_ibus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 325.760 500.000 326.360 ;
    END
  END io_ibus_addr[3]
  PIN io_ibus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 331.200 500.000 331.800 ;
    END
  END io_ibus_addr[4]
  PIN io_ibus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 337.320 500.000 337.920 ;
    END
  END io_ibus_addr[5]
  PIN io_ibus_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 342.760 500.000 343.360 ;
    END
  END io_ibus_addr[6]
  PIN io_ibus_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 348.880 500.000 349.480 ;
    END
  END io_ibus_addr[7]
  PIN io_ibus_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 355.000 500.000 355.600 ;
    END
  END io_ibus_addr[8]
  PIN io_ibus_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 360.440 500.000 361.040 ;
    END
  END io_ibus_addr[9]
  PIN io_ibus_inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 310.800 500.000 311.400 ;
    END
  END io_ibus_inst[0]
  PIN io_ibus_inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 369.280 500.000 369.880 ;
    END
  END io_ibus_inst[10]
  PIN io_ibus_inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 375.400 500.000 376.000 ;
    END
  END io_ibus_inst[11]
  PIN io_ibus_inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 380.840 500.000 381.440 ;
    END
  END io_ibus_inst[12]
  PIN io_ibus_inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 386.960 500.000 387.560 ;
    END
  END io_ibus_inst[13]
  PIN io_ibus_inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 392.400 500.000 393.000 ;
    END
  END io_ibus_inst[14]
  PIN io_ibus_inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 398.520 500.000 399.120 ;
    END
  END io_ibus_inst[15]
  PIN io_ibus_inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 404.640 500.000 405.240 ;
    END
  END io_ibus_inst[16]
  PIN io_ibus_inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 410.080 500.000 410.680 ;
    END
  END io_ibus_inst[17]
  PIN io_ibus_inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 416.200 500.000 416.800 ;
    END
  END io_ibus_inst[18]
  PIN io_ibus_inst[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 421.640 500.000 422.240 ;
    END
  END io_ibus_inst[19]
  PIN io_ibus_inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 316.920 500.000 317.520 ;
    END
  END io_ibus_inst[1]
  PIN io_ibus_inst[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 427.760 500.000 428.360 ;
    END
  END io_ibus_inst[20]
  PIN io_ibus_inst[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 433.880 500.000 434.480 ;
    END
  END io_ibus_inst[21]
  PIN io_ibus_inst[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 439.320 500.000 439.920 ;
    END
  END io_ibus_inst[22]
  PIN io_ibus_inst[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 445.440 500.000 446.040 ;
    END
  END io_ibus_inst[23]
  PIN io_ibus_inst[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 450.880 500.000 451.480 ;
    END
  END io_ibus_inst[24]
  PIN io_ibus_inst[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 457.000 500.000 457.600 ;
    END
  END io_ibus_inst[25]
  PIN io_ibus_inst[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 463.120 500.000 463.720 ;
    END
  END io_ibus_inst[26]
  PIN io_ibus_inst[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 468.560 500.000 469.160 ;
    END
  END io_ibus_inst[27]
  PIN io_ibus_inst[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 474.680 500.000 475.280 ;
    END
  END io_ibus_inst[28]
  PIN io_ibus_inst[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 480.120 500.000 480.720 ;
    END
  END io_ibus_inst[29]
  PIN io_ibus_inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 322.360 500.000 322.960 ;
    END
  END io_ibus_inst[2]
  PIN io_ibus_inst[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 486.240 500.000 486.840 ;
    END
  END io_ibus_inst[30]
  PIN io_ibus_inst[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 492.360 500.000 492.960 ;
    END
  END io_ibus_inst[31]
  PIN io_ibus_inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 328.480 500.000 329.080 ;
    END
  END io_ibus_inst[3]
  PIN io_ibus_inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 334.600 500.000 335.200 ;
    END
  END io_ibus_inst[4]
  PIN io_ibus_inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.040 500.000 340.640 ;
    END
  END io_ibus_inst[5]
  PIN io_ibus_inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 346.160 500.000 346.760 ;
    END
  END io_ibus_inst[6]
  PIN io_ibus_inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 351.600 500.000 352.200 ;
    END
  END io_ibus_inst[7]
  PIN io_ibus_inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 357.720 500.000 358.320 ;
    END
  END io_ibus_inst[8]
  PIN io_ibus_inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 363.160 500.000 363.760 ;
    END
  END io_ibus_inst[9]
  PIN io_ibus_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 305.360 500.000 305.960 ;
    END
  END io_ibus_valid
  PIN io_irq_motor_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 496.000 250.150 500.000 ;
    END
  END io_irq_motor_irq
  PIN io_irq_spi_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 495.080 500.000 495.680 ;
    END
  END io_irq_spi_irq
  PIN io_irq_uart_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 497.800 500.000 498.400 ;
    END
  END io_irq_uart_irq
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 485.465 494.230 487.070 ;
        RECT 5.330 480.025 494.230 482.855 ;
        RECT 5.330 474.585 494.230 477.415 ;
        RECT 5.330 469.145 494.230 471.975 ;
        RECT 5.330 463.705 494.230 466.535 ;
        RECT 5.330 458.265 494.230 461.095 ;
        RECT 5.330 452.825 494.230 455.655 ;
        RECT 5.330 447.385 494.230 450.215 ;
        RECT 5.330 441.945 494.230 444.775 ;
        RECT 5.330 436.505 494.230 439.335 ;
        RECT 5.330 431.065 494.230 433.895 ;
        RECT 5.330 425.625 494.230 428.455 ;
        RECT 5.330 420.185 494.230 423.015 ;
        RECT 5.330 414.745 494.230 417.575 ;
        RECT 5.330 409.305 494.230 412.135 ;
        RECT 5.330 403.865 494.230 406.695 ;
        RECT 5.330 398.425 494.230 401.255 ;
        RECT 5.330 392.985 494.230 395.815 ;
        RECT 5.330 387.545 494.230 390.375 ;
        RECT 5.330 382.105 494.230 384.935 ;
        RECT 5.330 376.665 494.230 379.495 ;
        RECT 5.330 371.225 494.230 374.055 ;
        RECT 5.330 365.785 494.230 368.615 ;
        RECT 5.330 360.345 494.230 363.175 ;
        RECT 5.330 354.905 494.230 357.735 ;
        RECT 5.330 349.465 494.230 352.295 ;
        RECT 5.330 344.025 494.230 346.855 ;
        RECT 5.330 338.585 494.230 341.415 ;
        RECT 5.330 333.145 494.230 335.975 ;
        RECT 5.330 327.705 494.230 330.535 ;
        RECT 5.330 322.265 494.230 325.095 ;
        RECT 5.330 316.825 494.230 319.655 ;
        RECT 5.330 311.385 494.230 314.215 ;
        RECT 5.330 305.945 494.230 308.775 ;
        RECT 5.330 300.505 494.230 303.335 ;
        RECT 5.330 295.065 494.230 297.895 ;
        RECT 5.330 289.625 494.230 292.455 ;
        RECT 5.330 284.185 494.230 287.015 ;
        RECT 5.330 278.745 494.230 281.575 ;
        RECT 5.330 273.305 494.230 276.135 ;
        RECT 5.330 267.865 494.230 270.695 ;
        RECT 5.330 262.425 494.230 265.255 ;
        RECT 5.330 256.985 494.230 259.815 ;
        RECT 5.330 251.545 494.230 254.375 ;
        RECT 5.330 246.105 494.230 248.935 ;
        RECT 5.330 240.665 494.230 243.495 ;
        RECT 5.330 235.225 494.230 238.055 ;
        RECT 5.330 229.785 494.230 232.615 ;
        RECT 5.330 224.345 494.230 227.175 ;
        RECT 5.330 218.905 494.230 221.735 ;
        RECT 5.330 213.465 494.230 216.295 ;
        RECT 5.330 208.025 494.230 210.855 ;
        RECT 5.330 202.585 494.230 205.415 ;
        RECT 5.330 197.145 494.230 199.975 ;
        RECT 5.330 191.705 494.230 194.535 ;
        RECT 5.330 186.265 494.230 189.095 ;
        RECT 5.330 180.825 494.230 183.655 ;
        RECT 5.330 175.385 494.230 178.215 ;
        RECT 5.330 169.945 494.230 172.775 ;
        RECT 5.330 164.505 494.230 167.335 ;
        RECT 5.330 159.065 494.230 161.895 ;
        RECT 5.330 153.625 494.230 156.455 ;
        RECT 5.330 148.185 494.230 151.015 ;
        RECT 5.330 142.745 494.230 145.575 ;
        RECT 5.330 137.305 494.230 140.135 ;
        RECT 5.330 131.865 494.230 134.695 ;
        RECT 5.330 126.425 494.230 129.255 ;
        RECT 5.330 120.985 494.230 123.815 ;
        RECT 5.330 115.545 494.230 118.375 ;
        RECT 5.330 110.105 494.230 112.935 ;
        RECT 5.330 104.665 494.230 107.495 ;
        RECT 5.330 99.225 494.230 102.055 ;
        RECT 5.330 93.785 494.230 96.615 ;
        RECT 5.330 88.345 494.230 91.175 ;
        RECT 5.330 82.905 494.230 85.735 ;
        RECT 5.330 77.465 494.230 80.295 ;
        RECT 5.330 72.025 494.230 74.855 ;
        RECT 5.330 66.585 494.230 69.415 ;
        RECT 5.330 61.145 494.230 63.975 ;
        RECT 5.330 55.705 494.230 58.535 ;
        RECT 5.330 50.265 494.230 53.095 ;
        RECT 5.330 44.825 494.230 47.655 ;
        RECT 5.330 39.385 494.230 42.215 ;
        RECT 5.330 33.945 494.230 36.775 ;
        RECT 5.330 28.505 494.230 31.335 ;
        RECT 5.330 23.065 494.230 25.895 ;
        RECT 5.330 17.625 494.230 20.455 ;
        RECT 5.330 12.185 494.230 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.240 499.950 488.540 ;
      LAYER met2 ;
        RECT 7.000 495.720 249.590 498.285 ;
        RECT 250.430 495.720 499.930 498.285 ;
        RECT 7.000 4.280 499.930 495.720 ;
        RECT 7.000 1.515 124.470 4.280 ;
        RECT 125.310 1.515 374.250 4.280 ;
        RECT 375.090 1.515 499.930 4.280 ;
      LAYER met3 ;
        RECT 15.705 497.400 495.600 498.265 ;
        RECT 15.705 496.080 499.955 497.400 ;
        RECT 15.705 494.680 495.600 496.080 ;
        RECT 15.705 493.360 499.955 494.680 ;
        RECT 15.705 491.960 495.600 493.360 ;
        RECT 15.705 489.960 499.955 491.960 ;
        RECT 15.705 488.560 495.600 489.960 ;
        RECT 15.705 487.240 499.955 488.560 ;
        RECT 15.705 485.840 495.600 487.240 ;
        RECT 15.705 484.520 499.955 485.840 ;
        RECT 15.705 483.120 495.600 484.520 ;
        RECT 15.705 481.120 499.955 483.120 ;
        RECT 15.705 479.720 495.600 481.120 ;
        RECT 15.705 478.400 499.955 479.720 ;
        RECT 15.705 477.000 495.600 478.400 ;
        RECT 15.705 475.680 499.955 477.000 ;
        RECT 15.705 474.280 495.600 475.680 ;
        RECT 15.705 472.960 499.955 474.280 ;
        RECT 15.705 471.560 495.600 472.960 ;
        RECT 15.705 469.560 499.955 471.560 ;
        RECT 15.705 468.160 495.600 469.560 ;
        RECT 15.705 466.840 499.955 468.160 ;
        RECT 15.705 465.440 495.600 466.840 ;
        RECT 15.705 464.120 499.955 465.440 ;
        RECT 15.705 462.720 495.600 464.120 ;
        RECT 15.705 460.720 499.955 462.720 ;
        RECT 15.705 459.320 495.600 460.720 ;
        RECT 15.705 458.000 499.955 459.320 ;
        RECT 15.705 456.600 495.600 458.000 ;
        RECT 15.705 455.280 499.955 456.600 ;
        RECT 15.705 453.880 495.600 455.280 ;
        RECT 15.705 451.880 499.955 453.880 ;
        RECT 15.705 450.480 495.600 451.880 ;
        RECT 15.705 449.160 499.955 450.480 ;
        RECT 15.705 447.760 495.600 449.160 ;
        RECT 15.705 446.440 499.955 447.760 ;
        RECT 15.705 445.040 495.600 446.440 ;
        RECT 15.705 443.720 499.955 445.040 ;
        RECT 15.705 442.320 495.600 443.720 ;
        RECT 15.705 440.320 499.955 442.320 ;
        RECT 15.705 438.920 495.600 440.320 ;
        RECT 15.705 437.600 499.955 438.920 ;
        RECT 15.705 436.200 495.600 437.600 ;
        RECT 15.705 434.880 499.955 436.200 ;
        RECT 15.705 433.480 495.600 434.880 ;
        RECT 15.705 431.480 499.955 433.480 ;
        RECT 15.705 430.080 495.600 431.480 ;
        RECT 15.705 428.760 499.955 430.080 ;
        RECT 15.705 427.360 495.600 428.760 ;
        RECT 15.705 426.040 499.955 427.360 ;
        RECT 15.705 424.640 495.600 426.040 ;
        RECT 15.705 422.640 499.955 424.640 ;
        RECT 15.705 421.240 495.600 422.640 ;
        RECT 15.705 419.920 499.955 421.240 ;
        RECT 15.705 418.520 495.600 419.920 ;
        RECT 15.705 417.200 499.955 418.520 ;
        RECT 15.705 415.800 495.600 417.200 ;
        RECT 15.705 414.480 499.955 415.800 ;
        RECT 15.705 413.080 495.600 414.480 ;
        RECT 15.705 411.080 499.955 413.080 ;
        RECT 15.705 409.680 495.600 411.080 ;
        RECT 15.705 408.360 499.955 409.680 ;
        RECT 15.705 406.960 495.600 408.360 ;
        RECT 15.705 405.640 499.955 406.960 ;
        RECT 15.705 404.240 495.600 405.640 ;
        RECT 15.705 402.240 499.955 404.240 ;
        RECT 15.705 400.840 495.600 402.240 ;
        RECT 15.705 399.520 499.955 400.840 ;
        RECT 15.705 398.120 495.600 399.520 ;
        RECT 15.705 396.800 499.955 398.120 ;
        RECT 15.705 395.400 495.600 396.800 ;
        RECT 15.705 393.400 499.955 395.400 ;
        RECT 15.705 392.000 495.600 393.400 ;
        RECT 15.705 390.680 499.955 392.000 ;
        RECT 15.705 389.280 495.600 390.680 ;
        RECT 15.705 387.960 499.955 389.280 ;
        RECT 15.705 386.560 495.600 387.960 ;
        RECT 15.705 385.240 499.955 386.560 ;
        RECT 15.705 383.840 495.600 385.240 ;
        RECT 15.705 381.840 499.955 383.840 ;
        RECT 15.705 380.440 495.600 381.840 ;
        RECT 15.705 379.120 499.955 380.440 ;
        RECT 15.705 377.720 495.600 379.120 ;
        RECT 15.705 376.400 499.955 377.720 ;
        RECT 15.705 375.000 495.600 376.400 ;
        RECT 15.705 373.000 499.955 375.000 ;
        RECT 15.705 371.600 495.600 373.000 ;
        RECT 15.705 370.280 499.955 371.600 ;
        RECT 15.705 368.880 495.600 370.280 ;
        RECT 15.705 367.560 499.955 368.880 ;
        RECT 15.705 366.160 495.600 367.560 ;
        RECT 15.705 364.160 499.955 366.160 ;
        RECT 15.705 362.760 495.600 364.160 ;
        RECT 15.705 361.440 499.955 362.760 ;
        RECT 15.705 360.040 495.600 361.440 ;
        RECT 15.705 358.720 499.955 360.040 ;
        RECT 15.705 357.320 495.600 358.720 ;
        RECT 15.705 356.000 499.955 357.320 ;
        RECT 15.705 354.600 495.600 356.000 ;
        RECT 15.705 352.600 499.955 354.600 ;
        RECT 15.705 351.200 495.600 352.600 ;
        RECT 15.705 349.880 499.955 351.200 ;
        RECT 15.705 348.480 495.600 349.880 ;
        RECT 15.705 347.160 499.955 348.480 ;
        RECT 15.705 345.760 495.600 347.160 ;
        RECT 15.705 343.760 499.955 345.760 ;
        RECT 15.705 342.360 495.600 343.760 ;
        RECT 15.705 341.040 499.955 342.360 ;
        RECT 15.705 339.640 495.600 341.040 ;
        RECT 15.705 338.320 499.955 339.640 ;
        RECT 15.705 336.920 495.600 338.320 ;
        RECT 15.705 335.600 499.955 336.920 ;
        RECT 15.705 334.200 495.600 335.600 ;
        RECT 15.705 332.200 499.955 334.200 ;
        RECT 15.705 330.800 495.600 332.200 ;
        RECT 15.705 329.480 499.955 330.800 ;
        RECT 15.705 328.080 495.600 329.480 ;
        RECT 15.705 326.760 499.955 328.080 ;
        RECT 15.705 325.360 495.600 326.760 ;
        RECT 15.705 323.360 499.955 325.360 ;
        RECT 15.705 321.960 495.600 323.360 ;
        RECT 15.705 320.640 499.955 321.960 ;
        RECT 15.705 319.240 495.600 320.640 ;
        RECT 15.705 317.920 499.955 319.240 ;
        RECT 15.705 316.520 495.600 317.920 ;
        RECT 15.705 314.520 499.955 316.520 ;
        RECT 15.705 313.120 495.600 314.520 ;
        RECT 15.705 311.800 499.955 313.120 ;
        RECT 15.705 310.400 495.600 311.800 ;
        RECT 15.705 309.080 499.955 310.400 ;
        RECT 15.705 307.680 495.600 309.080 ;
        RECT 15.705 306.360 499.955 307.680 ;
        RECT 15.705 304.960 495.600 306.360 ;
        RECT 15.705 302.960 499.955 304.960 ;
        RECT 15.705 301.560 495.600 302.960 ;
        RECT 15.705 300.240 499.955 301.560 ;
        RECT 15.705 298.840 495.600 300.240 ;
        RECT 15.705 297.520 499.955 298.840 ;
        RECT 15.705 296.120 495.600 297.520 ;
        RECT 15.705 294.120 499.955 296.120 ;
        RECT 15.705 292.720 495.600 294.120 ;
        RECT 15.705 291.400 499.955 292.720 ;
        RECT 15.705 290.000 495.600 291.400 ;
        RECT 15.705 288.680 499.955 290.000 ;
        RECT 15.705 287.280 495.600 288.680 ;
        RECT 15.705 285.280 499.955 287.280 ;
        RECT 15.705 283.880 495.600 285.280 ;
        RECT 15.705 282.560 499.955 283.880 ;
        RECT 15.705 281.160 495.600 282.560 ;
        RECT 15.705 279.840 499.955 281.160 ;
        RECT 15.705 278.440 495.600 279.840 ;
        RECT 15.705 277.120 499.955 278.440 ;
        RECT 15.705 275.720 495.600 277.120 ;
        RECT 15.705 273.720 499.955 275.720 ;
        RECT 15.705 272.320 495.600 273.720 ;
        RECT 15.705 271.000 499.955 272.320 ;
        RECT 15.705 269.600 495.600 271.000 ;
        RECT 15.705 268.280 499.955 269.600 ;
        RECT 15.705 266.880 495.600 268.280 ;
        RECT 15.705 264.880 499.955 266.880 ;
        RECT 15.705 263.480 495.600 264.880 ;
        RECT 15.705 262.160 499.955 263.480 ;
        RECT 15.705 260.760 495.600 262.160 ;
        RECT 15.705 259.440 499.955 260.760 ;
        RECT 15.705 258.040 495.600 259.440 ;
        RECT 15.705 256.040 499.955 258.040 ;
        RECT 15.705 254.640 495.600 256.040 ;
        RECT 15.705 253.320 499.955 254.640 ;
        RECT 15.705 251.920 495.600 253.320 ;
        RECT 15.705 250.600 499.955 251.920 ;
        RECT 15.705 249.200 495.600 250.600 ;
        RECT 15.705 247.880 499.955 249.200 ;
        RECT 15.705 246.480 495.600 247.880 ;
        RECT 15.705 244.480 499.955 246.480 ;
        RECT 15.705 243.080 495.600 244.480 ;
        RECT 15.705 241.760 499.955 243.080 ;
        RECT 15.705 240.360 495.600 241.760 ;
        RECT 15.705 239.040 499.955 240.360 ;
        RECT 15.705 237.640 495.600 239.040 ;
        RECT 15.705 235.640 499.955 237.640 ;
        RECT 15.705 234.240 495.600 235.640 ;
        RECT 15.705 232.920 499.955 234.240 ;
        RECT 15.705 231.520 495.600 232.920 ;
        RECT 15.705 230.200 499.955 231.520 ;
        RECT 15.705 228.800 495.600 230.200 ;
        RECT 15.705 226.800 499.955 228.800 ;
        RECT 15.705 225.400 495.600 226.800 ;
        RECT 15.705 224.080 499.955 225.400 ;
        RECT 15.705 222.680 495.600 224.080 ;
        RECT 15.705 221.360 499.955 222.680 ;
        RECT 15.705 219.960 495.600 221.360 ;
        RECT 15.705 218.640 499.955 219.960 ;
        RECT 15.705 217.240 495.600 218.640 ;
        RECT 15.705 215.240 499.955 217.240 ;
        RECT 15.705 213.840 495.600 215.240 ;
        RECT 15.705 212.520 499.955 213.840 ;
        RECT 15.705 211.120 495.600 212.520 ;
        RECT 15.705 209.800 499.955 211.120 ;
        RECT 15.705 208.400 495.600 209.800 ;
        RECT 15.705 206.400 499.955 208.400 ;
        RECT 15.705 205.000 495.600 206.400 ;
        RECT 15.705 203.680 499.955 205.000 ;
        RECT 15.705 202.280 495.600 203.680 ;
        RECT 15.705 200.960 499.955 202.280 ;
        RECT 15.705 199.560 495.600 200.960 ;
        RECT 15.705 197.560 499.955 199.560 ;
        RECT 15.705 196.160 495.600 197.560 ;
        RECT 15.705 194.840 499.955 196.160 ;
        RECT 15.705 193.440 495.600 194.840 ;
        RECT 15.705 192.120 499.955 193.440 ;
        RECT 15.705 190.720 495.600 192.120 ;
        RECT 15.705 189.400 499.955 190.720 ;
        RECT 15.705 188.000 495.600 189.400 ;
        RECT 15.705 186.000 499.955 188.000 ;
        RECT 15.705 184.600 495.600 186.000 ;
        RECT 15.705 183.280 499.955 184.600 ;
        RECT 15.705 181.880 495.600 183.280 ;
        RECT 15.705 180.560 499.955 181.880 ;
        RECT 15.705 179.160 495.600 180.560 ;
        RECT 15.705 177.160 499.955 179.160 ;
        RECT 15.705 175.760 495.600 177.160 ;
        RECT 15.705 174.440 499.955 175.760 ;
        RECT 15.705 173.040 495.600 174.440 ;
        RECT 15.705 171.720 499.955 173.040 ;
        RECT 15.705 170.320 495.600 171.720 ;
        RECT 15.705 169.000 499.955 170.320 ;
        RECT 15.705 167.600 495.600 169.000 ;
        RECT 15.705 165.600 499.955 167.600 ;
        RECT 15.705 164.200 495.600 165.600 ;
        RECT 15.705 162.880 499.955 164.200 ;
        RECT 15.705 161.480 495.600 162.880 ;
        RECT 15.705 160.160 499.955 161.480 ;
        RECT 15.705 158.760 495.600 160.160 ;
        RECT 15.705 156.760 499.955 158.760 ;
        RECT 15.705 155.360 495.600 156.760 ;
        RECT 15.705 154.040 499.955 155.360 ;
        RECT 15.705 152.640 495.600 154.040 ;
        RECT 15.705 151.320 499.955 152.640 ;
        RECT 15.705 149.920 495.600 151.320 ;
        RECT 15.705 147.920 499.955 149.920 ;
        RECT 15.705 146.520 495.600 147.920 ;
        RECT 15.705 145.200 499.955 146.520 ;
        RECT 15.705 143.800 495.600 145.200 ;
        RECT 15.705 142.480 499.955 143.800 ;
        RECT 15.705 141.080 495.600 142.480 ;
        RECT 15.705 139.760 499.955 141.080 ;
        RECT 15.705 138.360 495.600 139.760 ;
        RECT 15.705 136.360 499.955 138.360 ;
        RECT 15.705 134.960 495.600 136.360 ;
        RECT 15.705 133.640 499.955 134.960 ;
        RECT 15.705 132.240 495.600 133.640 ;
        RECT 15.705 130.920 499.955 132.240 ;
        RECT 15.705 129.520 495.600 130.920 ;
        RECT 15.705 127.520 499.955 129.520 ;
        RECT 15.705 126.120 495.600 127.520 ;
        RECT 15.705 124.800 499.955 126.120 ;
        RECT 15.705 123.400 495.600 124.800 ;
        RECT 15.705 122.080 499.955 123.400 ;
        RECT 15.705 120.680 495.600 122.080 ;
        RECT 15.705 118.680 499.955 120.680 ;
        RECT 15.705 117.280 495.600 118.680 ;
        RECT 15.705 115.960 499.955 117.280 ;
        RECT 15.705 114.560 495.600 115.960 ;
        RECT 15.705 113.240 499.955 114.560 ;
        RECT 15.705 111.840 495.600 113.240 ;
        RECT 15.705 110.520 499.955 111.840 ;
        RECT 15.705 109.120 495.600 110.520 ;
        RECT 15.705 107.120 499.955 109.120 ;
        RECT 15.705 105.720 495.600 107.120 ;
        RECT 15.705 104.400 499.955 105.720 ;
        RECT 15.705 103.000 495.600 104.400 ;
        RECT 15.705 101.680 499.955 103.000 ;
        RECT 15.705 100.280 495.600 101.680 ;
        RECT 15.705 98.280 499.955 100.280 ;
        RECT 15.705 96.880 495.600 98.280 ;
        RECT 15.705 95.560 499.955 96.880 ;
        RECT 15.705 94.160 495.600 95.560 ;
        RECT 15.705 92.840 499.955 94.160 ;
        RECT 15.705 91.440 495.600 92.840 ;
        RECT 15.705 89.440 499.955 91.440 ;
        RECT 15.705 88.040 495.600 89.440 ;
        RECT 15.705 86.720 499.955 88.040 ;
        RECT 15.705 85.320 495.600 86.720 ;
        RECT 15.705 84.000 499.955 85.320 ;
        RECT 15.705 82.600 495.600 84.000 ;
        RECT 15.705 81.280 499.955 82.600 ;
        RECT 15.705 79.880 495.600 81.280 ;
        RECT 15.705 77.880 499.955 79.880 ;
        RECT 15.705 76.480 495.600 77.880 ;
        RECT 15.705 75.160 499.955 76.480 ;
        RECT 15.705 73.760 495.600 75.160 ;
        RECT 15.705 72.440 499.955 73.760 ;
        RECT 15.705 71.040 495.600 72.440 ;
        RECT 15.705 69.040 499.955 71.040 ;
        RECT 15.705 67.640 495.600 69.040 ;
        RECT 15.705 66.320 499.955 67.640 ;
        RECT 15.705 64.920 495.600 66.320 ;
        RECT 15.705 63.600 499.955 64.920 ;
        RECT 15.705 62.200 495.600 63.600 ;
        RECT 15.705 60.200 499.955 62.200 ;
        RECT 15.705 58.800 495.600 60.200 ;
        RECT 15.705 57.480 499.955 58.800 ;
        RECT 15.705 56.080 495.600 57.480 ;
        RECT 15.705 54.760 499.955 56.080 ;
        RECT 15.705 53.360 495.600 54.760 ;
        RECT 15.705 52.040 499.955 53.360 ;
        RECT 15.705 50.640 495.600 52.040 ;
        RECT 15.705 48.640 499.955 50.640 ;
        RECT 15.705 47.240 495.600 48.640 ;
        RECT 15.705 45.920 499.955 47.240 ;
        RECT 15.705 44.520 495.600 45.920 ;
        RECT 15.705 43.200 499.955 44.520 ;
        RECT 15.705 41.800 495.600 43.200 ;
        RECT 15.705 39.800 499.955 41.800 ;
        RECT 15.705 38.400 495.600 39.800 ;
        RECT 15.705 37.080 499.955 38.400 ;
        RECT 15.705 35.680 495.600 37.080 ;
        RECT 15.705 34.360 499.955 35.680 ;
        RECT 15.705 32.960 495.600 34.360 ;
        RECT 15.705 30.960 499.955 32.960 ;
        RECT 15.705 29.560 495.600 30.960 ;
        RECT 15.705 28.240 499.955 29.560 ;
        RECT 15.705 26.840 495.600 28.240 ;
        RECT 15.705 25.520 499.955 26.840 ;
        RECT 15.705 24.120 495.600 25.520 ;
        RECT 15.705 22.800 499.955 24.120 ;
        RECT 15.705 21.400 495.600 22.800 ;
        RECT 15.705 19.400 499.955 21.400 ;
        RECT 15.705 18.000 495.600 19.400 ;
        RECT 15.705 16.680 499.955 18.000 ;
        RECT 15.705 15.280 495.600 16.680 ;
        RECT 15.705 13.960 499.955 15.280 ;
        RECT 15.705 12.560 495.600 13.960 ;
        RECT 15.705 10.560 499.955 12.560 ;
        RECT 15.705 9.160 495.600 10.560 ;
        RECT 15.705 7.840 499.955 9.160 ;
        RECT 15.705 6.440 495.600 7.840 ;
        RECT 15.705 5.120 499.955 6.440 ;
        RECT 15.705 3.720 495.600 5.120 ;
        RECT 15.705 2.400 499.955 3.720 ;
        RECT 15.705 1.535 495.600 2.400 ;
      LAYER met4 ;
        RECT 41.695 13.095 97.440 486.025 ;
        RECT 99.840 13.095 174.240 486.025 ;
        RECT 176.640 13.095 251.040 486.025 ;
        RECT 253.440 13.095 327.840 486.025 ;
        RECT 330.240 13.095 404.640 486.025 ;
        RECT 407.040 13.095 481.440 486.025 ;
        RECT 483.840 13.095 490.985 486.025 ;
  END
END Core
END LIBRARY

