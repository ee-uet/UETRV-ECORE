magic
tech sky130A
magscale 1 2
timestamp 1647754903
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 14 1708 99898 97640
<< metal2 >>
rect 1306 99200 1362 100000
rect 3882 99200 3938 100000
rect 5814 99200 5870 100000
rect 8390 99200 8446 100000
rect 10322 99200 10378 100000
rect 12898 99200 12954 100000
rect 14830 99200 14886 100000
rect 17406 99200 17462 100000
rect 19338 99200 19394 100000
rect 21914 99200 21970 100000
rect 23846 99200 23902 100000
rect 26422 99200 26478 100000
rect 28354 99200 28410 100000
rect 30930 99200 30986 100000
rect 32862 99200 32918 100000
rect 34794 99200 34850 100000
rect 37370 99200 37426 100000
rect 39302 99200 39358 100000
rect 41878 99200 41934 100000
rect 43810 99200 43866 100000
rect 46386 99200 46442 100000
rect 48318 99200 48374 100000
rect 50894 99200 50950 100000
rect 52826 99200 52882 100000
rect 55402 99200 55458 100000
rect 57334 99200 57390 100000
rect 59910 99200 59966 100000
rect 61842 99200 61898 100000
rect 64418 99200 64474 100000
rect 66350 99200 66406 100000
rect 68926 99200 68982 100000
rect 70858 99200 70914 100000
rect 73434 99200 73490 100000
rect 75366 99200 75422 100000
rect 77942 99200 77998 100000
rect 79874 99200 79930 100000
rect 82450 99200 82506 100000
rect 84382 99200 84438 100000
rect 86958 99200 87014 100000
rect 88890 99200 88946 100000
rect 91466 99200 91522 100000
rect 93398 99200 93454 100000
rect 95974 99200 96030 100000
rect 97906 99200 97962 100000
rect 99838 99200 99894 100000
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 15474 0 15530 800
rect 17406 0 17462 800
rect 19982 0 20038 800
rect 21914 0 21970 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 28998 0 29054 800
rect 30930 0 30986 800
rect 33506 0 33562 800
rect 35438 0 35494 800
rect 38014 0 38070 800
rect 39946 0 40002 800
rect 42522 0 42578 800
rect 44454 0 44510 800
rect 47030 0 47086 800
rect 48962 0 49018 800
rect 51538 0 51594 800
rect 53470 0 53526 800
rect 56046 0 56102 800
rect 57978 0 58034 800
rect 60554 0 60610 800
rect 62486 0 62542 800
rect 65062 0 65118 800
rect 66994 0 67050 800
rect 68926 0 68982 800
rect 71502 0 71558 800
rect 73434 0 73490 800
rect 76010 0 76066 800
rect 77942 0 77998 800
rect 80518 0 80574 800
rect 82450 0 82506 800
rect 85026 0 85082 800
rect 86958 0 87014 800
rect 89534 0 89590 800
rect 91466 0 91522 800
rect 94042 0 94098 800
rect 95974 0 96030 800
rect 98550 0 98606 800
<< obsm2 >>
rect 20 99144 1250 99385
rect 1418 99144 3826 99385
rect 3994 99144 5758 99385
rect 5926 99144 8334 99385
rect 8502 99144 10266 99385
rect 10434 99144 12842 99385
rect 13010 99144 14774 99385
rect 14942 99144 17350 99385
rect 17518 99144 19282 99385
rect 19450 99144 21858 99385
rect 22026 99144 23790 99385
rect 23958 99144 26366 99385
rect 26534 99144 28298 99385
rect 28466 99144 30874 99385
rect 31042 99144 32806 99385
rect 32974 99144 34738 99385
rect 34906 99144 37314 99385
rect 37482 99144 39246 99385
rect 39414 99144 41822 99385
rect 41990 99144 43754 99385
rect 43922 99144 46330 99385
rect 46498 99144 48262 99385
rect 48430 99144 50838 99385
rect 51006 99144 52770 99385
rect 52938 99144 55346 99385
rect 55514 99144 57278 99385
rect 57446 99144 59854 99385
rect 60022 99144 61786 99385
rect 61954 99144 64362 99385
rect 64530 99144 66294 99385
rect 66462 99144 68870 99385
rect 69038 99144 70802 99385
rect 70970 99144 73378 99385
rect 73546 99144 75310 99385
rect 75478 99144 77886 99385
rect 78054 99144 79818 99385
rect 79986 99144 82394 99385
rect 82562 99144 84326 99385
rect 84494 99144 86902 99385
rect 87070 99144 88834 99385
rect 89002 99144 91410 99385
rect 91578 99144 93342 99385
rect 93510 99144 95918 99385
rect 96086 99144 97850 99385
rect 98018 99144 99782 99385
rect 20 856 99892 99144
rect 130 31 1894 856
rect 2062 31 3826 856
rect 3994 31 6402 856
rect 6570 31 8334 856
rect 8502 31 10910 856
rect 11078 31 12842 856
rect 13010 31 15418 856
rect 15586 31 17350 856
rect 17518 31 19926 856
rect 20094 31 21858 856
rect 22026 31 24434 856
rect 24602 31 26366 856
rect 26534 31 28942 856
rect 29110 31 30874 856
rect 31042 31 33450 856
rect 33618 31 35382 856
rect 35550 31 37958 856
rect 38126 31 39890 856
rect 40058 31 42466 856
rect 42634 31 44398 856
rect 44566 31 46974 856
rect 47142 31 48906 856
rect 49074 31 51482 856
rect 51650 31 53414 856
rect 53582 31 55990 856
rect 56158 31 57922 856
rect 58090 31 60498 856
rect 60666 31 62430 856
rect 62598 31 65006 856
rect 65174 31 66938 856
rect 67106 31 68870 856
rect 69038 31 71446 856
rect 71614 31 73378 856
rect 73546 31 75954 856
rect 76122 31 77886 856
rect 78054 31 80462 856
rect 80630 31 82394 856
rect 82562 31 84970 856
rect 85138 31 86902 856
rect 87070 31 89478 856
rect 89646 31 91410 856
rect 91578 31 93986 856
rect 94154 31 95918 856
rect 96086 31 98494 856
rect 98662 31 99892 856
<< metal3 >>
rect 0 99288 800 99408
rect 99200 97248 100000 97368
rect 0 96568 800 96688
rect 99200 95208 100000 95328
rect 0 94528 800 94648
rect 99200 92488 100000 92608
rect 0 91808 800 91928
rect 99200 90448 100000 90568
rect 0 89768 800 89888
rect 99200 87728 100000 87848
rect 0 87048 800 87168
rect 99200 85688 100000 85808
rect 0 85008 800 85128
rect 99200 82968 100000 83088
rect 0 82288 800 82408
rect 99200 80928 100000 81048
rect 0 80248 800 80368
rect 99200 78208 100000 78328
rect 0 77528 800 77648
rect 99200 76168 100000 76288
rect 0 75488 800 75608
rect 99200 73448 100000 73568
rect 0 72768 800 72888
rect 99200 71408 100000 71528
rect 0 70728 800 70848
rect 99200 68688 100000 68808
rect 0 68008 800 68128
rect 99200 66648 100000 66768
rect 0 65968 800 66088
rect 0 63928 800 64048
rect 99200 63928 100000 64048
rect 99200 61888 100000 62008
rect 0 61208 800 61328
rect 0 59168 800 59288
rect 99200 59168 100000 59288
rect 99200 57128 100000 57248
rect 0 56448 800 56568
rect 0 54408 800 54528
rect 99200 54408 100000 54528
rect 99200 52368 100000 52488
rect 0 51688 800 51808
rect 0 49648 800 49768
rect 99200 49648 100000 49768
rect 99200 47608 100000 47728
rect 0 46928 800 47048
rect 0 44888 800 45008
rect 99200 44888 100000 45008
rect 99200 42848 100000 42968
rect 0 42168 800 42288
rect 0 40128 800 40248
rect 99200 40128 100000 40248
rect 99200 38088 100000 38208
rect 0 37408 800 37528
rect 0 35368 800 35488
rect 99200 35368 100000 35488
rect 99200 33328 100000 33448
rect 0 32648 800 32768
rect 99200 31288 100000 31408
rect 0 30608 800 30728
rect 99200 28568 100000 28688
rect 0 27888 800 28008
rect 99200 26528 100000 26648
rect 0 25848 800 25968
rect 99200 23808 100000 23928
rect 0 23128 800 23248
rect 99200 21768 100000 21888
rect 0 21088 800 21208
rect 99200 19048 100000 19168
rect 0 18368 800 18488
rect 99200 17008 100000 17128
rect 0 16328 800 16448
rect 99200 14288 100000 14408
rect 0 13608 800 13728
rect 99200 12248 100000 12368
rect 0 11568 800 11688
rect 99200 9528 100000 9648
rect 0 8848 800 8968
rect 99200 7488 100000 7608
rect 0 6808 800 6928
rect 99200 4768 100000 4888
rect 0 4088 800 4208
rect 99200 2728 100000 2848
rect 0 2048 800 2168
rect 99200 8 100000 128
<< obsm3 >>
rect 880 99208 99200 99381
rect 749 97448 99200 99208
rect 749 97168 99120 97448
rect 749 96768 99200 97168
rect 880 96488 99200 96768
rect 749 95408 99200 96488
rect 749 95128 99120 95408
rect 749 94728 99200 95128
rect 880 94448 99200 94728
rect 749 92688 99200 94448
rect 749 92408 99120 92688
rect 749 92008 99200 92408
rect 880 91728 99200 92008
rect 749 90648 99200 91728
rect 749 90368 99120 90648
rect 749 89968 99200 90368
rect 880 89688 99200 89968
rect 749 87928 99200 89688
rect 749 87648 99120 87928
rect 749 87248 99200 87648
rect 880 86968 99200 87248
rect 749 85888 99200 86968
rect 749 85608 99120 85888
rect 749 85208 99200 85608
rect 880 84928 99200 85208
rect 749 83168 99200 84928
rect 749 82888 99120 83168
rect 749 82488 99200 82888
rect 880 82208 99200 82488
rect 749 81128 99200 82208
rect 749 80848 99120 81128
rect 749 80448 99200 80848
rect 880 80168 99200 80448
rect 749 78408 99200 80168
rect 749 78128 99120 78408
rect 749 77728 99200 78128
rect 880 77448 99200 77728
rect 749 76368 99200 77448
rect 749 76088 99120 76368
rect 749 75688 99200 76088
rect 880 75408 99200 75688
rect 749 73648 99200 75408
rect 749 73368 99120 73648
rect 749 72968 99200 73368
rect 880 72688 99200 72968
rect 749 71608 99200 72688
rect 749 71328 99120 71608
rect 749 70928 99200 71328
rect 880 70648 99200 70928
rect 749 68888 99200 70648
rect 749 68608 99120 68888
rect 749 68208 99200 68608
rect 880 67928 99200 68208
rect 749 66848 99200 67928
rect 749 66568 99120 66848
rect 749 66168 99200 66568
rect 880 65888 99200 66168
rect 749 64128 99200 65888
rect 880 63848 99120 64128
rect 749 62088 99200 63848
rect 749 61808 99120 62088
rect 749 61408 99200 61808
rect 880 61128 99200 61408
rect 749 59368 99200 61128
rect 880 59088 99120 59368
rect 749 57328 99200 59088
rect 749 57048 99120 57328
rect 749 56648 99200 57048
rect 880 56368 99200 56648
rect 749 54608 99200 56368
rect 880 54328 99120 54608
rect 749 52568 99200 54328
rect 749 52288 99120 52568
rect 749 51888 99200 52288
rect 880 51608 99200 51888
rect 749 49848 99200 51608
rect 880 49568 99120 49848
rect 749 47808 99200 49568
rect 749 47528 99120 47808
rect 749 47128 99200 47528
rect 880 46848 99200 47128
rect 749 45088 99200 46848
rect 880 44808 99120 45088
rect 749 43048 99200 44808
rect 749 42768 99120 43048
rect 749 42368 99200 42768
rect 880 42088 99200 42368
rect 749 40328 99200 42088
rect 880 40048 99120 40328
rect 749 38288 99200 40048
rect 749 38008 99120 38288
rect 749 37608 99200 38008
rect 880 37328 99200 37608
rect 749 35568 99200 37328
rect 880 35288 99120 35568
rect 749 33528 99200 35288
rect 749 33248 99120 33528
rect 749 32848 99200 33248
rect 880 32568 99200 32848
rect 749 31488 99200 32568
rect 749 31208 99120 31488
rect 749 30808 99200 31208
rect 880 30528 99200 30808
rect 749 28768 99200 30528
rect 749 28488 99120 28768
rect 749 28088 99200 28488
rect 880 27808 99200 28088
rect 749 26728 99200 27808
rect 749 26448 99120 26728
rect 749 26048 99200 26448
rect 880 25768 99200 26048
rect 749 24008 99200 25768
rect 749 23728 99120 24008
rect 749 23328 99200 23728
rect 880 23048 99200 23328
rect 749 21968 99200 23048
rect 749 21688 99120 21968
rect 749 21288 99200 21688
rect 880 21008 99200 21288
rect 749 19248 99200 21008
rect 749 18968 99120 19248
rect 749 18568 99200 18968
rect 880 18288 99200 18568
rect 749 17208 99200 18288
rect 749 16928 99120 17208
rect 749 16528 99200 16928
rect 880 16248 99200 16528
rect 749 14488 99200 16248
rect 749 14208 99120 14488
rect 749 13808 99200 14208
rect 880 13528 99200 13808
rect 749 12448 99200 13528
rect 749 12168 99120 12448
rect 749 11768 99200 12168
rect 880 11488 99200 11768
rect 749 9728 99200 11488
rect 749 9448 99120 9728
rect 749 9048 99200 9448
rect 880 8768 99200 9048
rect 749 7688 99200 8768
rect 749 7408 99120 7688
rect 749 7008 99200 7408
rect 880 6728 99200 7008
rect 749 4968 99200 6728
rect 749 4688 99120 4968
rect 749 4288 99200 4688
rect 880 4008 99200 4288
rect 749 2928 99200 4008
rect 749 2648 99120 2928
rect 749 2248 99200 2648
rect 880 1968 99200 2248
rect 749 208 99200 1968
rect 749 35 99120 208
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 1163 97504 97645 97613
rect 1163 2048 4128 97504
rect 4608 2048 19488 97504
rect 19968 2048 34848 97504
rect 35328 2048 50208 97504
rect 50688 2048 65568 97504
rect 66048 2048 80928 97504
rect 81408 2048 96288 97504
rect 96768 2048 97645 97504
rect 1163 1803 97645 2048
<< labels >>
rlabel metal2 s 19338 99200 19394 100000 6 clock
port 1 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 io_dbus_addr[0]
port 2 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_dbus_addr[10]
port 3 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 io_dbus_addr[11]
port 4 nsew signal output
rlabel metal3 s 99200 42848 100000 42968 6 io_dbus_addr[12]
port 5 nsew signal output
rlabel metal2 s 64418 99200 64474 100000 6 io_dbus_addr[13]
port 6 nsew signal output
rlabel metal2 s 5814 99200 5870 100000 6 io_dbus_addr[14]
port 7 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 io_dbus_addr[15]
port 8 nsew signal output
rlabel metal3 s 99200 7488 100000 7608 6 io_dbus_addr[16]
port 9 nsew signal output
rlabel metal2 s 95974 99200 96030 100000 6 io_dbus_addr[17]
port 10 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 io_dbus_addr[18]
port 11 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 io_dbus_addr[19]
port 12 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 io_dbus_addr[1]
port 13 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 io_dbus_addr[20]
port 14 nsew signal output
rlabel metal3 s 99200 17008 100000 17128 6 io_dbus_addr[21]
port 15 nsew signal output
rlabel metal2 s 46386 99200 46442 100000 6 io_dbus_addr[22]
port 16 nsew signal output
rlabel metal3 s 99200 76168 100000 76288 6 io_dbus_addr[23]
port 17 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 io_dbus_addr[24]
port 18 nsew signal output
rlabel metal2 s 43810 99200 43866 100000 6 io_dbus_addr[25]
port 19 nsew signal output
rlabel metal2 s 57334 99200 57390 100000 6 io_dbus_addr[26]
port 20 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 io_dbus_addr[27]
port 21 nsew signal output
rlabel metal3 s 99200 78208 100000 78328 6 io_dbus_addr[28]
port 22 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 io_dbus_addr[29]
port 23 nsew signal output
rlabel metal2 s 23846 99200 23902 100000 6 io_dbus_addr[2]
port 24 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 io_dbus_addr[30]
port 25 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 io_dbus_addr[31]
port 26 nsew signal output
rlabel metal3 s 99200 9528 100000 9648 6 io_dbus_addr[3]
port 27 nsew signal output
rlabel metal3 s 99200 95208 100000 95328 6 io_dbus_addr[4]
port 28 nsew signal output
rlabel metal2 s 12898 99200 12954 100000 6 io_dbus_addr[5]
port 29 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 io_dbus_addr[6]
port 30 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 io_dbus_addr[7]
port 31 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 io_dbus_addr[8]
port 32 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 io_dbus_addr[9]
port 33 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 io_dbus_ld_type[0]
port 34 nsew signal output
rlabel metal3 s 99200 14288 100000 14408 6 io_dbus_ld_type[1]
port 35 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 io_dbus_ld_type[2]
port 36 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 io_dbus_rd_en
port 37 nsew signal output
rlabel metal2 s 8390 99200 8446 100000 6 io_dbus_rdata[0]
port 38 nsew signal input
rlabel metal2 s 3882 99200 3938 100000 6 io_dbus_rdata[10]
port 39 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 io_dbus_rdata[11]
port 40 nsew signal input
rlabel metal2 s 88890 99200 88946 100000 6 io_dbus_rdata[12]
port 41 nsew signal input
rlabel metal3 s 99200 63928 100000 64048 6 io_dbus_rdata[13]
port 42 nsew signal input
rlabel metal2 s 61842 99200 61898 100000 6 io_dbus_rdata[14]
port 43 nsew signal input
rlabel metal2 s 79874 99200 79930 100000 6 io_dbus_rdata[15]
port 44 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 io_dbus_rdata[16]
port 45 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 io_dbus_rdata[17]
port 46 nsew signal input
rlabel metal2 s 91466 99200 91522 100000 6 io_dbus_rdata[18]
port 47 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 io_dbus_rdata[19]
port 48 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 io_dbus_rdata[1]
port 49 nsew signal input
rlabel metal3 s 99200 80928 100000 81048 6 io_dbus_rdata[20]
port 50 nsew signal input
rlabel metal3 s 99200 54408 100000 54528 6 io_dbus_rdata[21]
port 51 nsew signal input
rlabel metal2 s 93398 99200 93454 100000 6 io_dbus_rdata[22]
port 52 nsew signal input
rlabel metal2 s 41878 99200 41934 100000 6 io_dbus_rdata[23]
port 53 nsew signal input
rlabel metal3 s 99200 49648 100000 49768 6 io_dbus_rdata[24]
port 54 nsew signal input
rlabel metal2 s 26422 99200 26478 100000 6 io_dbus_rdata[25]
port 55 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 io_dbus_rdata[26]
port 56 nsew signal input
rlabel metal2 s 34794 99200 34850 100000 6 io_dbus_rdata[27]
port 57 nsew signal input
rlabel metal3 s 99200 68688 100000 68808 6 io_dbus_rdata[28]
port 58 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 io_dbus_rdata[29]
port 59 nsew signal input
rlabel metal2 s 86958 99200 87014 100000 6 io_dbus_rdata[2]
port 60 nsew signal input
rlabel metal2 s 99838 99200 99894 100000 6 io_dbus_rdata[30]
port 61 nsew signal input
rlabel metal2 s 37370 99200 37426 100000 6 io_dbus_rdata[31]
port 62 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 io_dbus_rdata[3]
port 63 nsew signal input
rlabel metal3 s 99200 31288 100000 31408 6 io_dbus_rdata[4]
port 64 nsew signal input
rlabel metal3 s 99200 4768 100000 4888 6 io_dbus_rdata[5]
port 65 nsew signal input
rlabel metal2 s 59910 99200 59966 100000 6 io_dbus_rdata[6]
port 66 nsew signal input
rlabel metal3 s 99200 87728 100000 87848 6 io_dbus_rdata[7]
port 67 nsew signal input
rlabel metal3 s 99200 35368 100000 35488 6 io_dbus_rdata[8]
port 68 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 io_dbus_rdata[9]
port 69 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 io_dbus_st_type[0]
port 70 nsew signal output
rlabel metal2 s 68926 99200 68982 100000 6 io_dbus_st_type[1]
port 71 nsew signal output
rlabel metal3 s 99200 90448 100000 90568 6 io_dbus_valid
port 72 nsew signal input
rlabel metal2 s 28354 99200 28410 100000 6 io_dbus_wdata[0]
port 73 nsew signal output
rlabel metal3 s 99200 61888 100000 62008 6 io_dbus_wdata[10]
port 74 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 io_dbus_wdata[11]
port 75 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 io_dbus_wdata[12]
port 76 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 io_dbus_wdata[13]
port 77 nsew signal output
rlabel metal2 s 82450 99200 82506 100000 6 io_dbus_wdata[14]
port 78 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 io_dbus_wdata[15]
port 79 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 io_dbus_wdata[16]
port 80 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 io_dbus_wdata[17]
port 81 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 io_dbus_wdata[18]
port 82 nsew signal output
rlabel metal3 s 99200 40128 100000 40248 6 io_dbus_wdata[19]
port 83 nsew signal output
rlabel metal3 s 99200 23808 100000 23928 6 io_dbus_wdata[1]
port 84 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 io_dbus_wdata[20]
port 85 nsew signal output
rlabel metal2 s 39302 99200 39358 100000 6 io_dbus_wdata[21]
port 86 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 io_dbus_wdata[22]
port 87 nsew signal output
rlabel metal3 s 99200 82968 100000 83088 6 io_dbus_wdata[23]
port 88 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 io_dbus_wdata[24]
port 89 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 io_dbus_wdata[25]
port 90 nsew signal output
rlabel metal3 s 99200 71408 100000 71528 6 io_dbus_wdata[26]
port 91 nsew signal output
rlabel metal3 s 99200 8 100000 128 6 io_dbus_wdata[27]
port 92 nsew signal output
rlabel metal3 s 99200 26528 100000 26648 6 io_dbus_wdata[28]
port 93 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 io_dbus_wdata[29]
port 94 nsew signal output
rlabel metal3 s 99200 44888 100000 45008 6 io_dbus_wdata[2]
port 95 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 io_dbus_wdata[30]
port 96 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 io_dbus_wdata[31]
port 97 nsew signal output
rlabel metal3 s 99200 52368 100000 52488 6 io_dbus_wdata[3]
port 98 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 io_dbus_wdata[4]
port 99 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 io_dbus_wdata[5]
port 100 nsew signal output
rlabel metal2 s 52826 99200 52882 100000 6 io_dbus_wdata[6]
port 101 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 io_dbus_wdata[7]
port 102 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 io_dbus_wdata[8]
port 103 nsew signal output
rlabel metal3 s 99200 92488 100000 92608 6 io_dbus_wdata[9]
port 104 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 io_dbus_wr_en
port 105 nsew signal output
rlabel metal2 s 55402 99200 55458 100000 6 io_ibus_addr[0]
port 106 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 io_ibus_addr[10]
port 107 nsew signal output
rlabel metal2 s 66350 99200 66406 100000 6 io_ibus_addr[11]
port 108 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 io_ibus_addr[12]
port 109 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 io_ibus_addr[13]
port 110 nsew signal output
rlabel metal3 s 99200 12248 100000 12368 6 io_ibus_addr[14]
port 111 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 io_ibus_addr[15]
port 112 nsew signal output
rlabel metal2 s 21914 99200 21970 100000 6 io_ibus_addr[16]
port 113 nsew signal output
rlabel metal2 s 30930 99200 30986 100000 6 io_ibus_addr[17]
port 114 nsew signal output
rlabel metal2 s 75366 99200 75422 100000 6 io_ibus_addr[18]
port 115 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 io_ibus_addr[19]
port 116 nsew signal output
rlabel metal3 s 99200 21768 100000 21888 6 io_ibus_addr[1]
port 117 nsew signal output
rlabel metal3 s 99200 57128 100000 57248 6 io_ibus_addr[20]
port 118 nsew signal output
rlabel metal2 s 32862 99200 32918 100000 6 io_ibus_addr[21]
port 119 nsew signal output
rlabel metal3 s 99200 38088 100000 38208 6 io_ibus_addr[22]
port 120 nsew signal output
rlabel metal2 s 10322 99200 10378 100000 6 io_ibus_addr[23]
port 121 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 io_ibus_addr[24]
port 122 nsew signal output
rlabel metal3 s 99200 73448 100000 73568 6 io_ibus_addr[25]
port 123 nsew signal output
rlabel metal2 s 77942 99200 77998 100000 6 io_ibus_addr[26]
port 124 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 io_ibus_addr[27]
port 125 nsew signal output
rlabel metal3 s 99200 28568 100000 28688 6 io_ibus_addr[28]
port 126 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 io_ibus_addr[29]
port 127 nsew signal output
rlabel metal3 s 99200 2728 100000 2848 6 io_ibus_addr[2]
port 128 nsew signal output
rlabel metal2 s 14830 99200 14886 100000 6 io_ibus_addr[30]
port 129 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 io_ibus_addr[31]
port 130 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 io_ibus_addr[3]
port 131 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 io_ibus_addr[4]
port 132 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 io_ibus_addr[5]
port 133 nsew signal output
rlabel metal3 s 99200 85688 100000 85808 6 io_ibus_addr[6]
port 134 nsew signal output
rlabel metal3 s 99200 59168 100000 59288 6 io_ibus_addr[7]
port 135 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 io_ibus_addr[8]
port 136 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 io_ibus_addr[9]
port 137 nsew signal output
rlabel metal3 s 99200 33328 100000 33448 6 io_ibus_inst[0]
port 138 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 io_ibus_inst[10]
port 139 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 io_ibus_inst[11]
port 140 nsew signal input
rlabel metal3 s 99200 97248 100000 97368 6 io_ibus_inst[12]
port 141 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 io_ibus_inst[13]
port 142 nsew signal input
rlabel metal2 s 97906 99200 97962 100000 6 io_ibus_inst[14]
port 143 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 io_ibus_inst[15]
port 144 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 io_ibus_inst[16]
port 145 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 io_ibus_inst[17]
port 146 nsew signal input
rlabel metal2 s 18 0 74 800 6 io_ibus_inst[18]
port 147 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 io_ibus_inst[19]
port 148 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 io_ibus_inst[1]
port 149 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 io_ibus_inst[20]
port 150 nsew signal input
rlabel metal2 s 50894 99200 50950 100000 6 io_ibus_inst[21]
port 151 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 io_ibus_inst[22]
port 152 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 io_ibus_inst[23]
port 153 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_ibus_inst[24]
port 154 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 io_ibus_inst[25]
port 155 nsew signal input
rlabel metal2 s 48318 99200 48374 100000 6 io_ibus_inst[26]
port 156 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 io_ibus_inst[27]
port 157 nsew signal input
rlabel metal2 s 84382 99200 84438 100000 6 io_ibus_inst[28]
port 158 nsew signal input
rlabel metal3 s 99200 19048 100000 19168 6 io_ibus_inst[29]
port 159 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 io_ibus_inst[2]
port 160 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 io_ibus_inst[30]
port 161 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 io_ibus_inst[31]
port 162 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 io_ibus_inst[3]
port 163 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 io_ibus_inst[4]
port 164 nsew signal input
rlabel metal3 s 99200 66648 100000 66768 6 io_ibus_inst[5]
port 165 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 io_ibus_inst[6]
port 166 nsew signal input
rlabel metal2 s 73434 99200 73490 100000 6 io_ibus_inst[7]
port 167 nsew signal input
rlabel metal2 s 70858 99200 70914 100000 6 io_ibus_inst[8]
port 168 nsew signal input
rlabel metal2 s 1306 99200 1362 100000 6 io_ibus_inst[9]
port 169 nsew signal input
rlabel metal2 s 17406 99200 17462 100000 6 io_ibus_valid
port 170 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 io_irq_motor_irq
port 171 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 io_irq_spi_irq
port 172 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 io_irq_uart_irq
port 173 nsew signal input
rlabel metal3 s 99200 47608 100000 47728 6 reset
port 174 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 175 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 175 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 175 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 175 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 176 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 176 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 176 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35185740
string GDS_FILE /home/ali11-2000/FYP/mpw/UETRV-ECORE/openlane/Core/runs/Core/results/finishing/Core.magic.gds
string GDS_START 1448936
<< end >>

