VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO WB_InterConnect
  CLASS BLOCK ;
  FOREIGN WB_InterConnect ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 700.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END clock
  PIN io_dbus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END io_dbus_addr[0]
  PIN io_dbus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END io_dbus_addr[10]
  PIN io_dbus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END io_dbus_addr[11]
  PIN io_dbus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END io_dbus_addr[12]
  PIN io_dbus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END io_dbus_addr[13]
  PIN io_dbus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END io_dbus_addr[14]
  PIN io_dbus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END io_dbus_addr[15]
  PIN io_dbus_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END io_dbus_addr[16]
  PIN io_dbus_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END io_dbus_addr[17]
  PIN io_dbus_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END io_dbus_addr[18]
  PIN io_dbus_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END io_dbus_addr[19]
  PIN io_dbus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END io_dbus_addr[1]
  PIN io_dbus_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END io_dbus_addr[20]
  PIN io_dbus_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END io_dbus_addr[21]
  PIN io_dbus_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END io_dbus_addr[22]
  PIN io_dbus_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END io_dbus_addr[23]
  PIN io_dbus_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END io_dbus_addr[24]
  PIN io_dbus_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END io_dbus_addr[25]
  PIN io_dbus_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END io_dbus_addr[26]
  PIN io_dbus_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END io_dbus_addr[27]
  PIN io_dbus_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END io_dbus_addr[28]
  PIN io_dbus_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END io_dbus_addr[29]
  PIN io_dbus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END io_dbus_addr[2]
  PIN io_dbus_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END io_dbus_addr[30]
  PIN io_dbus_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END io_dbus_addr[31]
  PIN io_dbus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END io_dbus_addr[3]
  PIN io_dbus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_dbus_addr[4]
  PIN io_dbus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_dbus_addr[5]
  PIN io_dbus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END io_dbus_addr[6]
  PIN io_dbus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END io_dbus_addr[7]
  PIN io_dbus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END io_dbus_addr[8]
  PIN io_dbus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END io_dbus_addr[9]
  PIN io_dbus_ld_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END io_dbus_ld_type[0]
  PIN io_dbus_ld_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_dbus_ld_type[1]
  PIN io_dbus_ld_type[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END io_dbus_ld_type[2]
  PIN io_dbus_rd_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END io_dbus_rd_en
  PIN io_dbus_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END io_dbus_rdata[0]
  PIN io_dbus_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END io_dbus_rdata[10]
  PIN io_dbus_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END io_dbus_rdata[11]
  PIN io_dbus_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END io_dbus_rdata[12]
  PIN io_dbus_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END io_dbus_rdata[13]
  PIN io_dbus_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END io_dbus_rdata[14]
  PIN io_dbus_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END io_dbus_rdata[15]
  PIN io_dbus_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END io_dbus_rdata[16]
  PIN io_dbus_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END io_dbus_rdata[17]
  PIN io_dbus_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END io_dbus_rdata[18]
  PIN io_dbus_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END io_dbus_rdata[19]
  PIN io_dbus_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END io_dbus_rdata[1]
  PIN io_dbus_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END io_dbus_rdata[20]
  PIN io_dbus_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END io_dbus_rdata[21]
  PIN io_dbus_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END io_dbus_rdata[22]
  PIN io_dbus_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END io_dbus_rdata[23]
  PIN io_dbus_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END io_dbus_rdata[24]
  PIN io_dbus_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END io_dbus_rdata[25]
  PIN io_dbus_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END io_dbus_rdata[26]
  PIN io_dbus_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END io_dbus_rdata[27]
  PIN io_dbus_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END io_dbus_rdata[28]
  PIN io_dbus_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END io_dbus_rdata[29]
  PIN io_dbus_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END io_dbus_rdata[2]
  PIN io_dbus_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END io_dbus_rdata[30]
  PIN io_dbus_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END io_dbus_rdata[31]
  PIN io_dbus_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END io_dbus_rdata[3]
  PIN io_dbus_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END io_dbus_rdata[4]
  PIN io_dbus_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END io_dbus_rdata[5]
  PIN io_dbus_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END io_dbus_rdata[6]
  PIN io_dbus_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END io_dbus_rdata[7]
  PIN io_dbus_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END io_dbus_rdata[8]
  PIN io_dbus_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_dbus_rdata[9]
  PIN io_dbus_st_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END io_dbus_st_type[0]
  PIN io_dbus_st_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END io_dbus_st_type[1]
  PIN io_dbus_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END io_dbus_valid
  PIN io_dbus_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END io_dbus_wdata[0]
  PIN io_dbus_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END io_dbus_wdata[10]
  PIN io_dbus_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END io_dbus_wdata[11]
  PIN io_dbus_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END io_dbus_wdata[12]
  PIN io_dbus_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END io_dbus_wdata[13]
  PIN io_dbus_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END io_dbus_wdata[14]
  PIN io_dbus_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END io_dbus_wdata[15]
  PIN io_dbus_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END io_dbus_wdata[16]
  PIN io_dbus_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END io_dbus_wdata[17]
  PIN io_dbus_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 4.000 247.480 ;
    END
  END io_dbus_wdata[18]
  PIN io_dbus_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END io_dbus_wdata[19]
  PIN io_dbus_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END io_dbus_wdata[1]
  PIN io_dbus_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END io_dbus_wdata[20]
  PIN io_dbus_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END io_dbus_wdata[21]
  PIN io_dbus_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END io_dbus_wdata[22]
  PIN io_dbus_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END io_dbus_wdata[23]
  PIN io_dbus_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END io_dbus_wdata[24]
  PIN io_dbus_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END io_dbus_wdata[25]
  PIN io_dbus_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END io_dbus_wdata[26]
  PIN io_dbus_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END io_dbus_wdata[27]
  PIN io_dbus_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END io_dbus_wdata[28]
  PIN io_dbus_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END io_dbus_wdata[29]
  PIN io_dbus_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END io_dbus_wdata[2]
  PIN io_dbus_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END io_dbus_wdata[30]
  PIN io_dbus_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END io_dbus_wdata[31]
  PIN io_dbus_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END io_dbus_wdata[3]
  PIN io_dbus_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END io_dbus_wdata[4]
  PIN io_dbus_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END io_dbus_wdata[5]
  PIN io_dbus_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END io_dbus_wdata[6]
  PIN io_dbus_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END io_dbus_wdata[7]
  PIN io_dbus_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END io_dbus_wdata[8]
  PIN io_dbus_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END io_dbus_wdata[9]
  PIN io_dbus_wr_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END io_dbus_wr_en
  PIN io_dmem_io_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 696.000 16.470 700.000 ;
    END
  END io_dmem_io_addr[0]
  PIN io_dmem_io_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 696.000 42.230 700.000 ;
    END
  END io_dmem_io_addr[1]
  PIN io_dmem_io_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 696.000 67.990 700.000 ;
    END
  END io_dmem_io_addr[2]
  PIN io_dmem_io_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 696.000 94.210 700.000 ;
    END
  END io_dmem_io_addr[3]
  PIN io_dmem_io_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 696.000 119.970 700.000 ;
    END
  END io_dmem_io_addr[4]
  PIN io_dmem_io_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 696.000 139.290 700.000 ;
    END
  END io_dmem_io_addr[5]
  PIN io_dmem_io_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 696.000 159.070 700.000 ;
    END
  END io_dmem_io_addr[6]
  PIN io_dmem_io_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 696.000 178.390 700.000 ;
    END
  END io_dmem_io_addr[7]
  PIN io_dmem_io_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 696.000 3.590 700.000 ;
    END
  END io_dmem_io_cs
  PIN io_dmem_io_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 696.000 22.910 700.000 ;
    END
  END io_dmem_io_rdata[0]
  PIN io_dmem_io_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 696.000 223.930 700.000 ;
    END
  END io_dmem_io_rdata[10]
  PIN io_dmem_io_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 696.000 236.810 700.000 ;
    END
  END io_dmem_io_rdata[11]
  PIN io_dmem_io_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 696.000 249.690 700.000 ;
    END
  END io_dmem_io_rdata[12]
  PIN io_dmem_io_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 696.000 262.570 700.000 ;
    END
  END io_dmem_io_rdata[13]
  PIN io_dmem_io_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 696.000 275.450 700.000 ;
    END
  END io_dmem_io_rdata[14]
  PIN io_dmem_io_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 696.000 288.790 700.000 ;
    END
  END io_dmem_io_rdata[15]
  PIN io_dmem_io_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 696.000 301.670 700.000 ;
    END
  END io_dmem_io_rdata[16]
  PIN io_dmem_io_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 696.000 314.550 700.000 ;
    END
  END io_dmem_io_rdata[17]
  PIN io_dmem_io_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 696.000 327.430 700.000 ;
    END
  END io_dmem_io_rdata[18]
  PIN io_dmem_io_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 696.000 340.310 700.000 ;
    END
  END io_dmem_io_rdata[19]
  PIN io_dmem_io_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 696.000 48.670 700.000 ;
    END
  END io_dmem_io_rdata[1]
  PIN io_dmem_io_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 696.000 353.650 700.000 ;
    END
  END io_dmem_io_rdata[20]
  PIN io_dmem_io_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 696.000 366.530 700.000 ;
    END
  END io_dmem_io_rdata[21]
  PIN io_dmem_io_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 696.000 379.410 700.000 ;
    END
  END io_dmem_io_rdata[22]
  PIN io_dmem_io_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 696.000 392.290 700.000 ;
    END
  END io_dmem_io_rdata[23]
  PIN io_dmem_io_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 696.000 405.170 700.000 ;
    END
  END io_dmem_io_rdata[24]
  PIN io_dmem_io_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 696.000 418.050 700.000 ;
    END
  END io_dmem_io_rdata[25]
  PIN io_dmem_io_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 696.000 431.390 700.000 ;
    END
  END io_dmem_io_rdata[26]
  PIN io_dmem_io_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 696.000 444.270 700.000 ;
    END
  END io_dmem_io_rdata[27]
  PIN io_dmem_io_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 696.000 457.150 700.000 ;
    END
  END io_dmem_io_rdata[28]
  PIN io_dmem_io_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 696.000 470.030 700.000 ;
    END
  END io_dmem_io_rdata[29]
  PIN io_dmem_io_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 696.000 74.890 700.000 ;
    END
  END io_dmem_io_rdata[2]
  PIN io_dmem_io_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 696.000 482.910 700.000 ;
    END
  END io_dmem_io_rdata[30]
  PIN io_dmem_io_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 696.000 496.250 700.000 ;
    END
  END io_dmem_io_rdata[31]
  PIN io_dmem_io_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 696.000 100.650 700.000 ;
    END
  END io_dmem_io_rdata[3]
  PIN io_dmem_io_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 696.000 126.410 700.000 ;
    END
  END io_dmem_io_rdata[4]
  PIN io_dmem_io_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 696.000 146.190 700.000 ;
    END
  END io_dmem_io_rdata[5]
  PIN io_dmem_io_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 696.000 165.510 700.000 ;
    END
  END io_dmem_io_rdata[6]
  PIN io_dmem_io_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 696.000 184.830 700.000 ;
    END
  END io_dmem_io_rdata[7]
  PIN io_dmem_io_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 696.000 197.710 700.000 ;
    END
  END io_dmem_io_rdata[8]
  PIN io_dmem_io_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 696.000 210.590 700.000 ;
    END
  END io_dmem_io_rdata[9]
  PIN io_dmem_io_st_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 696.000 29.350 700.000 ;
    END
  END io_dmem_io_st_type[0]
  PIN io_dmem_io_st_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 696.000 55.110 700.000 ;
    END
  END io_dmem_io_st_type[1]
  PIN io_dmem_io_st_type[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 696.000 81.330 700.000 ;
    END
  END io_dmem_io_st_type[2]
  PIN io_dmem_io_st_type[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 696.000 107.090 700.000 ;
    END
  END io_dmem_io_st_type[3]
  PIN io_dmem_io_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 696.000 35.790 700.000 ;
    END
  END io_dmem_io_wdata[0]
  PIN io_dmem_io_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 696.000 230.370 700.000 ;
    END
  END io_dmem_io_wdata[10]
  PIN io_dmem_io_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 696.000 243.250 700.000 ;
    END
  END io_dmem_io_wdata[11]
  PIN io_dmem_io_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 696.000 256.130 700.000 ;
    END
  END io_dmem_io_wdata[12]
  PIN io_dmem_io_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 696.000 269.010 700.000 ;
    END
  END io_dmem_io_wdata[13]
  PIN io_dmem_io_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 696.000 281.890 700.000 ;
    END
  END io_dmem_io_wdata[14]
  PIN io_dmem_io_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 696.000 295.230 700.000 ;
    END
  END io_dmem_io_wdata[15]
  PIN io_dmem_io_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 696.000 308.110 700.000 ;
    END
  END io_dmem_io_wdata[16]
  PIN io_dmem_io_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 696.000 320.990 700.000 ;
    END
  END io_dmem_io_wdata[17]
  PIN io_dmem_io_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 696.000 333.870 700.000 ;
    END
  END io_dmem_io_wdata[18]
  PIN io_dmem_io_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 696.000 346.750 700.000 ;
    END
  END io_dmem_io_wdata[19]
  PIN io_dmem_io_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 696.000 61.550 700.000 ;
    END
  END io_dmem_io_wdata[1]
  PIN io_dmem_io_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 696.000 360.090 700.000 ;
    END
  END io_dmem_io_wdata[20]
  PIN io_dmem_io_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 696.000 372.970 700.000 ;
    END
  END io_dmem_io_wdata[21]
  PIN io_dmem_io_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 696.000 385.850 700.000 ;
    END
  END io_dmem_io_wdata[22]
  PIN io_dmem_io_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 696.000 398.730 700.000 ;
    END
  END io_dmem_io_wdata[23]
  PIN io_dmem_io_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 696.000 411.610 700.000 ;
    END
  END io_dmem_io_wdata[24]
  PIN io_dmem_io_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 696.000 424.950 700.000 ;
    END
  END io_dmem_io_wdata[25]
  PIN io_dmem_io_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 696.000 437.830 700.000 ;
    END
  END io_dmem_io_wdata[26]
  PIN io_dmem_io_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 696.000 450.710 700.000 ;
    END
  END io_dmem_io_wdata[27]
  PIN io_dmem_io_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 696.000 463.590 700.000 ;
    END
  END io_dmem_io_wdata[28]
  PIN io_dmem_io_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 696.000 476.470 700.000 ;
    END
  END io_dmem_io_wdata[29]
  PIN io_dmem_io_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 696.000 87.770 700.000 ;
    END
  END io_dmem_io_wdata[2]
  PIN io_dmem_io_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 696.000 489.350 700.000 ;
    END
  END io_dmem_io_wdata[30]
  PIN io_dmem_io_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 696.000 502.690 700.000 ;
    END
  END io_dmem_io_wdata[31]
  PIN io_dmem_io_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 696.000 113.530 700.000 ;
    END
  END io_dmem_io_wdata[3]
  PIN io_dmem_io_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 696.000 132.850 700.000 ;
    END
  END io_dmem_io_wdata[4]
  PIN io_dmem_io_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 696.000 152.630 700.000 ;
    END
  END io_dmem_io_wdata[5]
  PIN io_dmem_io_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 696.000 171.950 700.000 ;
    END
  END io_dmem_io_wdata[6]
  PIN io_dmem_io_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 696.000 191.270 700.000 ;
    END
  END io_dmem_io_wdata[7]
  PIN io_dmem_io_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 696.000 204.150 700.000 ;
    END
  END io_dmem_io_wdata[8]
  PIN io_dmem_io_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 696.000 217.490 700.000 ;
    END
  END io_dmem_io_wdata[9]
  PIN io_dmem_io_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 696.000 10.030 700.000 ;
    END
  END io_dmem_io_wr_en
  PIN io_ibus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END io_ibus_addr[0]
  PIN io_ibus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END io_ibus_addr[10]
  PIN io_ibus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END io_ibus_addr[11]
  PIN io_ibus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END io_ibus_addr[12]
  PIN io_ibus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END io_ibus_addr[13]
  PIN io_ibus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.080 4.000 512.680 ;
    END
  END io_ibus_addr[14]
  PIN io_ibus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END io_ibus_addr[15]
  PIN io_ibus_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END io_ibus_addr[16]
  PIN io_ibus_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END io_ibus_addr[17]
  PIN io_ibus_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END io_ibus_addr[18]
  PIN io_ibus_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END io_ibus_addr[19]
  PIN io_ibus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END io_ibus_addr[1]
  PIN io_ibus_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 558.320 4.000 558.920 ;
    END
  END io_ibus_addr[20]
  PIN io_ibus_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 4.000 567.080 ;
    END
  END io_ibus_addr[21]
  PIN io_ibus_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END io_ibus_addr[22]
  PIN io_ibus_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END io_ibus_addr[23]
  PIN io_ibus_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.600 4.000 590.200 ;
    END
  END io_ibus_addr[24]
  PIN io_ibus_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END io_ibus_addr[25]
  PIN io_ibus_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END io_ibus_addr[26]
  PIN io_ibus_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END io_ibus_addr[27]
  PIN io_ibus_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END io_ibus_addr[28]
  PIN io_ibus_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END io_ibus_addr[29]
  PIN io_ibus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END io_ibus_addr[2]
  PIN io_ibus_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END io_ibus_addr[30]
  PIN io_ibus_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END io_ibus_addr[31]
  PIN io_ibus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END io_ibus_addr[3]
  PIN io_ibus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END io_ibus_addr[4]
  PIN io_ibus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END io_ibus_addr[5]
  PIN io_ibus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.880 4.000 451.480 ;
    END
  END io_ibus_addr[6]
  PIN io_ibus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END io_ibus_addr[7]
  PIN io_ibus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END io_ibus_addr[8]
  PIN io_ibus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END io_ibus_addr[9]
  PIN io_ibus_inst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END io_ibus_inst[0]
  PIN io_ibus_inst[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END io_ibus_inst[10]
  PIN io_ibus_inst[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END io_ibus_inst[11]
  PIN io_ibus_inst[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END io_ibus_inst[12]
  PIN io_ibus_inst[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END io_ibus_inst[13]
  PIN io_ibus_inst[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.160 4.000 516.760 ;
    END
  END io_ibus_inst[14]
  PIN io_ibus_inst[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END io_ibus_inst[15]
  PIN io_ibus_inst[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END io_ibus_inst[16]
  PIN io_ibus_inst[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.280 4.000 539.880 ;
    END
  END io_ibus_inst[17]
  PIN io_ibus_inst[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END io_ibus_inst[18]
  PIN io_ibus_inst[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END io_ibus_inst[19]
  PIN io_ibus_inst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END io_ibus_inst[1]
  PIN io_ibus_inst[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END io_ibus_inst[20]
  PIN io_ibus_inst[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END io_ibus_inst[21]
  PIN io_ibus_inst[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END io_ibus_inst[22]
  PIN io_ibus_inst[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END io_ibus_inst[23]
  PIN io_ibus_inst[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END io_ibus_inst[24]
  PIN io_ibus_inst[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END io_ibus_inst[25]
  PIN io_ibus_inst[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END io_ibus_inst[26]
  PIN io_ibus_inst[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END io_ibus_inst[27]
  PIN io_ibus_inst[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END io_ibus_inst[28]
  PIN io_ibus_inst[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END io_ibus_inst[29]
  PIN io_ibus_inst[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END io_ibus_inst[2]
  PIN io_ibus_inst[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END io_ibus_inst[30]
  PIN io_ibus_inst[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END io_ibus_inst[31]
  PIN io_ibus_inst[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END io_ibus_inst[3]
  PIN io_ibus_inst[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END io_ibus_inst[4]
  PIN io_ibus_inst[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.800 4.000 447.400 ;
    END
  END io_ibus_inst[5]
  PIN io_ibus_inst[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.960 4.000 455.560 ;
    END
  END io_ibus_inst[6]
  PIN io_ibus_inst[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END io_ibus_inst[7]
  PIN io_ibus_inst[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END io_ibus_inst[8]
  PIN io_ibus_inst[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END io_ibus_inst[9]
  PIN io_ibus_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END io_ibus_valid
  PIN io_imem_io_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END io_imem_io_addr[0]
  PIN io_imem_io_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 696.000 515.570 700.000 ;
    END
  END io_imem_io_addr[1]
  PIN io_imem_io_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 696.000 522.010 700.000 ;
    END
  END io_imem_io_addr[2]
  PIN io_imem_io_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 606.600 700.000 607.200 ;
    END
  END io_imem_io_addr[3]
  PIN io_imem_io_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 696.000 541.330 700.000 ;
    END
  END io_imem_io_addr[4]
  PIN io_imem_io_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END io_imem_io_addr[5]
  PIN io_imem_io_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 696.000 560.650 700.000 ;
    END
  END io_imem_io_addr[6]
  PIN io_imem_io_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END io_imem_io_addr[7]
  PIN io_imem_io_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END io_imem_io_addr[8]
  PIN io_imem_io_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 587.560 700.000 588.160 ;
    END
  END io_imem_io_cs
  PIN io_imem_io_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END io_imem_io_rdata[0]
  PIN io_imem_io_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 644.680 700.000 645.280 ;
    END
  END io_imem_io_rdata[10]
  PIN io_imem_io_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 696.000 573.990 700.000 ;
    END
  END io_imem_io_rdata[11]
  PIN io_imem_io_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 696.000 580.430 700.000 ;
    END
  END io_imem_io_rdata[12]
  PIN io_imem_io_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 696.000 586.870 700.000 ;
    END
  END io_imem_io_rdata[13]
  PIN io_imem_io_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END io_imem_io_rdata[14]
  PIN io_imem_io_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 696.000 599.750 700.000 ;
    END
  END io_imem_io_rdata[15]
  PIN io_imem_io_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 696.000 612.630 700.000 ;
    END
  END io_imem_io_rdata[16]
  PIN io_imem_io_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END io_imem_io_rdata[17]
  PIN io_imem_io_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 670.520 700.000 671.120 ;
    END
  END io_imem_io_rdata[18]
  PIN io_imem_io_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 696.000 619.070 700.000 ;
    END
  END io_imem_io_rdata[19]
  PIN io_imem_io_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 593.680 700.000 594.280 ;
    END
  END io_imem_io_rdata[1]
  PIN io_imem_io_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 682.760 700.000 683.360 ;
    END
  END io_imem_io_rdata[20]
  PIN io_imem_io_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 696.000 631.950 700.000 ;
    END
  END io_imem_io_rdata[21]
  PIN io_imem_io_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END io_imem_io_rdata[22]
  PIN io_imem_io_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 689.560 700.000 690.160 ;
    END
  END io_imem_io_rdata[23]
  PIN io_imem_io_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 696.000 658.170 700.000 ;
    END
  END io_imem_io_rdata[24]
  PIN io_imem_io_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END io_imem_io_rdata[25]
  PIN io_imem_io_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.960 4.000 693.560 ;
    END
  END io_imem_io_rdata[26]
  PIN io_imem_io_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 695.680 700.000 696.280 ;
    END
  END io_imem_io_rdata[27]
  PIN io_imem_io_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END io_imem_io_rdata[28]
  PIN io_imem_io_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 696.000 677.490 700.000 ;
    END
  END io_imem_io_rdata[29]
  PIN io_imem_io_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 696.000 528.450 700.000 ;
    END
  END io_imem_io_rdata[2]
  PIN io_imem_io_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END io_imem_io_rdata[30]
  PIN io_imem_io_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 696.000 696.810 700.000 ;
    END
  END io_imem_io_rdata[31]
  PIN io_imem_io_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END io_imem_io_rdata[3]
  PIN io_imem_io_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 696.000 547.770 700.000 ;
    END
  END io_imem_io_rdata[4]
  PIN io_imem_io_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END io_imem_io_rdata[5]
  PIN io_imem_io_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 625.640 700.000 626.240 ;
    END
  END io_imem_io_rdata[6]
  PIN io_imem_io_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 632.440 700.000 633.040 ;
    END
  END io_imem_io_rdata[7]
  PIN io_imem_io_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END io_imem_io_rdata[8]
  PIN io_imem_io_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 696.000 567.550 700.000 ;
    END
  END io_imem_io_rdata[9]
  PIN io_imem_io_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END io_imem_io_wdata[0]
  PIN io_imem_io_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 651.480 700.000 652.080 ;
    END
  END io_imem_io_wdata[10]
  PIN io_imem_io_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END io_imem_io_wdata[11]
  PIN io_imem_io_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 657.600 700.000 658.200 ;
    END
  END io_imem_io_wdata[12]
  PIN io_imem_io_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 696.000 593.310 700.000 ;
    END
  END io_imem_io_wdata[13]
  PIN io_imem_io_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 663.720 700.000 664.320 ;
    END
  END io_imem_io_wdata[14]
  PIN io_imem_io_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 696.000 606.190 700.000 ;
    END
  END io_imem_io_wdata[15]
  PIN io_imem_io_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END io_imem_io_wdata[16]
  PIN io_imem_io_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END io_imem_io_wdata[17]
  PIN io_imem_io_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 676.640 700.000 677.240 ;
    END
  END io_imem_io_wdata[18]
  PIN io_imem_io_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END io_imem_io_wdata[19]
  PIN io_imem_io_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 600.480 700.000 601.080 ;
    END
  END io_imem_io_wdata[1]
  PIN io_imem_io_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 696.000 625.510 700.000 ;
    END
  END io_imem_io_wdata[20]
  PIN io_imem_io_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 696.000 638.850 700.000 ;
    END
  END io_imem_io_wdata[21]
  PIN io_imem_io_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 696.000 645.290 700.000 ;
    END
  END io_imem_io_wdata[22]
  PIN io_imem_io_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 696.000 651.730 700.000 ;
    END
  END io_imem_io_wdata[23]
  PIN io_imem_io_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 696.000 664.610 700.000 ;
    END
  END io_imem_io_wdata[24]
  PIN io_imem_io_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END io_imem_io_wdata[25]
  PIN io_imem_io_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 696.000 671.050 700.000 ;
    END
  END io_imem_io_wdata[26]
  PIN io_imem_io_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END io_imem_io_wdata[27]
  PIN io_imem_io_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END io_imem_io_wdata[28]
  PIN io_imem_io_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 696.000 683.930 700.000 ;
    END
  END io_imem_io_wdata[29]
  PIN io_imem_io_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 696.000 534.890 700.000 ;
    END
  END io_imem_io_wdata[2]
  PIN io_imem_io_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 696.000 690.370 700.000 ;
    END
  END io_imem_io_wdata[30]
  PIN io_imem_io_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END io_imem_io_wdata[31]
  PIN io_imem_io_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 613.400 700.000 614.000 ;
    END
  END io_imem_io_wdata[3]
  PIN io_imem_io_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 619.520 700.000 620.120 ;
    END
  END io_imem_io_wdata[4]
  PIN io_imem_io_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 696.000 554.210 700.000 ;
    END
  END io_imem_io_wdata[5]
  PIN io_imem_io_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END io_imem_io_wdata[6]
  PIN io_imem_io_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END io_imem_io_wdata[7]
  PIN io_imem_io_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 638.560 700.000 639.160 ;
    END
  END io_imem_io_wdata[8]
  PIN io_imem_io_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END io_imem_io_wdata[9]
  PIN io_imem_io_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 696.000 509.130 700.000 ;
    END
  END io_imem_io_wr_en
  PIN io_motor_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 2.760 700.000 3.360 ;
    END
  END io_motor_ack_i
  PIN io_motor_addr_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 8.880 700.000 9.480 ;
    END
  END io_motor_addr_sel
  PIN io_motor_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 15.000 700.000 15.600 ;
    END
  END io_motor_data_i[0]
  PIN io_motor_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 78.920 700.000 79.520 ;
    END
  END io_motor_data_i[10]
  PIN io_motor_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 85.040 700.000 85.640 ;
    END
  END io_motor_data_i[11]
  PIN io_motor_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 91.160 700.000 91.760 ;
    END
  END io_motor_data_i[12]
  PIN io_motor_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 97.960 700.000 98.560 ;
    END
  END io_motor_data_i[13]
  PIN io_motor_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 104.080 700.000 104.680 ;
    END
  END io_motor_data_i[14]
  PIN io_motor_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 110.880 700.000 111.480 ;
    END
  END io_motor_data_i[15]
  PIN io_motor_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 117.000 700.000 117.600 ;
    END
  END io_motor_data_i[16]
  PIN io_motor_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 123.120 700.000 123.720 ;
    END
  END io_motor_data_i[17]
  PIN io_motor_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 129.920 700.000 130.520 ;
    END
  END io_motor_data_i[18]
  PIN io_motor_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 136.040 700.000 136.640 ;
    END
  END io_motor_data_i[19]
  PIN io_motor_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 21.800 700.000 22.400 ;
    END
  END io_motor_data_i[1]
  PIN io_motor_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 142.160 700.000 142.760 ;
    END
  END io_motor_data_i[20]
  PIN io_motor_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 148.960 700.000 149.560 ;
    END
  END io_motor_data_i[21]
  PIN io_motor_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 155.080 700.000 155.680 ;
    END
  END io_motor_data_i[22]
  PIN io_motor_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 161.200 700.000 161.800 ;
    END
  END io_motor_data_i[23]
  PIN io_motor_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 168.000 700.000 168.600 ;
    END
  END io_motor_data_i[24]
  PIN io_motor_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 174.120 700.000 174.720 ;
    END
  END io_motor_data_i[25]
  PIN io_motor_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 180.240 700.000 180.840 ;
    END
  END io_motor_data_i[26]
  PIN io_motor_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 187.040 700.000 187.640 ;
    END
  END io_motor_data_i[27]
  PIN io_motor_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 193.160 700.000 193.760 ;
    END
  END io_motor_data_i[28]
  PIN io_motor_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 199.280 700.000 199.880 ;
    END
  END io_motor_data_i[29]
  PIN io_motor_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 27.920 700.000 28.520 ;
    END
  END io_motor_data_i[2]
  PIN io_motor_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 206.080 700.000 206.680 ;
    END
  END io_motor_data_i[30]
  PIN io_motor_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 212.200 700.000 212.800 ;
    END
  END io_motor_data_i[31]
  PIN io_motor_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 34.040 700.000 34.640 ;
    END
  END io_motor_data_i[3]
  PIN io_motor_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 40.840 700.000 41.440 ;
    END
  END io_motor_data_i[4]
  PIN io_motor_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 46.960 700.000 47.560 ;
    END
  END io_motor_data_i[5]
  PIN io_motor_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 53.080 700.000 53.680 ;
    END
  END io_motor_data_i[6]
  PIN io_motor_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 59.880 700.000 60.480 ;
    END
  END io_motor_data_i[7]
  PIN io_motor_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 66.000 700.000 66.600 ;
    END
  END io_motor_data_i[8]
  PIN io_motor_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 72.120 700.000 72.720 ;
    END
  END io_motor_data_i[9]
  PIN io_spi_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 562.400 700.000 563.000 ;
    END
  END io_spi_clk
  PIN io_spi_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 568.520 700.000 569.120 ;
    END
  END io_spi_cs
  PIN io_spi_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END io_spi_irq
  PIN io_spi_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_spi_miso
  PIN io_spi_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 574.640 700.000 575.240 ;
    END
  END io_spi_mosi
  PIN io_uart_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.880 4.000 655.480 ;
    END
  END io_uart_irq
  PIN io_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END io_uart_rx
  PIN io_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 581.440 700.000 582.040 ;
    END
  END io_uart_tx
  PIN io_wbm_m2s_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 231.240 700.000 231.840 ;
    END
  END io_wbm_m2s_addr[0]
  PIN io_wbm_m2s_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 384.240 700.000 384.840 ;
    END
  END io_wbm_m2s_addr[10]
  PIN io_wbm_m2s_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 396.480 700.000 397.080 ;
    END
  END io_wbm_m2s_addr[11]
  PIN io_wbm_m2s_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 409.400 700.000 410.000 ;
    END
  END io_wbm_m2s_addr[12]
  PIN io_wbm_m2s_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 422.320 700.000 422.920 ;
    END
  END io_wbm_m2s_addr[13]
  PIN io_wbm_m2s_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 435.240 700.000 435.840 ;
    END
  END io_wbm_m2s_addr[14]
  PIN io_wbm_m2s_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 447.480 700.000 448.080 ;
    END
  END io_wbm_m2s_addr[15]
  PIN io_wbm_m2s_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 250.280 700.000 250.880 ;
    END
  END io_wbm_m2s_addr[1]
  PIN io_wbm_m2s_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 269.320 700.000 269.920 ;
    END
  END io_wbm_m2s_addr[2]
  PIN io_wbm_m2s_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 288.360 700.000 288.960 ;
    END
  END io_wbm_m2s_addr[3]
  PIN io_wbm_m2s_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 308.080 700.000 308.680 ;
    END
  END io_wbm_m2s_addr[4]
  PIN io_wbm_m2s_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 320.320 700.000 320.920 ;
    END
  END io_wbm_m2s_addr[5]
  PIN io_wbm_m2s_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 333.240 700.000 333.840 ;
    END
  END io_wbm_m2s_addr[6]
  PIN io_wbm_m2s_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 346.160 700.000 346.760 ;
    END
  END io_wbm_m2s_addr[7]
  PIN io_wbm_m2s_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 358.400 700.000 359.000 ;
    END
  END io_wbm_m2s_addr[8]
  PIN io_wbm_m2s_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 371.320 700.000 371.920 ;
    END
  END io_wbm_m2s_addr[9]
  PIN io_wbm_m2s_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 238.040 700.000 238.640 ;
    END
  END io_wbm_m2s_data[0]
  PIN io_wbm_m2s_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 390.360 700.000 390.960 ;
    END
  END io_wbm_m2s_data[10]
  PIN io_wbm_m2s_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 403.280 700.000 403.880 ;
    END
  END io_wbm_m2s_data[11]
  PIN io_wbm_m2s_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 416.200 700.000 416.800 ;
    END
  END io_wbm_m2s_data[12]
  PIN io_wbm_m2s_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 428.440 700.000 429.040 ;
    END
  END io_wbm_m2s_data[13]
  PIN io_wbm_m2s_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 441.360 700.000 441.960 ;
    END
  END io_wbm_m2s_data[14]
  PIN io_wbm_m2s_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 454.280 700.000 454.880 ;
    END
  END io_wbm_m2s_data[15]
  PIN io_wbm_m2s_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 460.400 700.000 461.000 ;
    END
  END io_wbm_m2s_data[16]
  PIN io_wbm_m2s_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 466.520 700.000 467.120 ;
    END
  END io_wbm_m2s_data[17]
  PIN io_wbm_m2s_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 473.320 700.000 473.920 ;
    END
  END io_wbm_m2s_data[18]
  PIN io_wbm_m2s_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 479.440 700.000 480.040 ;
    END
  END io_wbm_m2s_data[19]
  PIN io_wbm_m2s_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 257.080 700.000 257.680 ;
    END
  END io_wbm_m2s_data[1]
  PIN io_wbm_m2s_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 485.560 700.000 486.160 ;
    END
  END io_wbm_m2s_data[20]
  PIN io_wbm_m2s_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 492.360 700.000 492.960 ;
    END
  END io_wbm_m2s_data[21]
  PIN io_wbm_m2s_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 498.480 700.000 499.080 ;
    END
  END io_wbm_m2s_data[22]
  PIN io_wbm_m2s_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 505.280 700.000 505.880 ;
    END
  END io_wbm_m2s_data[23]
  PIN io_wbm_m2s_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 511.400 700.000 512.000 ;
    END
  END io_wbm_m2s_data[24]
  PIN io_wbm_m2s_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 517.520 700.000 518.120 ;
    END
  END io_wbm_m2s_data[25]
  PIN io_wbm_m2s_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 524.320 700.000 524.920 ;
    END
  END io_wbm_m2s_data[26]
  PIN io_wbm_m2s_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 530.440 700.000 531.040 ;
    END
  END io_wbm_m2s_data[27]
  PIN io_wbm_m2s_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 536.560 700.000 537.160 ;
    END
  END io_wbm_m2s_data[28]
  PIN io_wbm_m2s_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 543.360 700.000 543.960 ;
    END
  END io_wbm_m2s_data[29]
  PIN io_wbm_m2s_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 276.120 700.000 276.720 ;
    END
  END io_wbm_m2s_data[2]
  PIN io_wbm_m2s_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 549.480 700.000 550.080 ;
    END
  END io_wbm_m2s_data[30]
  PIN io_wbm_m2s_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 555.600 700.000 556.200 ;
    END
  END io_wbm_m2s_data[31]
  PIN io_wbm_m2s_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 295.160 700.000 295.760 ;
    END
  END io_wbm_m2s_data[3]
  PIN io_wbm_m2s_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 314.200 700.000 314.800 ;
    END
  END io_wbm_m2s_data[4]
  PIN io_wbm_m2s_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 327.120 700.000 327.720 ;
    END
  END io_wbm_m2s_data[5]
  PIN io_wbm_m2s_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 339.360 700.000 339.960 ;
    END
  END io_wbm_m2s_data[6]
  PIN io_wbm_m2s_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 352.280 700.000 352.880 ;
    END
  END io_wbm_m2s_data[7]
  PIN io_wbm_m2s_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 365.200 700.000 365.800 ;
    END
  END io_wbm_m2s_data[8]
  PIN io_wbm_m2s_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 377.440 700.000 378.040 ;
    END
  END io_wbm_m2s_data[9]
  PIN io_wbm_m2s_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 244.160 700.000 244.760 ;
    END
  END io_wbm_m2s_sel[0]
  PIN io_wbm_m2s_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 263.200 700.000 263.800 ;
    END
  END io_wbm_m2s_sel[1]
  PIN io_wbm_m2s_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 282.240 700.000 282.840 ;
    END
  END io_wbm_m2s_sel[2]
  PIN io_wbm_m2s_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 301.280 700.000 301.880 ;
    END
  END io_wbm_m2s_sel[3]
  PIN io_wbm_m2s_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 219.000 700.000 219.600 ;
    END
  END io_wbm_m2s_stb
  PIN io_wbm_m2s_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 225.120 700.000 225.720 ;
    END
  END io_wbm_m2s_we
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 688.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 688.400 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 694.140 688.245 ;
      LAYER met1 ;
        RECT 5.130 10.640 696.830 689.140 ;
      LAYER met2 ;
        RECT 3.870 695.720 9.470 697.525 ;
        RECT 10.310 695.720 15.910 697.525 ;
        RECT 16.750 695.720 22.350 697.525 ;
        RECT 23.190 695.720 28.790 697.525 ;
        RECT 29.630 695.720 35.230 697.525 ;
        RECT 36.070 695.720 41.670 697.525 ;
        RECT 42.510 695.720 48.110 697.525 ;
        RECT 48.950 695.720 54.550 697.525 ;
        RECT 55.390 695.720 60.990 697.525 ;
        RECT 61.830 695.720 67.430 697.525 ;
        RECT 68.270 695.720 74.330 697.525 ;
        RECT 75.170 695.720 80.770 697.525 ;
        RECT 81.610 695.720 87.210 697.525 ;
        RECT 88.050 695.720 93.650 697.525 ;
        RECT 94.490 695.720 100.090 697.525 ;
        RECT 100.930 695.720 106.530 697.525 ;
        RECT 107.370 695.720 112.970 697.525 ;
        RECT 113.810 695.720 119.410 697.525 ;
        RECT 120.250 695.720 125.850 697.525 ;
        RECT 126.690 695.720 132.290 697.525 ;
        RECT 133.130 695.720 138.730 697.525 ;
        RECT 139.570 695.720 145.630 697.525 ;
        RECT 146.470 695.720 152.070 697.525 ;
        RECT 152.910 695.720 158.510 697.525 ;
        RECT 159.350 695.720 164.950 697.525 ;
        RECT 165.790 695.720 171.390 697.525 ;
        RECT 172.230 695.720 177.830 697.525 ;
        RECT 178.670 695.720 184.270 697.525 ;
        RECT 185.110 695.720 190.710 697.525 ;
        RECT 191.550 695.720 197.150 697.525 ;
        RECT 197.990 695.720 203.590 697.525 ;
        RECT 204.430 695.720 210.030 697.525 ;
        RECT 210.870 695.720 216.930 697.525 ;
        RECT 217.770 695.720 223.370 697.525 ;
        RECT 224.210 695.720 229.810 697.525 ;
        RECT 230.650 695.720 236.250 697.525 ;
        RECT 237.090 695.720 242.690 697.525 ;
        RECT 243.530 695.720 249.130 697.525 ;
        RECT 249.970 695.720 255.570 697.525 ;
        RECT 256.410 695.720 262.010 697.525 ;
        RECT 262.850 695.720 268.450 697.525 ;
        RECT 269.290 695.720 274.890 697.525 ;
        RECT 275.730 695.720 281.330 697.525 ;
        RECT 282.170 695.720 288.230 697.525 ;
        RECT 289.070 695.720 294.670 697.525 ;
        RECT 295.510 695.720 301.110 697.525 ;
        RECT 301.950 695.720 307.550 697.525 ;
        RECT 308.390 695.720 313.990 697.525 ;
        RECT 314.830 695.720 320.430 697.525 ;
        RECT 321.270 695.720 326.870 697.525 ;
        RECT 327.710 695.720 333.310 697.525 ;
        RECT 334.150 695.720 339.750 697.525 ;
        RECT 340.590 695.720 346.190 697.525 ;
        RECT 347.030 695.720 353.090 697.525 ;
        RECT 353.930 695.720 359.530 697.525 ;
        RECT 360.370 695.720 365.970 697.525 ;
        RECT 366.810 695.720 372.410 697.525 ;
        RECT 373.250 695.720 378.850 697.525 ;
        RECT 379.690 695.720 385.290 697.525 ;
        RECT 386.130 695.720 391.730 697.525 ;
        RECT 392.570 695.720 398.170 697.525 ;
        RECT 399.010 695.720 404.610 697.525 ;
        RECT 405.450 695.720 411.050 697.525 ;
        RECT 411.890 695.720 417.490 697.525 ;
        RECT 418.330 695.720 424.390 697.525 ;
        RECT 425.230 695.720 430.830 697.525 ;
        RECT 431.670 695.720 437.270 697.525 ;
        RECT 438.110 695.720 443.710 697.525 ;
        RECT 444.550 695.720 450.150 697.525 ;
        RECT 450.990 695.720 456.590 697.525 ;
        RECT 457.430 695.720 463.030 697.525 ;
        RECT 463.870 695.720 469.470 697.525 ;
        RECT 470.310 695.720 475.910 697.525 ;
        RECT 476.750 695.720 482.350 697.525 ;
        RECT 483.190 695.720 488.790 697.525 ;
        RECT 489.630 695.720 495.690 697.525 ;
        RECT 496.530 695.720 502.130 697.525 ;
        RECT 502.970 695.720 508.570 697.525 ;
        RECT 509.410 695.720 515.010 697.525 ;
        RECT 515.850 695.720 521.450 697.525 ;
        RECT 522.290 695.720 527.890 697.525 ;
        RECT 528.730 695.720 534.330 697.525 ;
        RECT 535.170 695.720 540.770 697.525 ;
        RECT 541.610 695.720 547.210 697.525 ;
        RECT 548.050 695.720 553.650 697.525 ;
        RECT 554.490 695.720 560.090 697.525 ;
        RECT 560.930 695.720 566.990 697.525 ;
        RECT 567.830 695.720 573.430 697.525 ;
        RECT 574.270 695.720 579.870 697.525 ;
        RECT 580.710 695.720 586.310 697.525 ;
        RECT 587.150 695.720 592.750 697.525 ;
        RECT 593.590 695.720 599.190 697.525 ;
        RECT 600.030 695.720 605.630 697.525 ;
        RECT 606.470 695.720 612.070 697.525 ;
        RECT 612.910 695.720 618.510 697.525 ;
        RECT 619.350 695.720 624.950 697.525 ;
        RECT 625.790 695.720 631.390 697.525 ;
        RECT 632.230 695.720 638.290 697.525 ;
        RECT 639.130 695.720 644.730 697.525 ;
        RECT 645.570 695.720 651.170 697.525 ;
        RECT 652.010 695.720 657.610 697.525 ;
        RECT 658.450 695.720 664.050 697.525 ;
        RECT 664.890 695.720 670.490 697.525 ;
        RECT 671.330 695.720 676.930 697.525 ;
        RECT 677.770 695.720 683.370 697.525 ;
        RECT 684.210 695.720 689.810 697.525 ;
        RECT 690.650 695.720 696.250 697.525 ;
        RECT 3.590 4.280 696.800 695.720 ;
        RECT 3.590 1.515 17.290 4.280 ;
        RECT 18.130 1.515 52.250 4.280 ;
        RECT 53.090 1.515 87.210 4.280 ;
        RECT 88.050 1.515 122.170 4.280 ;
        RECT 123.010 1.515 157.130 4.280 ;
        RECT 157.970 1.515 192.090 4.280 ;
        RECT 192.930 1.515 227.050 4.280 ;
        RECT 227.890 1.515 262.010 4.280 ;
        RECT 262.850 1.515 296.970 4.280 ;
        RECT 297.810 1.515 331.930 4.280 ;
        RECT 332.770 1.515 367.350 4.280 ;
        RECT 368.190 1.515 402.310 4.280 ;
        RECT 403.150 1.515 437.270 4.280 ;
        RECT 438.110 1.515 472.230 4.280 ;
        RECT 473.070 1.515 507.190 4.280 ;
        RECT 508.030 1.515 542.150 4.280 ;
        RECT 542.990 1.515 577.110 4.280 ;
        RECT 577.950 1.515 612.070 4.280 ;
        RECT 612.910 1.515 647.030 4.280 ;
        RECT 647.870 1.515 681.990 4.280 ;
        RECT 682.830 1.515 696.800 4.280 ;
      LAYER met3 ;
        RECT 4.400 696.680 696.000 697.505 ;
        RECT 4.400 696.640 695.600 696.680 ;
        RECT 4.000 695.280 695.600 696.640 ;
        RECT 4.000 693.960 696.000 695.280 ;
        RECT 4.400 692.560 696.000 693.960 ;
        RECT 4.000 690.560 696.000 692.560 ;
        RECT 4.400 689.160 695.600 690.560 ;
        RECT 4.000 686.480 696.000 689.160 ;
        RECT 4.400 685.080 696.000 686.480 ;
        RECT 4.000 683.760 696.000 685.080 ;
        RECT 4.000 682.400 695.600 683.760 ;
        RECT 4.400 682.360 695.600 682.400 ;
        RECT 4.400 681.000 696.000 682.360 ;
        RECT 4.000 679.000 696.000 681.000 ;
        RECT 4.400 677.640 696.000 679.000 ;
        RECT 4.400 677.600 695.600 677.640 ;
        RECT 4.000 676.240 695.600 677.600 ;
        RECT 4.000 674.920 696.000 676.240 ;
        RECT 4.400 673.520 696.000 674.920 ;
        RECT 4.000 671.520 696.000 673.520 ;
        RECT 4.000 670.840 695.600 671.520 ;
        RECT 4.400 670.120 695.600 670.840 ;
        RECT 4.400 669.440 696.000 670.120 ;
        RECT 4.000 667.440 696.000 669.440 ;
        RECT 4.400 666.040 696.000 667.440 ;
        RECT 4.000 664.720 696.000 666.040 ;
        RECT 4.000 663.360 695.600 664.720 ;
        RECT 4.400 663.320 695.600 663.360 ;
        RECT 4.400 661.960 696.000 663.320 ;
        RECT 4.000 659.280 696.000 661.960 ;
        RECT 4.400 658.600 696.000 659.280 ;
        RECT 4.400 657.880 695.600 658.600 ;
        RECT 4.000 657.200 695.600 657.880 ;
        RECT 4.000 655.880 696.000 657.200 ;
        RECT 4.400 654.480 696.000 655.880 ;
        RECT 4.000 652.480 696.000 654.480 ;
        RECT 4.000 651.800 695.600 652.480 ;
        RECT 4.400 651.080 695.600 651.800 ;
        RECT 4.400 650.400 696.000 651.080 ;
        RECT 4.000 647.720 696.000 650.400 ;
        RECT 4.400 646.320 696.000 647.720 ;
        RECT 4.000 645.680 696.000 646.320 ;
        RECT 4.000 644.320 695.600 645.680 ;
        RECT 4.400 644.280 695.600 644.320 ;
        RECT 4.400 642.920 696.000 644.280 ;
        RECT 4.000 640.240 696.000 642.920 ;
        RECT 4.400 639.560 696.000 640.240 ;
        RECT 4.400 638.840 695.600 639.560 ;
        RECT 4.000 638.160 695.600 638.840 ;
        RECT 4.000 636.160 696.000 638.160 ;
        RECT 4.400 634.760 696.000 636.160 ;
        RECT 4.000 633.440 696.000 634.760 ;
        RECT 4.000 632.760 695.600 633.440 ;
        RECT 4.400 632.040 695.600 632.760 ;
        RECT 4.400 631.360 696.000 632.040 ;
        RECT 4.000 628.680 696.000 631.360 ;
        RECT 4.400 627.280 696.000 628.680 ;
        RECT 4.000 626.640 696.000 627.280 ;
        RECT 4.000 625.240 695.600 626.640 ;
        RECT 4.000 624.600 696.000 625.240 ;
        RECT 4.400 623.200 696.000 624.600 ;
        RECT 4.000 621.200 696.000 623.200 ;
        RECT 4.400 620.520 696.000 621.200 ;
        RECT 4.400 619.800 695.600 620.520 ;
        RECT 4.000 619.120 695.600 619.800 ;
        RECT 4.000 617.120 696.000 619.120 ;
        RECT 4.400 615.720 696.000 617.120 ;
        RECT 4.000 614.400 696.000 615.720 ;
        RECT 4.000 613.040 695.600 614.400 ;
        RECT 4.400 613.000 695.600 613.040 ;
        RECT 4.400 611.640 696.000 613.000 ;
        RECT 4.000 609.640 696.000 611.640 ;
        RECT 4.400 608.240 696.000 609.640 ;
        RECT 4.000 607.600 696.000 608.240 ;
        RECT 4.000 606.200 695.600 607.600 ;
        RECT 4.000 605.560 696.000 606.200 ;
        RECT 4.400 604.160 696.000 605.560 ;
        RECT 4.000 602.160 696.000 604.160 ;
        RECT 4.400 601.480 696.000 602.160 ;
        RECT 4.400 600.760 695.600 601.480 ;
        RECT 4.000 600.080 695.600 600.760 ;
        RECT 4.000 598.080 696.000 600.080 ;
        RECT 4.400 596.680 696.000 598.080 ;
        RECT 4.000 594.680 696.000 596.680 ;
        RECT 4.000 594.000 695.600 594.680 ;
        RECT 4.400 593.280 695.600 594.000 ;
        RECT 4.400 592.600 696.000 593.280 ;
        RECT 4.000 590.600 696.000 592.600 ;
        RECT 4.400 589.200 696.000 590.600 ;
        RECT 4.000 588.560 696.000 589.200 ;
        RECT 4.000 587.160 695.600 588.560 ;
        RECT 4.000 586.520 696.000 587.160 ;
        RECT 4.400 585.120 696.000 586.520 ;
        RECT 4.000 582.440 696.000 585.120 ;
        RECT 4.400 581.040 695.600 582.440 ;
        RECT 4.000 579.040 696.000 581.040 ;
        RECT 4.400 577.640 696.000 579.040 ;
        RECT 4.000 575.640 696.000 577.640 ;
        RECT 4.000 574.960 695.600 575.640 ;
        RECT 4.400 574.240 695.600 574.960 ;
        RECT 4.400 573.560 696.000 574.240 ;
        RECT 4.000 570.880 696.000 573.560 ;
        RECT 4.400 569.520 696.000 570.880 ;
        RECT 4.400 569.480 695.600 569.520 ;
        RECT 4.000 568.120 695.600 569.480 ;
        RECT 4.000 567.480 696.000 568.120 ;
        RECT 4.400 566.080 696.000 567.480 ;
        RECT 4.000 563.400 696.000 566.080 ;
        RECT 4.400 562.000 695.600 563.400 ;
        RECT 4.000 559.320 696.000 562.000 ;
        RECT 4.400 557.920 696.000 559.320 ;
        RECT 4.000 556.600 696.000 557.920 ;
        RECT 4.000 555.920 695.600 556.600 ;
        RECT 4.400 555.200 695.600 555.920 ;
        RECT 4.400 554.520 696.000 555.200 ;
        RECT 4.000 551.840 696.000 554.520 ;
        RECT 4.400 550.480 696.000 551.840 ;
        RECT 4.400 550.440 695.600 550.480 ;
        RECT 4.000 549.080 695.600 550.440 ;
        RECT 4.000 547.760 696.000 549.080 ;
        RECT 4.400 546.360 696.000 547.760 ;
        RECT 4.000 544.360 696.000 546.360 ;
        RECT 4.400 542.960 695.600 544.360 ;
        RECT 4.000 540.280 696.000 542.960 ;
        RECT 4.400 538.880 696.000 540.280 ;
        RECT 4.000 537.560 696.000 538.880 ;
        RECT 4.000 536.200 695.600 537.560 ;
        RECT 4.400 536.160 695.600 536.200 ;
        RECT 4.400 534.800 696.000 536.160 ;
        RECT 4.000 532.800 696.000 534.800 ;
        RECT 4.400 531.440 696.000 532.800 ;
        RECT 4.400 531.400 695.600 531.440 ;
        RECT 4.000 530.040 695.600 531.400 ;
        RECT 4.000 528.720 696.000 530.040 ;
        RECT 4.400 527.320 696.000 528.720 ;
        RECT 4.000 525.320 696.000 527.320 ;
        RECT 4.000 524.640 695.600 525.320 ;
        RECT 4.400 523.920 695.600 524.640 ;
        RECT 4.400 523.240 696.000 523.920 ;
        RECT 4.000 521.240 696.000 523.240 ;
        RECT 4.400 519.840 696.000 521.240 ;
        RECT 4.000 518.520 696.000 519.840 ;
        RECT 4.000 517.160 695.600 518.520 ;
        RECT 4.400 517.120 695.600 517.160 ;
        RECT 4.400 515.760 696.000 517.120 ;
        RECT 4.000 513.080 696.000 515.760 ;
        RECT 4.400 512.400 696.000 513.080 ;
        RECT 4.400 511.680 695.600 512.400 ;
        RECT 4.000 511.000 695.600 511.680 ;
        RECT 4.000 509.680 696.000 511.000 ;
        RECT 4.400 508.280 696.000 509.680 ;
        RECT 4.000 506.280 696.000 508.280 ;
        RECT 4.000 505.600 695.600 506.280 ;
        RECT 4.400 504.880 695.600 505.600 ;
        RECT 4.400 504.200 696.000 504.880 ;
        RECT 4.000 502.200 696.000 504.200 ;
        RECT 4.400 500.800 696.000 502.200 ;
        RECT 4.000 499.480 696.000 500.800 ;
        RECT 4.000 498.120 695.600 499.480 ;
        RECT 4.400 498.080 695.600 498.120 ;
        RECT 4.400 496.720 696.000 498.080 ;
        RECT 4.000 494.040 696.000 496.720 ;
        RECT 4.400 493.360 696.000 494.040 ;
        RECT 4.400 492.640 695.600 493.360 ;
        RECT 4.000 491.960 695.600 492.640 ;
        RECT 4.000 490.640 696.000 491.960 ;
        RECT 4.400 489.240 696.000 490.640 ;
        RECT 4.000 486.560 696.000 489.240 ;
        RECT 4.400 485.160 695.600 486.560 ;
        RECT 4.000 482.480 696.000 485.160 ;
        RECT 4.400 481.080 696.000 482.480 ;
        RECT 4.000 480.440 696.000 481.080 ;
        RECT 4.000 479.080 695.600 480.440 ;
        RECT 4.400 479.040 695.600 479.080 ;
        RECT 4.400 477.680 696.000 479.040 ;
        RECT 4.000 475.000 696.000 477.680 ;
        RECT 4.400 474.320 696.000 475.000 ;
        RECT 4.400 473.600 695.600 474.320 ;
        RECT 4.000 472.920 695.600 473.600 ;
        RECT 4.000 470.920 696.000 472.920 ;
        RECT 4.400 469.520 696.000 470.920 ;
        RECT 4.000 467.520 696.000 469.520 ;
        RECT 4.400 466.120 695.600 467.520 ;
        RECT 4.000 463.440 696.000 466.120 ;
        RECT 4.400 462.040 696.000 463.440 ;
        RECT 4.000 461.400 696.000 462.040 ;
        RECT 4.000 460.000 695.600 461.400 ;
        RECT 4.000 459.360 696.000 460.000 ;
        RECT 4.400 457.960 696.000 459.360 ;
        RECT 4.000 455.960 696.000 457.960 ;
        RECT 4.400 455.280 696.000 455.960 ;
        RECT 4.400 454.560 695.600 455.280 ;
        RECT 4.000 453.880 695.600 454.560 ;
        RECT 4.000 451.880 696.000 453.880 ;
        RECT 4.400 450.480 696.000 451.880 ;
        RECT 4.000 448.480 696.000 450.480 ;
        RECT 4.000 447.800 695.600 448.480 ;
        RECT 4.400 447.080 695.600 447.800 ;
        RECT 4.400 446.400 696.000 447.080 ;
        RECT 4.000 444.400 696.000 446.400 ;
        RECT 4.400 443.000 696.000 444.400 ;
        RECT 4.000 442.360 696.000 443.000 ;
        RECT 4.000 440.960 695.600 442.360 ;
        RECT 4.000 440.320 696.000 440.960 ;
        RECT 4.400 438.920 696.000 440.320 ;
        RECT 4.000 436.240 696.000 438.920 ;
        RECT 4.400 434.840 695.600 436.240 ;
        RECT 4.000 432.840 696.000 434.840 ;
        RECT 4.400 431.440 696.000 432.840 ;
        RECT 4.000 429.440 696.000 431.440 ;
        RECT 4.000 428.760 695.600 429.440 ;
        RECT 4.400 428.040 695.600 428.760 ;
        RECT 4.400 427.360 696.000 428.040 ;
        RECT 4.000 424.680 696.000 427.360 ;
        RECT 4.400 423.320 696.000 424.680 ;
        RECT 4.400 423.280 695.600 423.320 ;
        RECT 4.000 421.920 695.600 423.280 ;
        RECT 4.000 421.280 696.000 421.920 ;
        RECT 4.400 419.880 696.000 421.280 ;
        RECT 4.000 417.200 696.000 419.880 ;
        RECT 4.400 415.800 695.600 417.200 ;
        RECT 4.000 413.120 696.000 415.800 ;
        RECT 4.400 411.720 696.000 413.120 ;
        RECT 4.000 410.400 696.000 411.720 ;
        RECT 4.000 409.720 695.600 410.400 ;
        RECT 4.400 409.000 695.600 409.720 ;
        RECT 4.400 408.320 696.000 409.000 ;
        RECT 4.000 405.640 696.000 408.320 ;
        RECT 4.400 404.280 696.000 405.640 ;
        RECT 4.400 404.240 695.600 404.280 ;
        RECT 4.000 402.880 695.600 404.240 ;
        RECT 4.000 402.240 696.000 402.880 ;
        RECT 4.400 400.840 696.000 402.240 ;
        RECT 4.000 398.160 696.000 400.840 ;
        RECT 4.400 397.480 696.000 398.160 ;
        RECT 4.400 396.760 695.600 397.480 ;
        RECT 4.000 396.080 695.600 396.760 ;
        RECT 4.000 394.080 696.000 396.080 ;
        RECT 4.400 392.680 696.000 394.080 ;
        RECT 4.000 391.360 696.000 392.680 ;
        RECT 4.000 390.680 695.600 391.360 ;
        RECT 4.400 389.960 695.600 390.680 ;
        RECT 4.400 389.280 696.000 389.960 ;
        RECT 4.000 386.600 696.000 389.280 ;
        RECT 4.400 385.240 696.000 386.600 ;
        RECT 4.400 385.200 695.600 385.240 ;
        RECT 4.000 383.840 695.600 385.200 ;
        RECT 4.000 382.520 696.000 383.840 ;
        RECT 4.400 381.120 696.000 382.520 ;
        RECT 4.000 379.120 696.000 381.120 ;
        RECT 4.400 378.440 696.000 379.120 ;
        RECT 4.400 377.720 695.600 378.440 ;
        RECT 4.000 377.040 695.600 377.720 ;
        RECT 4.000 375.040 696.000 377.040 ;
        RECT 4.400 373.640 696.000 375.040 ;
        RECT 4.000 372.320 696.000 373.640 ;
        RECT 4.000 370.960 695.600 372.320 ;
        RECT 4.400 370.920 695.600 370.960 ;
        RECT 4.400 369.560 696.000 370.920 ;
        RECT 4.000 367.560 696.000 369.560 ;
        RECT 4.400 366.200 696.000 367.560 ;
        RECT 4.400 366.160 695.600 366.200 ;
        RECT 4.000 364.800 695.600 366.160 ;
        RECT 4.000 363.480 696.000 364.800 ;
        RECT 4.400 362.080 696.000 363.480 ;
        RECT 4.000 359.400 696.000 362.080 ;
        RECT 4.400 358.000 695.600 359.400 ;
        RECT 4.000 356.000 696.000 358.000 ;
        RECT 4.400 354.600 696.000 356.000 ;
        RECT 4.000 353.280 696.000 354.600 ;
        RECT 4.000 351.920 695.600 353.280 ;
        RECT 4.400 351.880 695.600 351.920 ;
        RECT 4.400 350.520 696.000 351.880 ;
        RECT 4.000 347.840 696.000 350.520 ;
        RECT 4.400 347.160 696.000 347.840 ;
        RECT 4.400 346.440 695.600 347.160 ;
        RECT 4.000 345.760 695.600 346.440 ;
        RECT 4.000 344.440 696.000 345.760 ;
        RECT 4.400 343.040 696.000 344.440 ;
        RECT 4.000 340.360 696.000 343.040 ;
        RECT 4.400 338.960 695.600 340.360 ;
        RECT 4.000 336.280 696.000 338.960 ;
        RECT 4.400 334.880 696.000 336.280 ;
        RECT 4.000 334.240 696.000 334.880 ;
        RECT 4.000 332.880 695.600 334.240 ;
        RECT 4.400 332.840 695.600 332.880 ;
        RECT 4.400 331.480 696.000 332.840 ;
        RECT 4.000 328.800 696.000 331.480 ;
        RECT 4.400 328.120 696.000 328.800 ;
        RECT 4.400 327.400 695.600 328.120 ;
        RECT 4.000 326.720 695.600 327.400 ;
        RECT 4.000 324.720 696.000 326.720 ;
        RECT 4.400 323.320 696.000 324.720 ;
        RECT 4.000 321.320 696.000 323.320 ;
        RECT 4.400 319.920 695.600 321.320 ;
        RECT 4.000 317.240 696.000 319.920 ;
        RECT 4.400 315.840 696.000 317.240 ;
        RECT 4.000 315.200 696.000 315.840 ;
        RECT 4.000 313.800 695.600 315.200 ;
        RECT 4.000 313.160 696.000 313.800 ;
        RECT 4.400 311.760 696.000 313.160 ;
        RECT 4.000 309.760 696.000 311.760 ;
        RECT 4.400 309.080 696.000 309.760 ;
        RECT 4.400 308.360 695.600 309.080 ;
        RECT 4.000 307.680 695.600 308.360 ;
        RECT 4.000 305.680 696.000 307.680 ;
        RECT 4.400 304.280 696.000 305.680 ;
        RECT 4.000 302.280 696.000 304.280 ;
        RECT 4.400 300.880 695.600 302.280 ;
        RECT 4.000 298.200 696.000 300.880 ;
        RECT 4.400 296.800 696.000 298.200 ;
        RECT 4.000 296.160 696.000 296.800 ;
        RECT 4.000 294.760 695.600 296.160 ;
        RECT 4.000 294.120 696.000 294.760 ;
        RECT 4.400 292.720 696.000 294.120 ;
        RECT 4.000 290.720 696.000 292.720 ;
        RECT 4.400 289.360 696.000 290.720 ;
        RECT 4.400 289.320 695.600 289.360 ;
        RECT 4.000 287.960 695.600 289.320 ;
        RECT 4.000 286.640 696.000 287.960 ;
        RECT 4.400 285.240 696.000 286.640 ;
        RECT 4.000 283.240 696.000 285.240 ;
        RECT 4.000 282.560 695.600 283.240 ;
        RECT 4.400 281.840 695.600 282.560 ;
        RECT 4.400 281.160 696.000 281.840 ;
        RECT 4.000 279.160 696.000 281.160 ;
        RECT 4.400 277.760 696.000 279.160 ;
        RECT 4.000 277.120 696.000 277.760 ;
        RECT 4.000 275.720 695.600 277.120 ;
        RECT 4.000 275.080 696.000 275.720 ;
        RECT 4.400 273.680 696.000 275.080 ;
        RECT 4.000 271.000 696.000 273.680 ;
        RECT 4.400 270.320 696.000 271.000 ;
        RECT 4.400 269.600 695.600 270.320 ;
        RECT 4.000 268.920 695.600 269.600 ;
        RECT 4.000 267.600 696.000 268.920 ;
        RECT 4.400 266.200 696.000 267.600 ;
        RECT 4.000 264.200 696.000 266.200 ;
        RECT 4.000 263.520 695.600 264.200 ;
        RECT 4.400 262.800 695.600 263.520 ;
        RECT 4.400 262.120 696.000 262.800 ;
        RECT 4.000 259.440 696.000 262.120 ;
        RECT 4.400 258.080 696.000 259.440 ;
        RECT 4.400 258.040 695.600 258.080 ;
        RECT 4.000 256.680 695.600 258.040 ;
        RECT 4.000 256.040 696.000 256.680 ;
        RECT 4.400 254.640 696.000 256.040 ;
        RECT 4.000 251.960 696.000 254.640 ;
        RECT 4.400 251.280 696.000 251.960 ;
        RECT 4.400 250.560 695.600 251.280 ;
        RECT 4.000 249.880 695.600 250.560 ;
        RECT 4.000 247.880 696.000 249.880 ;
        RECT 4.400 246.480 696.000 247.880 ;
        RECT 4.000 245.160 696.000 246.480 ;
        RECT 4.000 244.480 695.600 245.160 ;
        RECT 4.400 243.760 695.600 244.480 ;
        RECT 4.400 243.080 696.000 243.760 ;
        RECT 4.000 240.400 696.000 243.080 ;
        RECT 4.400 239.040 696.000 240.400 ;
        RECT 4.400 239.000 695.600 239.040 ;
        RECT 4.000 237.640 695.600 239.000 ;
        RECT 4.000 236.320 696.000 237.640 ;
        RECT 4.400 234.920 696.000 236.320 ;
        RECT 4.000 232.920 696.000 234.920 ;
        RECT 4.400 232.240 696.000 232.920 ;
        RECT 4.400 231.520 695.600 232.240 ;
        RECT 4.000 230.840 695.600 231.520 ;
        RECT 4.000 228.840 696.000 230.840 ;
        RECT 4.400 227.440 696.000 228.840 ;
        RECT 4.000 226.120 696.000 227.440 ;
        RECT 4.000 224.760 695.600 226.120 ;
        RECT 4.400 224.720 695.600 224.760 ;
        RECT 4.400 223.360 696.000 224.720 ;
        RECT 4.000 221.360 696.000 223.360 ;
        RECT 4.400 220.000 696.000 221.360 ;
        RECT 4.400 219.960 695.600 220.000 ;
        RECT 4.000 218.600 695.600 219.960 ;
        RECT 4.000 217.280 696.000 218.600 ;
        RECT 4.400 215.880 696.000 217.280 ;
        RECT 4.000 213.200 696.000 215.880 ;
        RECT 4.400 211.800 695.600 213.200 ;
        RECT 4.000 209.800 696.000 211.800 ;
        RECT 4.400 208.400 696.000 209.800 ;
        RECT 4.000 207.080 696.000 208.400 ;
        RECT 4.000 205.720 695.600 207.080 ;
        RECT 4.400 205.680 695.600 205.720 ;
        RECT 4.400 204.320 696.000 205.680 ;
        RECT 4.000 202.320 696.000 204.320 ;
        RECT 4.400 200.920 696.000 202.320 ;
        RECT 4.000 200.280 696.000 200.920 ;
        RECT 4.000 198.880 695.600 200.280 ;
        RECT 4.000 198.240 696.000 198.880 ;
        RECT 4.400 196.840 696.000 198.240 ;
        RECT 4.000 194.160 696.000 196.840 ;
        RECT 4.400 192.760 695.600 194.160 ;
        RECT 4.000 190.760 696.000 192.760 ;
        RECT 4.400 189.360 696.000 190.760 ;
        RECT 4.000 188.040 696.000 189.360 ;
        RECT 4.000 186.680 695.600 188.040 ;
        RECT 4.400 186.640 695.600 186.680 ;
        RECT 4.400 185.280 696.000 186.640 ;
        RECT 4.000 182.600 696.000 185.280 ;
        RECT 4.400 181.240 696.000 182.600 ;
        RECT 4.400 181.200 695.600 181.240 ;
        RECT 4.000 179.840 695.600 181.200 ;
        RECT 4.000 179.200 696.000 179.840 ;
        RECT 4.400 177.800 696.000 179.200 ;
        RECT 4.000 175.120 696.000 177.800 ;
        RECT 4.400 173.720 695.600 175.120 ;
        RECT 4.000 171.040 696.000 173.720 ;
        RECT 4.400 169.640 696.000 171.040 ;
        RECT 4.000 169.000 696.000 169.640 ;
        RECT 4.000 167.640 695.600 169.000 ;
        RECT 4.400 167.600 695.600 167.640 ;
        RECT 4.400 166.240 696.000 167.600 ;
        RECT 4.000 163.560 696.000 166.240 ;
        RECT 4.400 162.200 696.000 163.560 ;
        RECT 4.400 162.160 695.600 162.200 ;
        RECT 4.000 160.800 695.600 162.160 ;
        RECT 4.000 159.480 696.000 160.800 ;
        RECT 4.400 158.080 696.000 159.480 ;
        RECT 4.000 156.080 696.000 158.080 ;
        RECT 4.400 154.680 695.600 156.080 ;
        RECT 4.000 152.000 696.000 154.680 ;
        RECT 4.400 150.600 696.000 152.000 ;
        RECT 4.000 149.960 696.000 150.600 ;
        RECT 4.000 148.560 695.600 149.960 ;
        RECT 4.000 147.920 696.000 148.560 ;
        RECT 4.400 146.520 696.000 147.920 ;
        RECT 4.000 144.520 696.000 146.520 ;
        RECT 4.400 143.160 696.000 144.520 ;
        RECT 4.400 143.120 695.600 143.160 ;
        RECT 4.000 141.760 695.600 143.120 ;
        RECT 4.000 140.440 696.000 141.760 ;
        RECT 4.400 139.040 696.000 140.440 ;
        RECT 4.000 137.040 696.000 139.040 ;
        RECT 4.000 136.360 695.600 137.040 ;
        RECT 4.400 135.640 695.600 136.360 ;
        RECT 4.400 134.960 696.000 135.640 ;
        RECT 4.000 132.960 696.000 134.960 ;
        RECT 4.400 131.560 696.000 132.960 ;
        RECT 4.000 130.920 696.000 131.560 ;
        RECT 4.000 129.520 695.600 130.920 ;
        RECT 4.000 128.880 696.000 129.520 ;
        RECT 4.400 127.480 696.000 128.880 ;
        RECT 4.000 124.800 696.000 127.480 ;
        RECT 4.400 124.120 696.000 124.800 ;
        RECT 4.400 123.400 695.600 124.120 ;
        RECT 4.000 122.720 695.600 123.400 ;
        RECT 4.000 121.400 696.000 122.720 ;
        RECT 4.400 120.000 696.000 121.400 ;
        RECT 4.000 118.000 696.000 120.000 ;
        RECT 4.000 117.320 695.600 118.000 ;
        RECT 4.400 116.600 695.600 117.320 ;
        RECT 4.400 115.920 696.000 116.600 ;
        RECT 4.000 113.240 696.000 115.920 ;
        RECT 4.400 111.880 696.000 113.240 ;
        RECT 4.400 111.840 695.600 111.880 ;
        RECT 4.000 110.480 695.600 111.840 ;
        RECT 4.000 109.840 696.000 110.480 ;
        RECT 4.400 108.440 696.000 109.840 ;
        RECT 4.000 105.760 696.000 108.440 ;
        RECT 4.400 105.080 696.000 105.760 ;
        RECT 4.400 104.360 695.600 105.080 ;
        RECT 4.000 103.680 695.600 104.360 ;
        RECT 4.000 102.360 696.000 103.680 ;
        RECT 4.400 100.960 696.000 102.360 ;
        RECT 4.000 98.960 696.000 100.960 ;
        RECT 4.000 98.280 695.600 98.960 ;
        RECT 4.400 97.560 695.600 98.280 ;
        RECT 4.400 96.880 696.000 97.560 ;
        RECT 4.000 94.200 696.000 96.880 ;
        RECT 4.400 92.800 696.000 94.200 ;
        RECT 4.000 92.160 696.000 92.800 ;
        RECT 4.000 90.800 695.600 92.160 ;
        RECT 4.400 90.760 695.600 90.800 ;
        RECT 4.400 89.400 696.000 90.760 ;
        RECT 4.000 86.720 696.000 89.400 ;
        RECT 4.400 86.040 696.000 86.720 ;
        RECT 4.400 85.320 695.600 86.040 ;
        RECT 4.000 84.640 695.600 85.320 ;
        RECT 4.000 82.640 696.000 84.640 ;
        RECT 4.400 81.240 696.000 82.640 ;
        RECT 4.000 79.920 696.000 81.240 ;
        RECT 4.000 79.240 695.600 79.920 ;
        RECT 4.400 78.520 695.600 79.240 ;
        RECT 4.400 77.840 696.000 78.520 ;
        RECT 4.000 75.160 696.000 77.840 ;
        RECT 4.400 73.760 696.000 75.160 ;
        RECT 4.000 73.120 696.000 73.760 ;
        RECT 4.000 71.720 695.600 73.120 ;
        RECT 4.000 71.080 696.000 71.720 ;
        RECT 4.400 69.680 696.000 71.080 ;
        RECT 4.000 67.680 696.000 69.680 ;
        RECT 4.400 67.000 696.000 67.680 ;
        RECT 4.400 66.280 695.600 67.000 ;
        RECT 4.000 65.600 695.600 66.280 ;
        RECT 4.000 63.600 696.000 65.600 ;
        RECT 4.400 62.200 696.000 63.600 ;
        RECT 4.000 60.880 696.000 62.200 ;
        RECT 4.000 59.520 695.600 60.880 ;
        RECT 4.400 59.480 695.600 59.520 ;
        RECT 4.400 58.120 696.000 59.480 ;
        RECT 4.000 56.120 696.000 58.120 ;
        RECT 4.400 54.720 696.000 56.120 ;
        RECT 4.000 54.080 696.000 54.720 ;
        RECT 4.000 52.680 695.600 54.080 ;
        RECT 4.000 52.040 696.000 52.680 ;
        RECT 4.400 50.640 696.000 52.040 ;
        RECT 4.000 47.960 696.000 50.640 ;
        RECT 4.400 46.560 695.600 47.960 ;
        RECT 4.000 44.560 696.000 46.560 ;
        RECT 4.400 43.160 696.000 44.560 ;
        RECT 4.000 41.840 696.000 43.160 ;
        RECT 4.000 40.480 695.600 41.840 ;
        RECT 4.400 40.440 695.600 40.480 ;
        RECT 4.400 39.080 696.000 40.440 ;
        RECT 4.000 36.400 696.000 39.080 ;
        RECT 4.400 35.040 696.000 36.400 ;
        RECT 4.400 35.000 695.600 35.040 ;
        RECT 4.000 33.640 695.600 35.000 ;
        RECT 4.000 33.000 696.000 33.640 ;
        RECT 4.400 31.600 696.000 33.000 ;
        RECT 4.000 28.920 696.000 31.600 ;
        RECT 4.400 27.520 695.600 28.920 ;
        RECT 4.000 24.840 696.000 27.520 ;
        RECT 4.400 23.440 696.000 24.840 ;
        RECT 4.000 22.800 696.000 23.440 ;
        RECT 4.000 21.440 695.600 22.800 ;
        RECT 4.400 21.400 695.600 21.440 ;
        RECT 4.400 20.040 696.000 21.400 ;
        RECT 4.000 17.360 696.000 20.040 ;
        RECT 4.400 16.000 696.000 17.360 ;
        RECT 4.400 15.960 695.600 16.000 ;
        RECT 4.000 14.600 695.600 15.960 ;
        RECT 4.000 13.280 696.000 14.600 ;
        RECT 4.400 11.880 696.000 13.280 ;
        RECT 4.000 9.880 696.000 11.880 ;
        RECT 4.400 8.480 695.600 9.880 ;
        RECT 4.000 5.800 696.000 8.480 ;
        RECT 4.400 4.400 696.000 5.800 ;
        RECT 4.000 3.760 696.000 4.400 ;
        RECT 4.000 2.400 695.600 3.760 ;
        RECT 4.400 2.360 695.600 2.400 ;
        RECT 4.400 1.535 696.000 2.360 ;
      LAYER met4 ;
        RECT 12.255 11.735 20.640 685.945 ;
        RECT 23.040 11.735 97.440 685.945 ;
        RECT 99.840 11.735 174.240 685.945 ;
        RECT 176.640 11.735 225.105 685.945 ;
  END
END WB_InterConnect
END LIBRARY

