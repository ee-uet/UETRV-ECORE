VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Core
  CLASS BLOCK ;
  FOREIGN Core ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 496.000 125.030 500.000 ;
    END
  END clock
  PIN io_dbus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 9.560 500.000 10.160 ;
    END
  END io_dbus_addr[0]
  PIN io_dbus_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 111.560 500.000 112.160 ;
    END
  END io_dbus_addr[10]
  PIN io_dbus_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 120.400 500.000 121.000 ;
    END
  END io_dbus_addr[11]
  PIN io_dbus_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 129.240 500.000 129.840 ;
    END
  END io_dbus_addr[12]
  PIN io_dbus_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 137.400 500.000 138.000 ;
    END
  END io_dbus_addr[13]
  PIN io_dbus_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 146.240 500.000 146.840 ;
    END
  END io_dbus_addr[14]
  PIN io_dbus_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 155.080 500.000 155.680 ;
    END
  END io_dbus_addr[15]
  PIN io_dbus_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 163.920 500.000 164.520 ;
    END
  END io_dbus_addr[16]
  PIN io_dbus_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 172.760 500.000 173.360 ;
    END
  END io_dbus_addr[17]
  PIN io_dbus_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 180.920 500.000 181.520 ;
    END
  END io_dbus_addr[18]
  PIN io_dbus_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 189.760 500.000 190.360 ;
    END
  END io_dbus_addr[19]
  PIN io_dbus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 24.520 500.000 25.120 ;
    END
  END io_dbus_addr[1]
  PIN io_dbus_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 198.600 500.000 199.200 ;
    END
  END io_dbus_addr[20]
  PIN io_dbus_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 207.440 500.000 208.040 ;
    END
  END io_dbus_addr[21]
  PIN io_dbus_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 216.280 500.000 216.880 ;
    END
  END io_dbus_addr[22]
  PIN io_dbus_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 225.120 500.000 225.720 ;
    END
  END io_dbus_addr[23]
  PIN io_dbus_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 233.280 500.000 233.880 ;
    END
  END io_dbus_addr[24]
  PIN io_dbus_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 242.120 500.000 242.720 ;
    END
  END io_dbus_addr[25]
  PIN io_dbus_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 250.960 500.000 251.560 ;
    END
  END io_dbus_addr[26]
  PIN io_dbus_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 259.800 500.000 260.400 ;
    END
  END io_dbus_addr[27]
  PIN io_dbus_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 268.640 500.000 269.240 ;
    END
  END io_dbus_addr[28]
  PIN io_dbus_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 276.800 500.000 277.400 ;
    END
  END io_dbus_addr[29]
  PIN io_dbus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 38.800 500.000 39.400 ;
    END
  END io_dbus_addr[2]
  PIN io_dbus_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 285.640 500.000 286.240 ;
    END
  END io_dbus_addr[30]
  PIN io_dbus_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 294.480 500.000 295.080 ;
    END
  END io_dbus_addr[31]
  PIN io_dbus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 50.360 500.000 50.960 ;
    END
  END io_dbus_addr[3]
  PIN io_dbus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 59.200 500.000 59.800 ;
    END
  END io_dbus_addr[4]
  PIN io_dbus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 68.040 500.000 68.640 ;
    END
  END io_dbus_addr[5]
  PIN io_dbus_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 76.880 500.000 77.480 ;
    END
  END io_dbus_addr[6]
  PIN io_dbus_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 85.040 500.000 85.640 ;
    END
  END io_dbus_addr[7]
  PIN io_dbus_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 93.880 500.000 94.480 ;
    END
  END io_dbus_addr[8]
  PIN io_dbus_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 102.720 500.000 103.320 ;
    END
  END io_dbus_addr[9]
  PIN io_dbus_ld_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 12.960 500.000 13.560 ;
    END
  END io_dbus_ld_type[0]
  PIN io_dbus_ld_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 27.240 500.000 27.840 ;
    END
  END io_dbus_ld_type[1]
  PIN io_dbus_ld_type[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 41.520 500.000 42.120 ;
    END
  END io_dbus_ld_type[2]
  PIN io_dbus_rd_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 1.400 500.000 2.000 ;
    END
  END io_dbus_rd_en
  PIN io_dbus_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 15.680 500.000 16.280 ;
    END
  END io_dbus_rdata[0]
  PIN io_dbus_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 114.280 500.000 114.880 ;
    END
  END io_dbus_rdata[10]
  PIN io_dbus_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 123.120 500.000 123.720 ;
    END
  END io_dbus_rdata[11]
  PIN io_dbus_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 131.960 500.000 132.560 ;
    END
  END io_dbus_rdata[12]
  PIN io_dbus_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 140.800 500.000 141.400 ;
    END
  END io_dbus_rdata[13]
  PIN io_dbus_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 148.960 500.000 149.560 ;
    END
  END io_dbus_rdata[14]
  PIN io_dbus_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 157.800 500.000 158.400 ;
    END
  END io_dbus_rdata[15]
  PIN io_dbus_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 166.640 500.000 167.240 ;
    END
  END io_dbus_rdata[16]
  PIN io_dbus_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 175.480 500.000 176.080 ;
    END
  END io_dbus_rdata[17]
  PIN io_dbus_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 184.320 500.000 184.920 ;
    END
  END io_dbus_rdata[18]
  PIN io_dbus_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 193.160 500.000 193.760 ;
    END
  END io_dbus_rdata[19]
  PIN io_dbus_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 29.960 500.000 30.560 ;
    END
  END io_dbus_rdata[1]
  PIN io_dbus_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 201.320 500.000 201.920 ;
    END
  END io_dbus_rdata[20]
  PIN io_dbus_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.160 500.000 210.760 ;
    END
  END io_dbus_rdata[21]
  PIN io_dbus_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 219.000 500.000 219.600 ;
    END
  END io_dbus_rdata[22]
  PIN io_dbus_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 227.840 500.000 228.440 ;
    END
  END io_dbus_rdata[23]
  PIN io_dbus_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 236.680 500.000 237.280 ;
    END
  END io_dbus_rdata[24]
  PIN io_dbus_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 244.840 500.000 245.440 ;
    END
  END io_dbus_rdata[25]
  PIN io_dbus_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 253.680 500.000 254.280 ;
    END
  END io_dbus_rdata[26]
  PIN io_dbus_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 262.520 500.000 263.120 ;
    END
  END io_dbus_rdata[27]
  PIN io_dbus_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 271.360 500.000 271.960 ;
    END
  END io_dbus_rdata[28]
  PIN io_dbus_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 280.200 500.000 280.800 ;
    END
  END io_dbus_rdata[29]
  PIN io_dbus_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.920 500.000 45.520 ;
    END
  END io_dbus_rdata[2]
  PIN io_dbus_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 289.040 500.000 289.640 ;
    END
  END io_dbus_rdata[30]
  PIN io_dbus_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 297.200 500.000 297.800 ;
    END
  END io_dbus_rdata[31]
  PIN io_dbus_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 53.080 500.000 53.680 ;
    END
  END io_dbus_rdata[3]
  PIN io_dbus_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 61.920 500.000 62.520 ;
    END
  END io_dbus_rdata[4]
  PIN io_dbus_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 70.760 500.000 71.360 ;
    END
  END io_dbus_rdata[5]
  PIN io_dbus_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 79.600 500.000 80.200 ;
    END
  END io_dbus_rdata[6]
  PIN io_dbus_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 88.440 500.000 89.040 ;
    END
  END io_dbus_rdata[7]
  PIN io_dbus_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 97.280 500.000 97.880 ;
    END
  END io_dbus_rdata[8]
  PIN io_dbus_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 105.440 500.000 106.040 ;
    END
  END io_dbus_rdata[9]
  PIN io_dbus_st_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 18.400 500.000 19.000 ;
    END
  END io_dbus_st_type[0]
  PIN io_dbus_st_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 33.360 500.000 33.960 ;
    END
  END io_dbus_st_type[1]
  PIN io_dbus_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 4.120 500.000 4.720 ;
    END
  END io_dbus_valid
  PIN io_dbus_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 21.120 500.000 21.720 ;
    END
  END io_dbus_wdata[0]
  PIN io_dbus_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 117.000 500.000 117.600 ;
    END
  END io_dbus_wdata[10]
  PIN io_dbus_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 125.840 500.000 126.440 ;
    END
  END io_dbus_wdata[11]
  PIN io_dbus_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 134.680 500.000 135.280 ;
    END
  END io_dbus_wdata[12]
  PIN io_dbus_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 143.520 500.000 144.120 ;
    END
  END io_dbus_wdata[13]
  PIN io_dbus_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 152.360 500.000 152.960 ;
    END
  END io_dbus_wdata[14]
  PIN io_dbus_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 161.200 500.000 161.800 ;
    END
  END io_dbus_wdata[15]
  PIN io_dbus_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 169.360 500.000 169.960 ;
    END
  END io_dbus_wdata[16]
  PIN io_dbus_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 178.200 500.000 178.800 ;
    END
  END io_dbus_wdata[17]
  PIN io_dbus_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 187.040 500.000 187.640 ;
    END
  END io_dbus_wdata[18]
  PIN io_dbus_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 195.880 500.000 196.480 ;
    END
  END io_dbus_wdata[19]
  PIN io_dbus_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 36.080 500.000 36.680 ;
    END
  END io_dbus_wdata[1]
  PIN io_dbus_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 204.720 500.000 205.320 ;
    END
  END io_dbus_wdata[20]
  PIN io_dbus_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 212.880 500.000 213.480 ;
    END
  END io_dbus_wdata[21]
  PIN io_dbus_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 221.720 500.000 222.320 ;
    END
  END io_dbus_wdata[22]
  PIN io_dbus_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 230.560 500.000 231.160 ;
    END
  END io_dbus_wdata[23]
  PIN io_dbus_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 239.400 500.000 240.000 ;
    END
  END io_dbus_wdata[24]
  PIN io_dbus_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 248.240 500.000 248.840 ;
    END
  END io_dbus_wdata[25]
  PIN io_dbus_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 257.080 500.000 257.680 ;
    END
  END io_dbus_wdata[26]
  PIN io_dbus_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 265.240 500.000 265.840 ;
    END
  END io_dbus_wdata[27]
  PIN io_dbus_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 274.080 500.000 274.680 ;
    END
  END io_dbus_wdata[28]
  PIN io_dbus_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 282.920 500.000 283.520 ;
    END
  END io_dbus_wdata[29]
  PIN io_dbus_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 47.640 500.000 48.240 ;
    END
  END io_dbus_wdata[2]
  PIN io_dbus_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 291.760 500.000 292.360 ;
    END
  END io_dbus_wdata[30]
  PIN io_dbus_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 300.600 500.000 301.200 ;
    END
  END io_dbus_wdata[31]
  PIN io_dbus_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 56.480 500.000 57.080 ;
    END
  END io_dbus_wdata[3]
  PIN io_dbus_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 65.320 500.000 65.920 ;
    END
  END io_dbus_wdata[4]
  PIN io_dbus_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 73.480 500.000 74.080 ;
    END
  END io_dbus_wdata[5]
  PIN io_dbus_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 82.320 500.000 82.920 ;
    END
  END io_dbus_wdata[6]
  PIN io_dbus_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 91.160 500.000 91.760 ;
    END
  END io_dbus_wdata[7]
  PIN io_dbus_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 100.000 500.000 100.600 ;
    END
  END io_dbus_wdata[8]
  PIN io_dbus_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 108.840 500.000 109.440 ;
    END
  END io_dbus_wdata[9]
  PIN io_dbus_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 6.840 500.000 7.440 ;
    END
  END io_dbus_wr_en
  PIN io_ibus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 306.040 500.000 306.640 ;
    END
  END io_ibus_addr[0]
  PIN io_ibus_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 364.520 500.000 365.120 ;
    END
  END io_ibus_addr[10]
  PIN io_ibus_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 369.960 500.000 370.560 ;
    END
  END io_ibus_addr[11]
  PIN io_ibus_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 376.080 500.000 376.680 ;
    END
  END io_ibus_addr[12]
  PIN io_ibus_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 381.520 500.000 382.120 ;
    END
  END io_ibus_addr[13]
  PIN io_ibus_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 387.640 500.000 388.240 ;
    END
  END io_ibus_addr[14]
  PIN io_ibus_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 393.080 500.000 393.680 ;
    END
  END io_ibus_addr[15]
  PIN io_ibus_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 399.200 500.000 399.800 ;
    END
  END io_ibus_addr[16]
  PIN io_ibus_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 404.640 500.000 405.240 ;
    END
  END io_ibus_addr[17]
  PIN io_ibus_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 410.760 500.000 411.360 ;
    END
  END io_ibus_addr[18]
  PIN io_ibus_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 416.880 500.000 417.480 ;
    END
  END io_ibus_addr[19]
  PIN io_ibus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 312.160 500.000 312.760 ;
    END
  END io_ibus_addr[1]
  PIN io_ibus_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 422.320 500.000 422.920 ;
    END
  END io_ibus_addr[20]
  PIN io_ibus_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 428.440 500.000 429.040 ;
    END
  END io_ibus_addr[21]
  PIN io_ibus_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 433.880 500.000 434.480 ;
    END
  END io_ibus_addr[22]
  PIN io_ibus_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 440.000 500.000 440.600 ;
    END
  END io_ibus_addr[23]
  PIN io_ibus_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 445.440 500.000 446.040 ;
    END
  END io_ibus_addr[24]
  PIN io_ibus_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 451.560 500.000 452.160 ;
    END
  END io_ibus_addr[25]
  PIN io_ibus_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 457.000 500.000 457.600 ;
    END
  END io_ibus_addr[26]
  PIN io_ibus_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 463.120 500.000 463.720 ;
    END
  END io_ibus_addr[27]
  PIN io_ibus_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 468.560 500.000 469.160 ;
    END
  END io_ibus_addr[28]
  PIN io_ibus_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 474.680 500.000 475.280 ;
    END
  END io_ibus_addr[29]
  PIN io_ibus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 317.600 500.000 318.200 ;
    END
  END io_ibus_addr[2]
  PIN io_ibus_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 480.800 500.000 481.400 ;
    END
  END io_ibus_addr[30]
  PIN io_ibus_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 486.240 500.000 486.840 ;
    END
  END io_ibus_addr[31]
  PIN io_ibus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 323.720 500.000 324.320 ;
    END
  END io_ibus_addr[3]
  PIN io_ibus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 329.160 500.000 329.760 ;
    END
  END io_ibus_addr[4]
  PIN io_ibus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 335.280 500.000 335.880 ;
    END
  END io_ibus_addr[5]
  PIN io_ibus_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.720 500.000 341.320 ;
    END
  END io_ibus_addr[6]
  PIN io_ibus_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 346.840 500.000 347.440 ;
    END
  END io_ibus_addr[7]
  PIN io_ibus_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 352.960 500.000 353.560 ;
    END
  END io_ibus_addr[8]
  PIN io_ibus_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 358.400 500.000 359.000 ;
    END
  END io_ibus_addr[9]
  PIN io_ibus_inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 308.760 500.000 309.360 ;
    END
  END io_ibus_inst[0]
  PIN io_ibus_inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 367.240 500.000 367.840 ;
    END
  END io_ibus_inst[10]
  PIN io_ibus_inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 372.680 500.000 373.280 ;
    END
  END io_ibus_inst[11]
  PIN io_ibus_inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 378.800 500.000 379.400 ;
    END
  END io_ibus_inst[12]
  PIN io_ibus_inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 384.920 500.000 385.520 ;
    END
  END io_ibus_inst[13]
  PIN io_ibus_inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 390.360 500.000 390.960 ;
    END
  END io_ibus_inst[14]
  PIN io_ibus_inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 396.480 500.000 397.080 ;
    END
  END io_ibus_inst[15]
  PIN io_ibus_inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 401.920 500.000 402.520 ;
    END
  END io_ibus_inst[16]
  PIN io_ibus_inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 408.040 500.000 408.640 ;
    END
  END io_ibus_inst[17]
  PIN io_ibus_inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 413.480 500.000 414.080 ;
    END
  END io_ibus_inst[18]
  PIN io_ibus_inst[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 419.600 500.000 420.200 ;
    END
  END io_ibus_inst[19]
  PIN io_ibus_inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 314.880 500.000 315.480 ;
    END
  END io_ibus_inst[1]
  PIN io_ibus_inst[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 425.040 500.000 425.640 ;
    END
  END io_ibus_inst[20]
  PIN io_ibus_inst[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 431.160 500.000 431.760 ;
    END
  END io_ibus_inst[21]
  PIN io_ibus_inst[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 436.600 500.000 437.200 ;
    END
  END io_ibus_inst[22]
  PIN io_ibus_inst[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 442.720 500.000 443.320 ;
    END
  END io_ibus_inst[23]
  PIN io_ibus_inst[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 448.840 500.000 449.440 ;
    END
  END io_ibus_inst[24]
  PIN io_ibus_inst[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 454.280 500.000 454.880 ;
    END
  END io_ibus_inst[25]
  PIN io_ibus_inst[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 460.400 500.000 461.000 ;
    END
  END io_ibus_inst[26]
  PIN io_ibus_inst[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 465.840 500.000 466.440 ;
    END
  END io_ibus_inst[27]
  PIN io_ibus_inst[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 471.960 500.000 472.560 ;
    END
  END io_ibus_inst[28]
  PIN io_ibus_inst[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 477.400 500.000 478.000 ;
    END
  END io_ibus_inst[29]
  PIN io_ibus_inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 321.000 500.000 321.600 ;
    END
  END io_ibus_inst[2]
  PIN io_ibus_inst[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 483.520 500.000 484.120 ;
    END
  END io_ibus_inst[30]
  PIN io_ibus_inst[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 488.960 500.000 489.560 ;
    END
  END io_ibus_inst[31]
  PIN io_ibus_inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 326.440 500.000 327.040 ;
    END
  END io_ibus_inst[3]
  PIN io_ibus_inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 332.560 500.000 333.160 ;
    END
  END io_ibus_inst[4]
  PIN io_ibus_inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 338.000 500.000 338.600 ;
    END
  END io_ibus_inst[5]
  PIN io_ibus_inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 344.120 500.000 344.720 ;
    END
  END io_ibus_inst[6]
  PIN io_ibus_inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 349.560 500.000 350.160 ;
    END
  END io_ibus_inst[7]
  PIN io_ibus_inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 355.680 500.000 356.280 ;
    END
  END io_ibus_inst[8]
  PIN io_ibus_inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 361.120 500.000 361.720 ;
    END
  END io_ibus_inst[9]
  PIN io_ibus_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 303.320 500.000 303.920 ;
    END
  END io_ibus_valid
  PIN io_irq_m1_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 497.800 500.000 498.400 ;
    END
  END io_irq_m1_irq
  PIN io_irq_m2_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END io_irq_m2_irq
  PIN io_irq_m3_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END io_irq_m3_irq
  PIN io_irq_spi_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 492.360 500.000 492.960 ;
    END
  END io_irq_spi_irq
  PIN io_irq_uart_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 495.080 500.000 495.680 ;
    END
  END io_irq_uart_irq
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 496.000 374.810 500.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.240 499.490 487.520 ;
      LAYER met2 ;
        RECT 6.990 495.720 124.470 498.285 ;
        RECT 125.310 495.720 374.250 498.285 ;
        RECT 375.090 495.720 499.470 498.285 ;
        RECT 6.990 4.280 499.470 495.720 ;
        RECT 6.990 1.515 249.590 4.280 ;
        RECT 250.430 1.515 499.470 4.280 ;
      LAYER met3 ;
        RECT 4.000 497.400 495.600 498.265 ;
        RECT 4.000 496.080 499.495 497.400 ;
        RECT 4.000 494.680 495.600 496.080 ;
        RECT 4.000 493.360 499.495 494.680 ;
        RECT 4.000 491.960 495.600 493.360 ;
        RECT 4.000 489.960 499.495 491.960 ;
        RECT 4.000 488.560 495.600 489.960 ;
        RECT 4.000 487.240 499.495 488.560 ;
        RECT 4.000 485.840 495.600 487.240 ;
        RECT 4.000 484.520 499.495 485.840 ;
        RECT 4.000 483.120 495.600 484.520 ;
        RECT 4.000 481.800 499.495 483.120 ;
        RECT 4.000 480.400 495.600 481.800 ;
        RECT 4.000 478.400 499.495 480.400 ;
        RECT 4.000 477.000 495.600 478.400 ;
        RECT 4.000 475.680 499.495 477.000 ;
        RECT 4.000 474.280 495.600 475.680 ;
        RECT 4.000 472.960 499.495 474.280 ;
        RECT 4.000 471.560 495.600 472.960 ;
        RECT 4.000 469.560 499.495 471.560 ;
        RECT 4.000 468.160 495.600 469.560 ;
        RECT 4.000 466.840 499.495 468.160 ;
        RECT 4.000 465.440 495.600 466.840 ;
        RECT 4.000 464.120 499.495 465.440 ;
        RECT 4.000 462.720 495.600 464.120 ;
        RECT 4.000 461.400 499.495 462.720 ;
        RECT 4.000 460.000 495.600 461.400 ;
        RECT 4.000 458.000 499.495 460.000 ;
        RECT 4.000 456.600 495.600 458.000 ;
        RECT 4.000 455.280 499.495 456.600 ;
        RECT 4.000 453.880 495.600 455.280 ;
        RECT 4.000 452.560 499.495 453.880 ;
        RECT 4.000 451.160 495.600 452.560 ;
        RECT 4.000 449.840 499.495 451.160 ;
        RECT 4.000 448.440 495.600 449.840 ;
        RECT 4.000 446.440 499.495 448.440 ;
        RECT 4.000 445.040 495.600 446.440 ;
        RECT 4.000 443.720 499.495 445.040 ;
        RECT 4.000 442.320 495.600 443.720 ;
        RECT 4.000 441.000 499.495 442.320 ;
        RECT 4.000 439.600 495.600 441.000 ;
        RECT 4.000 437.600 499.495 439.600 ;
        RECT 4.000 436.200 495.600 437.600 ;
        RECT 4.000 434.880 499.495 436.200 ;
        RECT 4.000 433.480 495.600 434.880 ;
        RECT 4.000 432.160 499.495 433.480 ;
        RECT 4.000 430.760 495.600 432.160 ;
        RECT 4.000 429.440 499.495 430.760 ;
        RECT 4.000 428.040 495.600 429.440 ;
        RECT 4.000 426.040 499.495 428.040 ;
        RECT 4.000 424.640 495.600 426.040 ;
        RECT 4.000 423.320 499.495 424.640 ;
        RECT 4.000 421.920 495.600 423.320 ;
        RECT 4.000 420.600 499.495 421.920 ;
        RECT 4.000 419.200 495.600 420.600 ;
        RECT 4.000 417.880 499.495 419.200 ;
        RECT 4.000 416.480 495.600 417.880 ;
        RECT 4.000 414.480 499.495 416.480 ;
        RECT 4.000 413.080 495.600 414.480 ;
        RECT 4.000 411.760 499.495 413.080 ;
        RECT 4.000 410.360 495.600 411.760 ;
        RECT 4.000 409.040 499.495 410.360 ;
        RECT 4.000 407.640 495.600 409.040 ;
        RECT 4.000 405.640 499.495 407.640 ;
        RECT 4.000 404.240 495.600 405.640 ;
        RECT 4.000 402.920 499.495 404.240 ;
        RECT 4.000 401.520 495.600 402.920 ;
        RECT 4.000 400.200 499.495 401.520 ;
        RECT 4.000 398.800 495.600 400.200 ;
        RECT 4.000 397.480 499.495 398.800 ;
        RECT 4.000 396.080 495.600 397.480 ;
        RECT 4.000 394.080 499.495 396.080 ;
        RECT 4.000 392.680 495.600 394.080 ;
        RECT 4.000 391.360 499.495 392.680 ;
        RECT 4.000 389.960 495.600 391.360 ;
        RECT 4.000 388.640 499.495 389.960 ;
        RECT 4.000 387.240 495.600 388.640 ;
        RECT 4.000 385.920 499.495 387.240 ;
        RECT 4.000 384.520 495.600 385.920 ;
        RECT 4.000 382.520 499.495 384.520 ;
        RECT 4.000 381.120 495.600 382.520 ;
        RECT 4.000 379.800 499.495 381.120 ;
        RECT 4.000 378.400 495.600 379.800 ;
        RECT 4.000 377.080 499.495 378.400 ;
        RECT 4.000 375.680 495.600 377.080 ;
        RECT 4.000 373.680 499.495 375.680 ;
        RECT 4.000 372.280 495.600 373.680 ;
        RECT 4.000 370.960 499.495 372.280 ;
        RECT 4.000 369.560 495.600 370.960 ;
        RECT 4.000 368.240 499.495 369.560 ;
        RECT 4.000 366.840 495.600 368.240 ;
        RECT 4.000 365.520 499.495 366.840 ;
        RECT 4.000 364.120 495.600 365.520 ;
        RECT 4.000 362.120 499.495 364.120 ;
        RECT 4.000 360.720 495.600 362.120 ;
        RECT 4.000 359.400 499.495 360.720 ;
        RECT 4.000 358.000 495.600 359.400 ;
        RECT 4.000 356.680 499.495 358.000 ;
        RECT 4.000 355.280 495.600 356.680 ;
        RECT 4.000 353.960 499.495 355.280 ;
        RECT 4.000 352.560 495.600 353.960 ;
        RECT 4.000 350.560 499.495 352.560 ;
        RECT 4.000 349.160 495.600 350.560 ;
        RECT 4.000 347.840 499.495 349.160 ;
        RECT 4.000 346.440 495.600 347.840 ;
        RECT 4.000 345.120 499.495 346.440 ;
        RECT 4.000 343.720 495.600 345.120 ;
        RECT 4.000 341.720 499.495 343.720 ;
        RECT 4.000 340.320 495.600 341.720 ;
        RECT 4.000 339.000 499.495 340.320 ;
        RECT 4.000 337.600 495.600 339.000 ;
        RECT 4.000 336.280 499.495 337.600 ;
        RECT 4.000 334.880 495.600 336.280 ;
        RECT 4.000 333.560 499.495 334.880 ;
        RECT 4.000 332.160 495.600 333.560 ;
        RECT 4.000 330.160 499.495 332.160 ;
        RECT 4.000 328.760 495.600 330.160 ;
        RECT 4.000 327.440 499.495 328.760 ;
        RECT 4.000 326.040 495.600 327.440 ;
        RECT 4.000 324.720 499.495 326.040 ;
        RECT 4.000 323.320 495.600 324.720 ;
        RECT 4.000 322.000 499.495 323.320 ;
        RECT 4.000 320.600 495.600 322.000 ;
        RECT 4.000 318.600 499.495 320.600 ;
        RECT 4.000 317.200 495.600 318.600 ;
        RECT 4.000 315.880 499.495 317.200 ;
        RECT 4.000 314.480 495.600 315.880 ;
        RECT 4.000 313.160 499.495 314.480 ;
        RECT 4.000 311.760 495.600 313.160 ;
        RECT 4.000 309.760 499.495 311.760 ;
        RECT 4.000 308.360 495.600 309.760 ;
        RECT 4.000 307.040 499.495 308.360 ;
        RECT 4.000 305.640 495.600 307.040 ;
        RECT 4.000 304.320 499.495 305.640 ;
        RECT 4.000 302.920 495.600 304.320 ;
        RECT 4.000 301.600 499.495 302.920 ;
        RECT 4.000 300.200 495.600 301.600 ;
        RECT 4.000 298.200 499.495 300.200 ;
        RECT 4.000 296.800 495.600 298.200 ;
        RECT 4.000 295.480 499.495 296.800 ;
        RECT 4.000 294.080 495.600 295.480 ;
        RECT 4.000 292.760 499.495 294.080 ;
        RECT 4.000 291.360 495.600 292.760 ;
        RECT 4.000 290.040 499.495 291.360 ;
        RECT 4.000 288.640 495.600 290.040 ;
        RECT 4.000 286.640 499.495 288.640 ;
        RECT 4.000 285.240 495.600 286.640 ;
        RECT 4.000 283.920 499.495 285.240 ;
        RECT 4.000 282.520 495.600 283.920 ;
        RECT 4.000 281.200 499.495 282.520 ;
        RECT 4.000 279.800 495.600 281.200 ;
        RECT 4.000 277.800 499.495 279.800 ;
        RECT 4.000 276.400 495.600 277.800 ;
        RECT 4.000 275.080 499.495 276.400 ;
        RECT 4.000 273.680 495.600 275.080 ;
        RECT 4.000 272.360 499.495 273.680 ;
        RECT 4.000 270.960 495.600 272.360 ;
        RECT 4.000 269.640 499.495 270.960 ;
        RECT 4.000 268.240 495.600 269.640 ;
        RECT 4.000 266.240 499.495 268.240 ;
        RECT 4.000 264.840 495.600 266.240 ;
        RECT 4.000 263.520 499.495 264.840 ;
        RECT 4.000 262.120 495.600 263.520 ;
        RECT 4.000 260.800 499.495 262.120 ;
        RECT 4.000 259.400 495.600 260.800 ;
        RECT 4.000 258.080 499.495 259.400 ;
        RECT 4.000 256.680 495.600 258.080 ;
        RECT 4.000 254.680 499.495 256.680 ;
        RECT 4.000 253.280 495.600 254.680 ;
        RECT 4.000 251.960 499.495 253.280 ;
        RECT 4.000 250.600 495.600 251.960 ;
        RECT 4.400 250.560 495.600 250.600 ;
        RECT 4.400 249.240 499.495 250.560 ;
        RECT 4.400 249.200 495.600 249.240 ;
        RECT 4.000 247.840 495.600 249.200 ;
        RECT 4.000 245.840 499.495 247.840 ;
        RECT 4.000 244.440 495.600 245.840 ;
        RECT 4.000 243.120 499.495 244.440 ;
        RECT 4.000 241.720 495.600 243.120 ;
        RECT 4.000 240.400 499.495 241.720 ;
        RECT 4.000 239.000 495.600 240.400 ;
        RECT 4.000 237.680 499.495 239.000 ;
        RECT 4.000 236.280 495.600 237.680 ;
        RECT 4.000 234.280 499.495 236.280 ;
        RECT 4.000 232.880 495.600 234.280 ;
        RECT 4.000 231.560 499.495 232.880 ;
        RECT 4.000 230.160 495.600 231.560 ;
        RECT 4.000 228.840 499.495 230.160 ;
        RECT 4.000 227.440 495.600 228.840 ;
        RECT 4.000 226.120 499.495 227.440 ;
        RECT 4.000 224.720 495.600 226.120 ;
        RECT 4.000 222.720 499.495 224.720 ;
        RECT 4.000 221.320 495.600 222.720 ;
        RECT 4.000 220.000 499.495 221.320 ;
        RECT 4.000 218.600 495.600 220.000 ;
        RECT 4.000 217.280 499.495 218.600 ;
        RECT 4.000 215.880 495.600 217.280 ;
        RECT 4.000 213.880 499.495 215.880 ;
        RECT 4.000 212.480 495.600 213.880 ;
        RECT 4.000 211.160 499.495 212.480 ;
        RECT 4.000 209.760 495.600 211.160 ;
        RECT 4.000 208.440 499.495 209.760 ;
        RECT 4.000 207.040 495.600 208.440 ;
        RECT 4.000 205.720 499.495 207.040 ;
        RECT 4.000 204.320 495.600 205.720 ;
        RECT 4.000 202.320 499.495 204.320 ;
        RECT 4.000 200.920 495.600 202.320 ;
        RECT 4.000 199.600 499.495 200.920 ;
        RECT 4.000 198.200 495.600 199.600 ;
        RECT 4.000 196.880 499.495 198.200 ;
        RECT 4.000 195.480 495.600 196.880 ;
        RECT 4.000 194.160 499.495 195.480 ;
        RECT 4.000 192.760 495.600 194.160 ;
        RECT 4.000 190.760 499.495 192.760 ;
        RECT 4.000 189.360 495.600 190.760 ;
        RECT 4.000 188.040 499.495 189.360 ;
        RECT 4.000 186.640 495.600 188.040 ;
        RECT 4.000 185.320 499.495 186.640 ;
        RECT 4.000 183.920 495.600 185.320 ;
        RECT 4.000 181.920 499.495 183.920 ;
        RECT 4.000 180.520 495.600 181.920 ;
        RECT 4.000 179.200 499.495 180.520 ;
        RECT 4.000 177.800 495.600 179.200 ;
        RECT 4.000 176.480 499.495 177.800 ;
        RECT 4.000 175.080 495.600 176.480 ;
        RECT 4.000 173.760 499.495 175.080 ;
        RECT 4.000 172.360 495.600 173.760 ;
        RECT 4.000 170.360 499.495 172.360 ;
        RECT 4.000 168.960 495.600 170.360 ;
        RECT 4.000 167.640 499.495 168.960 ;
        RECT 4.000 166.240 495.600 167.640 ;
        RECT 4.000 164.920 499.495 166.240 ;
        RECT 4.000 163.520 495.600 164.920 ;
        RECT 4.000 162.200 499.495 163.520 ;
        RECT 4.000 160.800 495.600 162.200 ;
        RECT 4.000 158.800 499.495 160.800 ;
        RECT 4.000 157.400 495.600 158.800 ;
        RECT 4.000 156.080 499.495 157.400 ;
        RECT 4.000 154.680 495.600 156.080 ;
        RECT 4.000 153.360 499.495 154.680 ;
        RECT 4.000 151.960 495.600 153.360 ;
        RECT 4.000 149.960 499.495 151.960 ;
        RECT 4.000 148.560 495.600 149.960 ;
        RECT 4.000 147.240 499.495 148.560 ;
        RECT 4.000 145.840 495.600 147.240 ;
        RECT 4.000 144.520 499.495 145.840 ;
        RECT 4.000 143.120 495.600 144.520 ;
        RECT 4.000 141.800 499.495 143.120 ;
        RECT 4.000 140.400 495.600 141.800 ;
        RECT 4.000 138.400 499.495 140.400 ;
        RECT 4.000 137.000 495.600 138.400 ;
        RECT 4.000 135.680 499.495 137.000 ;
        RECT 4.000 134.280 495.600 135.680 ;
        RECT 4.000 132.960 499.495 134.280 ;
        RECT 4.000 131.560 495.600 132.960 ;
        RECT 4.000 130.240 499.495 131.560 ;
        RECT 4.000 128.840 495.600 130.240 ;
        RECT 4.000 126.840 499.495 128.840 ;
        RECT 4.000 125.440 495.600 126.840 ;
        RECT 4.000 124.120 499.495 125.440 ;
        RECT 4.000 122.720 495.600 124.120 ;
        RECT 4.000 121.400 499.495 122.720 ;
        RECT 4.000 120.000 495.600 121.400 ;
        RECT 4.000 118.000 499.495 120.000 ;
        RECT 4.000 116.600 495.600 118.000 ;
        RECT 4.000 115.280 499.495 116.600 ;
        RECT 4.000 113.880 495.600 115.280 ;
        RECT 4.000 112.560 499.495 113.880 ;
        RECT 4.000 111.160 495.600 112.560 ;
        RECT 4.000 109.840 499.495 111.160 ;
        RECT 4.000 108.440 495.600 109.840 ;
        RECT 4.000 106.440 499.495 108.440 ;
        RECT 4.000 105.040 495.600 106.440 ;
        RECT 4.000 103.720 499.495 105.040 ;
        RECT 4.000 102.320 495.600 103.720 ;
        RECT 4.000 101.000 499.495 102.320 ;
        RECT 4.000 99.600 495.600 101.000 ;
        RECT 4.000 98.280 499.495 99.600 ;
        RECT 4.000 96.880 495.600 98.280 ;
        RECT 4.000 94.880 499.495 96.880 ;
        RECT 4.000 93.480 495.600 94.880 ;
        RECT 4.000 92.160 499.495 93.480 ;
        RECT 4.000 90.760 495.600 92.160 ;
        RECT 4.000 89.440 499.495 90.760 ;
        RECT 4.000 88.040 495.600 89.440 ;
        RECT 4.000 86.040 499.495 88.040 ;
        RECT 4.000 84.640 495.600 86.040 ;
        RECT 4.000 83.320 499.495 84.640 ;
        RECT 4.000 81.920 495.600 83.320 ;
        RECT 4.000 80.600 499.495 81.920 ;
        RECT 4.000 79.200 495.600 80.600 ;
        RECT 4.000 77.880 499.495 79.200 ;
        RECT 4.000 76.480 495.600 77.880 ;
        RECT 4.000 74.480 499.495 76.480 ;
        RECT 4.000 73.080 495.600 74.480 ;
        RECT 4.000 71.760 499.495 73.080 ;
        RECT 4.000 70.360 495.600 71.760 ;
        RECT 4.000 69.040 499.495 70.360 ;
        RECT 4.000 67.640 495.600 69.040 ;
        RECT 4.000 66.320 499.495 67.640 ;
        RECT 4.000 64.920 495.600 66.320 ;
        RECT 4.000 62.920 499.495 64.920 ;
        RECT 4.000 61.520 495.600 62.920 ;
        RECT 4.000 60.200 499.495 61.520 ;
        RECT 4.000 58.800 495.600 60.200 ;
        RECT 4.000 57.480 499.495 58.800 ;
        RECT 4.000 56.080 495.600 57.480 ;
        RECT 4.000 54.080 499.495 56.080 ;
        RECT 4.000 52.680 495.600 54.080 ;
        RECT 4.000 51.360 499.495 52.680 ;
        RECT 4.000 49.960 495.600 51.360 ;
        RECT 4.000 48.640 499.495 49.960 ;
        RECT 4.000 47.240 495.600 48.640 ;
        RECT 4.000 45.920 499.495 47.240 ;
        RECT 4.000 44.520 495.600 45.920 ;
        RECT 4.000 42.520 499.495 44.520 ;
        RECT 4.000 41.120 495.600 42.520 ;
        RECT 4.000 39.800 499.495 41.120 ;
        RECT 4.000 38.400 495.600 39.800 ;
        RECT 4.000 37.080 499.495 38.400 ;
        RECT 4.000 35.680 495.600 37.080 ;
        RECT 4.000 34.360 499.495 35.680 ;
        RECT 4.000 32.960 495.600 34.360 ;
        RECT 4.000 30.960 499.495 32.960 ;
        RECT 4.000 29.560 495.600 30.960 ;
        RECT 4.000 28.240 499.495 29.560 ;
        RECT 4.000 26.840 495.600 28.240 ;
        RECT 4.000 25.520 499.495 26.840 ;
        RECT 4.000 24.120 495.600 25.520 ;
        RECT 4.000 22.120 499.495 24.120 ;
        RECT 4.000 20.720 495.600 22.120 ;
        RECT 4.000 19.400 499.495 20.720 ;
        RECT 4.000 18.000 495.600 19.400 ;
        RECT 4.000 16.680 499.495 18.000 ;
        RECT 4.000 15.280 495.600 16.680 ;
        RECT 4.000 13.960 499.495 15.280 ;
        RECT 4.000 12.560 495.600 13.960 ;
        RECT 4.000 10.560 499.495 12.560 ;
        RECT 4.000 9.160 495.600 10.560 ;
        RECT 4.000 7.840 499.495 9.160 ;
        RECT 4.000 6.440 495.600 7.840 ;
        RECT 4.000 5.120 499.495 6.440 ;
        RECT 4.000 3.720 495.600 5.120 ;
        RECT 4.000 2.400 499.495 3.720 ;
        RECT 4.000 1.535 495.600 2.400 ;
      LAYER met4 ;
        RECT 17.775 11.735 20.640 483.305 ;
        RECT 23.040 11.735 97.440 483.305 ;
        RECT 99.840 11.735 174.240 483.305 ;
        RECT 176.640 11.735 251.040 483.305 ;
        RECT 253.440 11.735 327.840 483.305 ;
        RECT 330.240 11.735 404.640 483.305 ;
        RECT 407.040 11.735 481.440 483.305 ;
        RECT 483.840 11.735 490.985 483.305 ;
  END
END Core
END LIBRARY

