module WBM_DBus( // @[:@3196.2]
  input  [31:0] io_dbus_addr, // @[:@3199.4]
  input  [31:0] io_dbus_wdata, // @[:@3199.4]
  output [31:0] io_dbus_rdata, // @[:@3199.4]
  input         io_dbus_rd_en, // @[:@3199.4]
  input         io_dbus_wr_en, // @[:@3199.4]
  input  [1:0]  io_dbus_st_type, // @[:@3199.4]
  input  [2:0]  io_dbus_ld_type, // @[:@3199.4]
  output        io_dbus_valid, // @[:@3199.4]
  output [15:0] io_wbm_m2s_addr, // @[:@3199.4]
  output [31:0] io_wbm_m2s_data, // @[:@3199.4]
  output        io_wbm_m2s_we, // @[:@3199.4]
  output [3:0]  io_wbm_m2s_sel, // @[:@3199.4]
  output        io_wbm_m2s_stb, // @[:@3199.4]
  input         io_wbm_ack_i, // @[:@3199.4]
  input  [31:0] io_wbm_data_i // @[:@3199.4]
);
  wire  _T_39; // @[wbm_dbus.scala 35:19:@3203.4]
  wire  _T_40; // @[wbm_dbus.scala 38:26:@3208.6]
  wire  _T_41; // @[wbm_dbus.scala 41:26:@3213.8]
  wire [3:0] _GEN_0; // @[wbm_dbus.scala 41:46:@3214.8]
  wire [3:0] _GEN_1; // @[wbm_dbus.scala 38:47:@3209.6]
  wire [3:0] st_sel_vec; // @[wbm_dbus.scala 35:40:@3204.4]
  wire [1:0] ld_align; // @[wbm_dbus.scala 46:30:@3217.4]
  wire  _T_44; // @[wbm_dbus.scala 51:16:@3220.4]
  wire  _T_45; // @[wbm_dbus.scala 54:23:@3225.6]
  wire  _T_46; // @[wbm_dbus.scala 54:54:@3226.6]
  wire  _T_47; // @[wbm_dbus.scala 54:43:@3227.6]
  wire  _T_48; // @[wbm_dbus.scala 55:34:@3229.8]
  wire [3:0] _T_49; // @[wbm_dbus.scala 55:25:@3230.8]
  wire  _T_50; // @[wbm_dbus.scala 57:23:@3234.8]
  wire  _T_51; // @[wbm_dbus.scala 57:54:@3235.8]
  wire  _T_52; // @[wbm_dbus.scala 57:43:@3236.8]
  wire  _T_54; // @[wbm_dbus.scala 58:21:@3238.10]
  wire  _T_56; // @[wbm_dbus.scala 60:27:@3243.12]
  wire  _T_58; // @[wbm_dbus.scala 62:27:@3248.14]
  wire [3:0] _GEN_3; // @[wbm_dbus.scala 62:37:@3249.14]
  wire [3:0] _GEN_4; // @[wbm_dbus.scala 60:37:@3244.12]
  wire [3:0] _GEN_5; // @[wbm_dbus.scala 58:32:@3239.10]
  wire [3:0] _GEN_6; // @[wbm_dbus.scala 57:75:@3237.8]
  wire [3:0] _GEN_7; // @[wbm_dbus.scala 54:76:@3228.6]
  wire [3:0] ld_sel_vec; // @[wbm_dbus.scala 51:37:@3221.4]
  wire  _T_61; // @[wbm_dbus.scala 74:37:@3260.4]
  assign _T_39 = io_dbus_st_type == 2'h1; // @[wbm_dbus.scala 35:19:@3203.4]
  assign _T_40 = io_dbus_st_type == 2'h2; // @[wbm_dbus.scala 38:26:@3208.6]
  assign _T_41 = io_dbus_st_type == 2'h3; // @[wbm_dbus.scala 41:26:@3213.8]
  assign _GEN_0 = _T_41 ? 4'h1 : 4'h0; // @[wbm_dbus.scala 41:46:@3214.8]
  assign _GEN_1 = _T_40 ? 4'h3 : _GEN_0; // @[wbm_dbus.scala 38:47:@3209.6]
  assign st_sel_vec = _T_39 ? 4'hf : _GEN_1; // @[wbm_dbus.scala 35:40:@3204.4]
  assign ld_align = io_dbus_addr[1:0]; // @[wbm_dbus.scala 46:30:@3217.4]
  assign _T_44 = io_dbus_ld_type == 3'h1; // @[wbm_dbus.scala 51:16:@3220.4]
  assign _T_45 = io_dbus_ld_type == 3'h2; // @[wbm_dbus.scala 54:23:@3225.6]
  assign _T_46 = io_dbus_ld_type == 3'h4; // @[wbm_dbus.scala 54:54:@3226.6]
  assign _T_47 = _T_45 | _T_46; // @[wbm_dbus.scala 54:43:@3227.6]
  assign _T_48 = ld_align[1]; // @[wbm_dbus.scala 55:34:@3229.8]
  assign _T_49 = _T_48 ? 4'hc : 4'h3; // @[wbm_dbus.scala 55:25:@3230.8]
  assign _T_50 = io_dbus_ld_type == 3'h3; // @[wbm_dbus.scala 57:23:@3234.8]
  assign _T_51 = io_dbus_ld_type == 3'h5; // @[wbm_dbus.scala 57:54:@3235.8]
  assign _T_52 = _T_50 | _T_51; // @[wbm_dbus.scala 57:43:@3236.8]
  assign _T_54 = ld_align == 2'h3; // @[wbm_dbus.scala 58:21:@3238.10]
  assign _T_56 = ld_align == 2'h2; // @[wbm_dbus.scala 60:27:@3243.12]
  assign _T_58 = ld_align == 2'h1; // @[wbm_dbus.scala 62:27:@3248.14]
  assign _GEN_3 = _T_58 ? 4'h2 : 4'h1; // @[wbm_dbus.scala 62:37:@3249.14]
  assign _GEN_4 = _T_56 ? 4'h4 : _GEN_3; // @[wbm_dbus.scala 60:37:@3244.12]
  assign _GEN_5 = _T_54 ? 4'h8 : _GEN_4; // @[wbm_dbus.scala 58:32:@3239.10]
  assign _GEN_6 = _T_52 ? _GEN_5 : 4'h0; // @[wbm_dbus.scala 57:75:@3237.8]
  assign _GEN_7 = _T_47 ? _T_49 : _GEN_6; // @[wbm_dbus.scala 54:76:@3228.6]
  assign ld_sel_vec = _T_44 ? 4'hf : _GEN_7; // @[wbm_dbus.scala 51:37:@3221.4]
  assign _T_61 = io_dbus_st_type != 2'h0; // @[wbm_dbus.scala 74:37:@3260.4]
  assign io_dbus_rdata = io_wbm_data_i; // @[wbm_dbus.scala 78:19:@3268.4]
  assign io_dbus_valid = io_wbm_ack_i; // @[wbm_dbus.scala 79:19:@3269.4]
  assign io_wbm_m2s_addr = io_dbus_addr[15:0]; // @[wbm_dbus.scala 71:19:@3257.4]
  assign io_wbm_m2s_data = io_dbus_wdata; // @[wbm_dbus.scala 72:19:@3258.4]
  assign io_wbm_m2s_we = io_dbus_wr_en; // @[wbm_dbus.scala 73:19:@3259.4]
  assign io_wbm_m2s_sel = _T_61 ? st_sel_vec : ld_sel_vec; // @[wbm_dbus.scala 74:19:@3262.4]
  assign io_wbm_m2s_stb = io_dbus_rd_en | io_dbus_wr_en; // @[wbm_dbus.scala 75:19:@3266.4]
endmodule
